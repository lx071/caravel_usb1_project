magic
tech sky130A
magscale 1 2
timestamp 1698803719
<< viali >>
rect 432705 3485 432739 3519
rect 433901 3485 433935 3519
rect 337669 3417 337703 3451
rect 527189 3417 527223 3451
rect 248705 3349 248739 3383
rect 336289 3349 336323 3383
rect 338865 3349 338899 3383
rect 339877 3349 339911 3383
rect 433349 3349 433383 3383
rect 434453 3349 434487 3383
rect 78873 3145 78907 3179
rect 171609 3145 171643 3179
rect 218069 3145 218103 3179
rect 338405 3145 338439 3179
rect 357081 3145 357115 3179
rect 403449 3145 403483 3179
rect 588921 3145 588955 3179
rect 681749 3145 681783 3179
rect 278973 3077 279007 3111
rect 295717 3077 295751 3111
rect 387993 3077 388027 3111
rect 434269 3077 434303 3111
rect 449909 3077 449943 3111
rect 496185 3077 496219 3111
rect 525625 3077 525659 3111
rect 248981 3009 249015 3043
rect 264345 3009 264379 3043
rect 279617 3009 279651 3043
rect 279893 3009 279927 3043
rect 295165 3009 295199 3043
rect 310713 3009 310747 3043
rect 337393 3009 337427 3043
rect 339049 3009 339083 3043
rect 339601 3009 339635 3043
rect 342085 3009 342119 3043
rect 431417 3009 431451 3043
rect 432981 3009 433015 3043
rect 433533 3009 433567 3043
rect 434821 3009 434855 3043
rect 463893 3009 463927 3043
rect 479349 3009 479383 3043
rect 525901 3009 525935 3043
rect 527557 3009 527591 3043
rect 294429 2941 294463 2975
rect 336841 2941 336875 2975
rect 341533 2941 341567 2975
rect 431877 2941 431911 2975
rect 464445 2941 464479 2975
rect 479901 2941 479935 2975
rect 527005 2941 527039 2975
rect 573465 2941 573499 2975
rect 372629 2873 372663 2907
rect 136465 2805 136499 2839
rect 187709 2805 187743 2839
rect 203073 2805 203107 2839
rect 249257 2805 249291 2839
rect 277225 2805 277259 2839
rect 292681 2805 292715 2839
rect 323409 2805 323443 2839
rect 324513 2805 324547 2839
rect 326169 2805 326203 2839
rect 331689 2805 331723 2839
rect 333253 2805 333287 2839
rect 334817 2805 334851 2839
rect 335737 2805 335771 2839
rect 340245 2805 340279 2839
rect 342729 2805 342763 2839
rect 367477 2805 367511 2839
rect 370881 2805 370915 2839
rect 382841 2805 382875 2839
rect 386429 2805 386463 2839
rect 417341 2805 417375 2839
rect 418905 2805 418939 2839
rect 430773 2805 430807 2839
rect 435465 2805 435499 2839
rect 463249 2805 463283 2839
rect 465273 2805 465307 2839
rect 478705 2805 478739 2839
rect 480729 2805 480763 2839
rect 511641 2805 511675 2839
rect 528201 2805 528235 2839
rect 529029 2805 529063 2839
rect 558101 2805 558135 2839
rect 604469 2805 604503 2839
rect 619833 2805 619867 2839
rect 650745 2805 650779 2839
rect 666201 2805 666235 2839
rect 1869 2601 1903 2635
rect 17325 2601 17359 2635
rect 48237 2601 48271 2635
rect 63693 2601 63727 2635
rect 94605 2601 94639 2635
rect 98009 2601 98043 2635
rect 187341 2601 187375 2635
rect 202797 2601 202831 2635
rect 233709 2601 233743 2635
rect 248061 2601 248095 2635
rect 249165 2601 249199 2635
rect 295533 2601 295567 2635
rect 481005 2601 481039 2635
rect 511917 2601 511951 2635
rect 604653 2601 604687 2635
rect 620109 2601 620143 2635
rect 626089 2601 626123 2635
rect 681933 2601 681967 2635
rect 32965 2533 32999 2567
rect 48973 2533 49007 2567
rect 140973 2533 141007 2567
rect 156429 2533 156463 2567
rect 218253 2533 218287 2567
rect 372813 2533 372847 2567
rect 388269 2533 388303 2567
rect 525073 2533 525107 2567
rect 635749 2533 635783 2567
rect 651021 2533 651055 2567
rect 666477 2533 666511 2567
rect 41061 2465 41095 2499
rect 134717 2465 134751 2499
rect 190561 2465 190595 2499
rect 206753 2465 206787 2499
rect 385877 2465 385911 2499
rect 418077 2465 418111 2499
rect 478797 2465 478831 2499
rect 510813 2465 510847 2499
rect 570797 2465 570831 2499
rect 572545 2465 572579 2499
rect 2053 2397 2087 2431
rect 17509 2397 17543 2431
rect 32781 2397 32815 2431
rect 33425 2397 33459 2431
rect 40785 2397 40819 2431
rect 48421 2397 48455 2431
rect 63877 2397 63911 2431
rect 79333 2397 79367 2431
rect 94789 2397 94823 2431
rect 97365 2397 97399 2431
rect 110245 2397 110279 2431
rect 112821 2397 112855 2431
rect 125517 2397 125551 2431
rect 126161 2397 126195 2431
rect 135453 2397 135487 2431
rect 136557 2397 136591 2431
rect 138121 2397 138155 2431
rect 141157 2397 141191 2431
rect 143733 2397 143767 2431
rect 156613 2397 156647 2431
rect 159189 2397 159223 2431
rect 172069 2397 172103 2431
rect 187525 2397 187559 2431
rect 188905 2397 188939 2431
rect 189549 2397 189583 2431
rect 190837 2397 190871 2431
rect 202981 2397 203015 2431
rect 204177 2397 204211 2431
rect 206201 2397 206235 2431
rect 218437 2397 218471 2431
rect 233893 2397 233927 2431
rect 246773 2397 246807 2431
rect 249349 2397 249383 2431
rect 264805 2397 264839 2431
rect 273085 2397 273119 2431
rect 273361 2397 273395 2431
rect 275293 2397 275327 2431
rect 277409 2397 277443 2431
rect 280261 2397 280295 2431
rect 288541 2397 288575 2431
rect 290657 2397 290691 2431
rect 292865 2397 292899 2431
rect 294429 2397 294463 2431
rect 295717 2397 295751 2431
rect 311173 2397 311207 2431
rect 321569 2397 321603 2431
rect 323593 2397 323627 2431
rect 324789 2397 324823 2431
rect 326629 2397 326663 2431
rect 331597 2397 331631 2431
rect 333069 2397 333103 2431
rect 334633 2397 334667 2431
rect 335737 2397 335771 2431
rect 336473 2397 336507 2431
rect 338221 2397 338255 2431
rect 339601 2397 339635 2431
rect 340245 2397 340279 2431
rect 342085 2397 342119 2431
rect 342545 2397 342579 2431
rect 357449 2397 357483 2431
rect 367753 2397 367787 2431
rect 369869 2397 369903 2431
rect 371157 2397 371191 2431
rect 371709 2397 371743 2431
rect 372997 2397 373031 2431
rect 383117 2397 383151 2431
rect 385325 2397 385359 2431
rect 386613 2397 386647 2431
rect 388453 2397 388487 2431
rect 403909 2397 403943 2431
rect 416237 2397 416271 2431
rect 417525 2397 417559 2431
rect 419365 2397 419399 2431
rect 428473 2397 428507 2431
rect 430313 2397 430347 2431
rect 431693 2397 431727 2431
rect 432245 2397 432279 2431
rect 433441 2397 433475 2431
rect 434821 2397 434855 2431
rect 435925 2397 435959 2431
rect 462513 2397 462547 2431
rect 465733 2397 465767 2431
rect 477969 2397 478003 2431
rect 481189 2397 481223 2431
rect 496645 2397 496679 2431
rect 509709 2397 509743 2431
rect 510261 2397 510295 2431
rect 512101 2397 512135 2431
rect 525717 2397 525751 2431
rect 526269 2397 526303 2431
rect 527557 2397 527591 2431
rect 528845 2397 528879 2431
rect 530317 2397 530351 2431
rect 542829 2397 542863 2431
rect 543473 2397 543507 2431
rect 555893 2397 555927 2431
rect 558469 2397 558503 2431
rect 571349 2397 571383 2431
rect 573925 2397 573959 2431
rect 589381 2397 589415 2431
rect 604837 2397 604871 2431
rect 620293 2397 620327 2431
rect 623329 2397 623363 2431
rect 625445 2397 625479 2431
rect 635565 2397 635599 2431
rect 636209 2397 636243 2431
rect 651205 2397 651239 2431
rect 666661 2397 666695 2431
rect 682117 2397 682151 2431
rect 64429 2329 64463 2363
rect 96813 2329 96847 2363
rect 112269 2329 112303 2363
rect 136005 2329 136039 2363
rect 136833 2329 136867 2363
rect 143181 2329 143215 2363
rect 158637 2329 158671 2363
rect 188629 2329 188663 2363
rect 203901 2329 203935 2363
rect 205925 2329 205959 2363
rect 247049 2329 247083 2363
rect 275569 2329 275603 2363
rect 277685 2329 277719 2363
rect 288817 2329 288851 2363
rect 290197 2329 290231 2363
rect 290933 2329 290967 2363
rect 293417 2329 293451 2363
rect 322121 2329 322155 2363
rect 324145 2329 324179 2363
rect 325341 2329 325375 2363
rect 331321 2329 331355 2363
rect 332609 2329 332643 2363
rect 334081 2329 334115 2363
rect 335461 2329 335495 2363
rect 337025 2329 337059 2363
rect 337669 2329 337703 2363
rect 339049 2329 339083 2363
rect 340797 2329 340831 2363
rect 368305 2329 368339 2363
rect 370421 2329 370455 2363
rect 383669 2329 383703 2363
rect 387165 2329 387199 2363
rect 416789 2329 416823 2363
rect 428197 2329 428231 2363
rect 429761 2329 429795 2363
rect 432889 2329 432923 2363
rect 435373 2329 435407 2363
rect 450185 2329 450219 2363
rect 463341 2329 463375 2363
rect 528293 2329 528327 2363
rect 529765 2329 529799 2363
rect 557089 2329 557123 2363
rect 623053 2329 623087 2363
rect 624893 2329 624927 2363
rect 2605 2261 2639 2295
rect 18061 2261 18095 2295
rect 79149 2261 79183 2295
rect 95341 2261 95375 2295
rect 110061 2261 110095 2295
rect 110705 2261 110739 2295
rect 113465 2261 113499 2295
rect 125701 2261 125735 2295
rect 138305 2261 138339 2295
rect 141709 2261 141743 2295
rect 144377 2261 144411 2295
rect 157165 2261 157199 2295
rect 159833 2261 159867 2295
rect 171885 2261 171919 2295
rect 191389 2261 191423 2295
rect 205005 2261 205039 2295
rect 234353 2261 234387 2295
rect 246221 2261 246255 2295
rect 264621 2261 264655 2295
rect 272533 2261 272567 2295
rect 274741 2261 274775 2295
rect 278973 2261 279007 2295
rect 280077 2261 280111 2295
rect 287989 2261 288023 2295
rect 310989 2261 311023 2295
rect 320925 2261 320959 2295
rect 326445 2261 326479 2295
rect 341901 2261 341935 2295
rect 357357 2261 357391 2295
rect 369133 2261 369167 2295
rect 384589 2261 384623 2295
rect 403725 2261 403759 2295
rect 415501 2261 415535 2295
rect 419181 2261 419215 2295
rect 429117 2261 429151 2295
rect 430957 2261 430991 2295
rect 434637 2261 434671 2295
rect 436845 2261 436879 2295
rect 450093 2261 450127 2295
rect 461869 2261 461903 2295
rect 465549 2261 465583 2295
rect 477325 2261 477359 2295
rect 496461 2261 496495 2295
rect 527373 2261 527407 2295
rect 530961 2261 530995 2295
rect 543013 2261 543047 2295
rect 555341 2261 555375 2295
rect 558285 2261 558319 2295
rect 573741 2261 573775 2295
rect 589197 2261 589231 2295
<< metal1 >>
rect 74 9228 130 10000
rect 1854 9228 1860 9240
rect 74 9200 1860 9228
rect 1854 9188 1860 9200
rect 1912 9188 1918 9240
rect 15374 9228 15430 10000
rect 16574 9228 16580 9240
rect 15374 9200 16580 9228
rect 16574 9188 16580 9200
rect 16632 9188 16638 9240
rect 30674 9228 30730 10000
rect 31754 9228 31760 9240
rect 30674 9200 31760 9228
rect 31754 9188 31760 9200
rect 31812 9188 31818 9240
rect 45974 9228 46030 10000
rect 45940 9200 46030 9228
rect 61274 9228 61330 10000
rect 62022 9228 62028 9240
rect 61274 9200 62028 9228
rect 45940 9160 45968 9200
rect 62022 9188 62028 9200
rect 62080 9188 62086 9240
rect 76574 9228 76630 10000
rect 76926 9228 76932 9240
rect 76574 9200 76932 9228
rect 76926 9188 76932 9200
rect 76984 9188 76990 9240
rect 91874 9228 91930 10000
rect 107174 9228 107230 10000
rect 107562 9228 107568 9240
rect 91874 9200 91968 9228
rect 107174 9200 107568 9228
rect 91940 9160 91968 9200
rect 107562 9188 107568 9200
rect 107620 9188 107626 9240
rect 122474 9228 122530 10000
rect 122742 9228 122748 9240
rect 122474 9200 122748 9228
rect 122742 9188 122748 9200
rect 122800 9188 122806 9240
rect 137774 9228 137830 10000
rect 153074 9228 153130 10000
rect 168374 9228 168430 10000
rect 169662 9228 169668 9240
rect 137774 9200 137876 9228
rect 153074 9200 153148 9228
rect 168374 9200 169668 9228
rect 137848 9160 137876 9200
rect 153120 9160 153148 9200
rect 169662 9188 169668 9200
rect 169720 9188 169726 9240
rect 183674 9228 183730 10000
rect 184842 9228 184848 9240
rect 183674 9200 184848 9228
rect 184842 9188 184848 9200
rect 184900 9188 184906 9240
rect 198974 9228 199030 10000
rect 198936 9200 199030 9228
rect 214274 9228 214330 10000
rect 215202 9228 215208 9240
rect 214274 9200 215208 9228
rect 45940 9132 46014 9160
rect 45986 8956 46014 9132
rect 91894 9132 91968 9160
rect 137802 9132 137876 9160
rect 153074 9132 153148 9160
rect 198936 9160 198964 9200
rect 215202 9188 215208 9200
rect 215260 9188 215266 9240
rect 229574 9228 229630 10000
rect 230382 9228 230388 9240
rect 229574 9200 230388 9228
rect 230382 9188 230388 9200
rect 230440 9188 230446 9240
rect 244874 9228 244930 10000
rect 244844 9200 244930 9228
rect 260174 9228 260230 10000
rect 260466 9228 260472 9240
rect 260174 9200 260472 9228
rect 244844 9160 244872 9200
rect 260466 9188 260472 9200
rect 260524 9188 260530 9240
rect 275474 9228 275530 10000
rect 275922 9228 275928 9240
rect 275474 9200 275928 9228
rect 275922 9188 275928 9200
rect 275980 9188 275986 9240
rect 290774 9228 290830 10000
rect 306074 9228 306130 10000
rect 290752 9200 290830 9228
rect 306024 9200 306130 9228
rect 321374 9228 321430 10000
rect 321462 9228 321468 9240
rect 321374 9200 321468 9228
rect 290752 9160 290780 9200
rect 306024 9160 306052 9200
rect 321462 9188 321468 9200
rect 321520 9188 321526 9240
rect 336674 9228 336730 10000
rect 336826 9228 336832 9240
rect 336674 9200 336832 9228
rect 336826 9188 336832 9200
rect 336884 9188 336890 9240
rect 351974 9228 352030 10000
rect 367274 9228 367330 10000
rect 368382 9228 368388 9240
rect 351974 9200 352052 9228
rect 367274 9200 368388 9228
rect 352024 9160 352052 9200
rect 368382 9188 368388 9200
rect 368440 9188 368446 9240
rect 382574 9228 382630 10000
rect 383562 9228 383568 9240
rect 382574 9200 383568 9228
rect 383562 9188 383568 9200
rect 383620 9188 383626 9240
rect 397874 9228 397930 10000
rect 397840 9200 397930 9228
rect 413174 9228 413230 10000
rect 413922 9228 413928 9240
rect 413174 9200 413928 9228
rect 198936 9132 199010 9160
rect 244844 9132 244918 9160
rect 290752 9132 290826 9160
rect 306024 9132 306116 9160
rect 46934 8956 46940 8968
rect 45986 8928 46940 8956
rect 46934 8916 46940 8928
rect 46992 8916 46998 8968
rect 91894 8956 91922 9132
rect 92382 8956 92388 8968
rect 91894 8928 92388 8956
rect 92382 8916 92388 8928
rect 92440 8916 92446 8968
rect 137802 8956 137830 9132
rect 153074 8968 153102 9132
rect 137922 8956 137928 8968
rect 137802 8928 137928 8956
rect 137922 8916 137928 8928
rect 137980 8916 137986 8968
rect 153074 8928 153108 8968
rect 153102 8916 153108 8928
rect 153160 8916 153166 8968
rect 198982 8956 199010 9132
rect 200022 8956 200028 8968
rect 198982 8928 200028 8956
rect 200022 8916 200028 8928
rect 200080 8916 200086 8968
rect 244890 8956 244918 9132
rect 245562 8956 245568 8968
rect 244890 8928 245568 8956
rect 245562 8916 245568 8928
rect 245620 8916 245626 8968
rect 290798 8956 290826 9132
rect 291102 8956 291108 8968
rect 290798 8928 291108 8956
rect 291102 8916 291108 8928
rect 291160 8916 291166 8968
rect 306088 8956 306116 9132
rect 351978 9132 352052 9160
rect 397840 9160 397868 9200
rect 413922 9188 413928 9200
rect 413980 9188 413986 9240
rect 428474 9228 428530 10000
rect 429102 9228 429108 9240
rect 428474 9200 429108 9228
rect 429102 9188 429108 9200
rect 429160 9188 429166 9240
rect 443774 9228 443830 10000
rect 443748 9200 443830 9228
rect 459074 9228 459130 10000
rect 459462 9228 459468 9240
rect 459074 9200 459468 9228
rect 443748 9160 443776 9200
rect 459462 9188 459468 9200
rect 459520 9188 459526 9240
rect 474374 9228 474430 10000
rect 474642 9228 474648 9240
rect 474374 9200 474648 9228
rect 474642 9188 474648 9200
rect 474700 9188 474706 9240
rect 489674 9228 489730 10000
rect 504974 9228 505030 10000
rect 520274 9228 520330 10000
rect 520918 9228 520924 9240
rect 489674 9200 489776 9228
rect 504974 9200 505048 9228
rect 520274 9200 520924 9228
rect 489748 9160 489776 9200
rect 505020 9160 505048 9200
rect 520918 9188 520924 9200
rect 520976 9188 520982 9240
rect 535574 9228 535630 10000
rect 536742 9228 536748 9240
rect 535574 9200 536748 9228
rect 536742 9188 536748 9200
rect 536800 9188 536806 9240
rect 550874 9228 550930 10000
rect 550836 9200 550930 9228
rect 566174 9228 566230 10000
rect 567102 9228 567108 9240
rect 566174 9200 567108 9228
rect 397840 9132 397914 9160
rect 443748 9132 443822 9160
rect 306282 8956 306288 8968
rect 306088 8928 306288 8956
rect 306282 8916 306288 8928
rect 306340 8916 306346 8968
rect 351978 8888 352006 9132
rect 353202 8888 353208 8900
rect 351978 8860 353208 8888
rect 353202 8848 353208 8860
rect 353260 8848 353266 8900
rect 397886 8888 397914 9132
rect 443794 8956 443822 9132
rect 489702 9132 489776 9160
rect 504974 9132 505048 9160
rect 550836 9160 550864 9200
rect 567102 9188 567108 9200
rect 567160 9188 567166 9240
rect 581474 9228 581530 10000
rect 582282 9228 582288 9240
rect 581474 9200 582288 9228
rect 582282 9188 582288 9200
rect 582340 9188 582346 9240
rect 596774 9228 596830 10000
rect 612074 9228 612130 10000
rect 612642 9228 612648 9240
rect 596774 9200 596864 9228
rect 612074 9200 612648 9228
rect 596836 9160 596864 9200
rect 612642 9188 612648 9200
rect 612700 9188 612706 9240
rect 627374 9228 627430 10000
rect 627638 9228 627644 9240
rect 627374 9200 627644 9228
rect 627638 9188 627644 9200
rect 627696 9188 627702 9240
rect 642674 9228 642730 10000
rect 657974 9228 658030 10000
rect 642652 9200 642730 9228
rect 657924 9200 658030 9228
rect 673274 9228 673330 10000
rect 673362 9228 673368 9240
rect 673274 9200 673368 9228
rect 550836 9132 550910 9160
rect 444098 8956 444104 8968
rect 443794 8928 444104 8956
rect 444098 8916 444104 8928
rect 444156 8916 444162 8968
rect 489702 8956 489730 9132
rect 504974 8968 505002 9132
rect 489822 8956 489828 8968
rect 489702 8928 489828 8956
rect 489822 8916 489828 8928
rect 489880 8916 489886 8968
rect 504974 8928 505008 8968
rect 505002 8916 505008 8928
rect 505060 8916 505066 8968
rect 398742 8888 398748 8900
rect 397886 8860 398748 8888
rect 398742 8848 398748 8860
rect 398800 8848 398806 8900
rect 550882 8888 550910 9132
rect 596790 9132 596864 9160
rect 642652 9160 642680 9200
rect 657924 9160 657952 9200
rect 673362 9188 673368 9200
rect 673420 9188 673426 9240
rect 642652 9132 642726 9160
rect 657924 9132 658016 9160
rect 596790 8956 596818 9132
rect 597278 8956 597284 8968
rect 596790 8928 597284 8956
rect 597278 8916 597284 8928
rect 597336 8916 597342 8968
rect 642698 8956 642726 9132
rect 643002 8956 643008 8968
rect 642698 8928 643008 8956
rect 643002 8916 643008 8928
rect 643060 8916 643066 8968
rect 657988 8956 658016 9132
rect 658182 8956 658188 8968
rect 657988 8928 658188 8956
rect 658182 8916 658188 8928
rect 658240 8916 658246 8968
rect 551922 8888 551928 8900
rect 550882 8860 551928 8888
rect 551922 8848 551928 8860
rect 551980 8848 551986 8900
rect 1104 7642 682824 7664
rect 1104 7590 86825 7642
rect 86877 7590 86889 7642
rect 86941 7590 86953 7642
rect 87005 7590 87017 7642
rect 87069 7590 87081 7642
rect 87133 7590 257255 7642
rect 257307 7590 257319 7642
rect 257371 7590 257383 7642
rect 257435 7590 257447 7642
rect 257499 7590 257511 7642
rect 257563 7590 427685 7642
rect 427737 7590 427749 7642
rect 427801 7590 427813 7642
rect 427865 7590 427877 7642
rect 427929 7590 427941 7642
rect 427993 7590 598115 7642
rect 598167 7590 598179 7642
rect 598231 7590 598243 7642
rect 598295 7590 598307 7642
rect 598359 7590 598371 7642
rect 598423 7590 682824 7642
rect 1104 7568 682824 7590
rect 1104 7098 682824 7120
rect 1104 7046 86165 7098
rect 86217 7046 86229 7098
rect 86281 7046 86293 7098
rect 86345 7046 86357 7098
rect 86409 7046 86421 7098
rect 86473 7046 256595 7098
rect 256647 7046 256659 7098
rect 256711 7046 256723 7098
rect 256775 7046 256787 7098
rect 256839 7046 256851 7098
rect 256903 7046 427025 7098
rect 427077 7046 427089 7098
rect 427141 7046 427153 7098
rect 427205 7046 427217 7098
rect 427269 7046 427281 7098
rect 427333 7046 597455 7098
rect 597507 7046 597519 7098
rect 597571 7046 597583 7098
rect 597635 7046 597647 7098
rect 597699 7046 597711 7098
rect 597763 7046 682824 7098
rect 1104 7024 682824 7046
rect 62022 6808 62028 6860
rect 62080 6848 62086 6860
rect 63678 6848 63684 6860
rect 62080 6820 63684 6848
rect 62080 6808 62086 6820
rect 63678 6808 63684 6820
rect 63736 6808 63742 6860
rect 76926 6808 76932 6860
rect 76984 6848 76990 6860
rect 78858 6848 78864 6860
rect 76984 6820 78864 6848
rect 76984 6808 76990 6820
rect 78858 6808 78864 6820
rect 78916 6808 78922 6860
rect 92382 6808 92388 6860
rect 92440 6848 92446 6860
rect 94590 6848 94596 6860
rect 92440 6820 94596 6848
rect 92440 6808 92446 6820
rect 94590 6808 94596 6820
rect 94648 6808 94654 6860
rect 107562 6808 107568 6860
rect 107620 6848 107626 6860
rect 110046 6848 110052 6860
rect 107620 6820 110052 6848
rect 107620 6808 107626 6820
rect 110046 6808 110052 6820
rect 110104 6808 110110 6860
rect 122742 6808 122748 6860
rect 122800 6848 122806 6860
rect 125502 6848 125508 6860
rect 122800 6820 125508 6848
rect 122800 6808 122806 6820
rect 125502 6808 125508 6820
rect 125560 6808 125566 6860
rect 137922 6808 137928 6860
rect 137980 6848 137986 6860
rect 140682 6848 140688 6860
rect 137980 6820 140688 6848
rect 137980 6808 137986 6820
rect 140682 6808 140688 6820
rect 140740 6808 140746 6860
rect 153102 6808 153108 6860
rect 153160 6848 153166 6860
rect 155862 6848 155868 6860
rect 153160 6820 155868 6848
rect 153160 6808 153166 6820
rect 155862 6808 155868 6820
rect 155920 6808 155926 6860
rect 169662 6808 169668 6860
rect 169720 6848 169726 6860
rect 171594 6848 171600 6860
rect 169720 6820 171600 6848
rect 169720 6808 169726 6820
rect 171594 6808 171600 6820
rect 171652 6808 171658 6860
rect 184842 6808 184848 6860
rect 184900 6848 184906 6860
rect 187326 6848 187332 6860
rect 184900 6820 187332 6848
rect 184900 6808 184906 6820
rect 187326 6808 187332 6820
rect 187384 6808 187390 6860
rect 200022 6808 200028 6860
rect 200080 6848 200086 6860
rect 202782 6848 202788 6860
rect 200080 6820 202788 6848
rect 200080 6808 200086 6820
rect 202782 6808 202788 6820
rect 202840 6808 202846 6860
rect 215202 6808 215208 6860
rect 215260 6848 215266 6860
rect 218054 6848 218060 6860
rect 215260 6820 218060 6848
rect 215260 6808 215266 6820
rect 218054 6808 218060 6820
rect 218112 6808 218118 6860
rect 230382 6808 230388 6860
rect 230440 6848 230446 6860
rect 233050 6848 233056 6860
rect 230440 6820 233056 6848
rect 230440 6808 230446 6820
rect 233050 6808 233056 6820
rect 233108 6808 233114 6860
rect 245562 6808 245568 6860
rect 245620 6848 245626 6860
rect 249150 6848 249156 6860
rect 245620 6820 249156 6848
rect 245620 6808 245626 6820
rect 249150 6808 249156 6820
rect 249208 6808 249214 6860
rect 260466 6808 260472 6860
rect 260524 6848 260530 6860
rect 264330 6848 264336 6860
rect 260524 6820 264336 6848
rect 260524 6808 260530 6820
rect 264330 6808 264336 6820
rect 264388 6808 264394 6860
rect 275922 6808 275928 6860
rect 275980 6848 275986 6860
rect 280062 6848 280068 6860
rect 275980 6820 280068 6848
rect 275980 6808 275986 6820
rect 280062 6808 280068 6820
rect 280120 6808 280126 6860
rect 291102 6808 291108 6860
rect 291160 6848 291166 6860
rect 295518 6848 295524 6860
rect 291160 6820 295524 6848
rect 291160 6808 291166 6820
rect 295518 6808 295524 6820
rect 295576 6808 295582 6860
rect 321462 6808 321468 6860
rect 321520 6848 321526 6860
rect 326430 6848 326436 6860
rect 321520 6820 326436 6848
rect 321520 6808 321526 6820
rect 326430 6808 326436 6820
rect 326488 6808 326494 6860
rect 336826 6808 336832 6860
rect 336884 6848 336890 6860
rect 341886 6848 341892 6860
rect 336884 6820 341892 6848
rect 336884 6808 336890 6820
rect 341886 6808 341892 6820
rect 341944 6808 341950 6860
rect 353202 6808 353208 6860
rect 353260 6848 353266 6860
rect 357066 6848 357072 6860
rect 353260 6820 357072 6848
rect 353260 6808 353266 6820
rect 357066 6808 357072 6820
rect 357124 6808 357130 6860
rect 368382 6808 368388 6860
rect 368440 6848 368446 6860
rect 372798 6848 372804 6860
rect 368440 6820 372804 6848
rect 368440 6808 368446 6820
rect 372798 6808 372804 6820
rect 372856 6808 372862 6860
rect 398742 6808 398748 6860
rect 398800 6848 398806 6860
rect 403434 6848 403440 6860
rect 398800 6820 403440 6848
rect 398800 6808 398806 6820
rect 403434 6808 403440 6820
rect 403492 6808 403498 6860
rect 413922 6808 413928 6860
rect 413980 6848 413986 6860
rect 419166 6848 419172 6860
rect 413980 6820 419172 6848
rect 413980 6808 413986 6820
rect 419166 6808 419172 6820
rect 419224 6808 419230 6860
rect 429102 6808 429108 6860
rect 429160 6848 429166 6860
rect 434622 6848 434628 6860
rect 429160 6820 434628 6848
rect 429160 6808 429166 6820
rect 434622 6808 434628 6820
rect 434680 6808 434686 6860
rect 444098 6808 444104 6860
rect 444156 6848 444162 6860
rect 449894 6848 449900 6860
rect 444156 6820 449900 6848
rect 444156 6808 444162 6820
rect 449894 6808 449900 6820
rect 449952 6808 449958 6860
rect 474642 6808 474648 6860
rect 474700 6848 474706 6860
rect 478874 6848 478880 6860
rect 474700 6820 478880 6848
rect 474700 6808 474706 6820
rect 478874 6808 478880 6820
rect 478932 6808 478938 6860
rect 505002 6808 505008 6860
rect 505060 6848 505066 6860
rect 510522 6848 510528 6860
rect 505060 6820 510528 6848
rect 505060 6808 505066 6820
rect 510522 6808 510528 6820
rect 510580 6808 510586 6860
rect 520918 6808 520924 6860
rect 520976 6848 520982 6860
rect 527082 6848 527088 6860
rect 520976 6820 527088 6848
rect 520976 6808 520982 6820
rect 527082 6808 527088 6820
rect 527140 6808 527146 6860
rect 551922 6808 551928 6860
rect 551980 6848 551986 6860
rect 556154 6848 556160 6860
rect 551980 6820 556160 6848
rect 551980 6808 551986 6820
rect 556154 6808 556160 6820
rect 556212 6808 556218 6860
rect 582282 6808 582288 6860
rect 582340 6848 582346 6860
rect 588906 6848 588912 6860
rect 582340 6820 588912 6848
rect 582340 6808 582346 6820
rect 588906 6808 588912 6820
rect 588964 6808 588970 6860
rect 597278 6808 597284 6860
rect 597336 6848 597342 6860
rect 604638 6848 604644 6860
rect 597336 6820 604644 6848
rect 597336 6808 597342 6820
rect 604638 6808 604644 6820
rect 604696 6808 604702 6860
rect 658182 6808 658188 6860
rect 658240 6848 658246 6860
rect 666462 6848 666468 6860
rect 658240 6820 666468 6848
rect 658240 6808 658246 6820
rect 666462 6808 666468 6820
rect 666520 6808 666526 6860
rect 1104 6554 682824 6576
rect 1104 6502 86825 6554
rect 86877 6502 86889 6554
rect 86941 6502 86953 6554
rect 87005 6502 87017 6554
rect 87069 6502 87081 6554
rect 87133 6502 257255 6554
rect 257307 6502 257319 6554
rect 257371 6502 257383 6554
rect 257435 6502 257447 6554
rect 257499 6502 257511 6554
rect 257563 6502 427685 6554
rect 427737 6502 427749 6554
rect 427801 6502 427813 6554
rect 427865 6502 427877 6554
rect 427929 6502 427941 6554
rect 427993 6502 598115 6554
rect 598167 6502 598179 6554
rect 598231 6502 598243 6554
rect 598295 6502 598307 6554
rect 598359 6502 598371 6554
rect 598423 6502 682824 6554
rect 1104 6480 682824 6502
rect 306282 6128 306288 6180
rect 306340 6168 306346 6180
rect 310698 6168 310704 6180
rect 306340 6140 310704 6168
rect 306340 6128 306346 6140
rect 310698 6128 310704 6140
rect 310756 6128 310762 6180
rect 383562 6128 383568 6180
rect 383620 6168 383626 6180
rect 388254 6168 388260 6180
rect 383620 6140 388260 6168
rect 383620 6128 383626 6140
rect 388254 6128 388260 6140
rect 388312 6128 388318 6180
rect 459462 6128 459468 6180
rect 459520 6168 459526 6180
rect 464982 6168 464988 6180
rect 459520 6140 464988 6168
rect 459520 6128 459526 6140
rect 464982 6128 464988 6140
rect 465040 6128 465046 6180
rect 489822 6128 489828 6180
rect 489880 6168 489886 6180
rect 496170 6168 496176 6180
rect 489880 6140 496176 6168
rect 489880 6128 489886 6140
rect 496170 6128 496176 6140
rect 496228 6128 496234 6180
rect 536742 6128 536748 6180
rect 536800 6168 536806 6180
rect 542262 6168 542268 6180
rect 536800 6140 542268 6168
rect 536800 6128 536806 6140
rect 542262 6128 542268 6140
rect 542320 6128 542326 6180
rect 567102 6128 567108 6180
rect 567160 6168 567166 6180
rect 572622 6168 572628 6180
rect 567160 6140 572628 6168
rect 567160 6128 567166 6140
rect 572622 6128 572628 6140
rect 572680 6128 572686 6180
rect 612642 6128 612648 6180
rect 612700 6168 612706 6180
rect 620094 6168 620100 6180
rect 612700 6140 620100 6168
rect 612700 6128 612706 6140
rect 620094 6128 620100 6140
rect 620152 6128 620158 6180
rect 627638 6128 627644 6180
rect 627696 6168 627702 6180
rect 635550 6168 635556 6180
rect 627696 6140 635556 6168
rect 627696 6128 627702 6140
rect 635550 6128 635556 6140
rect 635608 6128 635614 6180
rect 643002 6128 643008 6180
rect 643060 6168 643066 6180
rect 651006 6168 651012 6180
rect 643060 6140 651012 6168
rect 643060 6128 643066 6140
rect 651006 6128 651012 6140
rect 651064 6128 651070 6180
rect 673362 6128 673368 6180
rect 673420 6168 673426 6180
rect 681734 6168 681740 6180
rect 673420 6140 681740 6168
rect 673420 6128 673426 6140
rect 681734 6128 681740 6140
rect 681792 6128 681798 6180
rect 1104 6010 682824 6032
rect 1104 5958 86165 6010
rect 86217 5958 86229 6010
rect 86281 5958 86293 6010
rect 86345 5958 86357 6010
rect 86409 5958 86421 6010
rect 86473 5958 256595 6010
rect 256647 5958 256659 6010
rect 256711 5958 256723 6010
rect 256775 5958 256787 6010
rect 256839 5958 256851 6010
rect 256903 5958 427025 6010
rect 427077 5958 427089 6010
rect 427141 5958 427153 6010
rect 427205 5958 427217 6010
rect 427269 5958 427281 6010
rect 427333 5958 597455 6010
rect 597507 5958 597519 6010
rect 597571 5958 597583 6010
rect 597635 5958 597647 6010
rect 597699 5958 597711 6010
rect 597763 5958 682824 6010
rect 1104 5936 682824 5958
rect 1104 5466 682824 5488
rect 1104 5414 86825 5466
rect 86877 5414 86889 5466
rect 86941 5414 86953 5466
rect 87005 5414 87017 5466
rect 87069 5414 87081 5466
rect 87133 5414 257255 5466
rect 257307 5414 257319 5466
rect 257371 5414 257383 5466
rect 257435 5414 257447 5466
rect 257499 5414 257511 5466
rect 257563 5414 427685 5466
rect 427737 5414 427749 5466
rect 427801 5414 427813 5466
rect 427865 5414 427877 5466
rect 427929 5414 427941 5466
rect 427993 5414 598115 5466
rect 598167 5414 598179 5466
rect 598231 5414 598243 5466
rect 598295 5414 598307 5466
rect 598359 5414 598371 5466
rect 598423 5414 682824 5466
rect 1104 5392 682824 5414
rect 1104 4922 682824 4944
rect 1104 4870 86165 4922
rect 86217 4870 86229 4922
rect 86281 4870 86293 4922
rect 86345 4870 86357 4922
rect 86409 4870 86421 4922
rect 86473 4870 256595 4922
rect 256647 4870 256659 4922
rect 256711 4870 256723 4922
rect 256775 4870 256787 4922
rect 256839 4870 256851 4922
rect 256903 4870 427025 4922
rect 427077 4870 427089 4922
rect 427141 4870 427153 4922
rect 427205 4870 427217 4922
rect 427269 4870 427281 4922
rect 427333 4870 597455 4922
rect 597507 4870 597519 4922
rect 597571 4870 597583 4922
rect 597635 4870 597647 4922
rect 597699 4870 597711 4922
rect 597763 4870 682824 4922
rect 1104 4848 682824 4870
rect 1104 4378 682824 4400
rect 1104 4326 86825 4378
rect 86877 4326 86889 4378
rect 86941 4326 86953 4378
rect 87005 4326 87017 4378
rect 87069 4326 87081 4378
rect 87133 4326 257255 4378
rect 257307 4326 257319 4378
rect 257371 4326 257383 4378
rect 257435 4326 257447 4378
rect 257499 4326 257511 4378
rect 257563 4326 427685 4378
rect 427737 4326 427749 4378
rect 427801 4326 427813 4378
rect 427865 4326 427877 4378
rect 427929 4326 427941 4378
rect 427993 4326 598115 4378
rect 598167 4326 598179 4378
rect 598231 4326 598243 4378
rect 598295 4326 598307 4378
rect 598359 4326 598371 4378
rect 598423 4326 682824 4378
rect 1104 4304 682824 4326
rect 1104 3834 682824 3856
rect 1104 3782 86165 3834
rect 86217 3782 86229 3834
rect 86281 3782 86293 3834
rect 86345 3782 86357 3834
rect 86409 3782 86421 3834
rect 86473 3782 256595 3834
rect 256647 3782 256659 3834
rect 256711 3782 256723 3834
rect 256775 3782 256787 3834
rect 256839 3782 256851 3834
rect 256903 3782 427025 3834
rect 427077 3782 427089 3834
rect 427141 3782 427153 3834
rect 427205 3782 427217 3834
rect 427269 3782 427281 3834
rect 427333 3782 597455 3834
rect 597507 3782 597519 3834
rect 597571 3782 597583 3834
rect 597635 3782 597647 3834
rect 597699 3782 597711 3834
rect 597763 3782 682824 3834
rect 1104 3760 682824 3782
rect 339586 3476 339592 3528
rect 339644 3516 339650 3528
rect 432693 3519 432751 3525
rect 432693 3516 432705 3519
rect 339644 3488 432705 3516
rect 339644 3476 339650 3488
rect 432693 3485 432705 3488
rect 432739 3516 432751 3519
rect 432966 3516 432972 3528
rect 432739 3488 432972 3516
rect 432739 3485 432751 3488
rect 432693 3479 432751 3485
rect 432966 3476 432972 3488
rect 433024 3476 433030 3528
rect 433426 3476 433432 3528
rect 433484 3516 433490 3528
rect 433889 3519 433947 3525
rect 433889 3516 433901 3519
rect 433484 3488 433901 3516
rect 433484 3476 433490 3488
rect 433889 3485 433901 3488
rect 433935 3516 433947 3519
rect 526990 3516 526996 3528
rect 433935 3488 526996 3516
rect 433935 3485 433947 3488
rect 433889 3479 433947 3485
rect 526990 3476 526996 3488
rect 527048 3476 527054 3528
rect 337378 3408 337384 3460
rect 337436 3448 337442 3460
rect 337657 3451 337715 3457
rect 337657 3448 337669 3451
rect 337436 3420 337669 3448
rect 337436 3408 337442 3420
rect 337657 3417 337669 3420
rect 337703 3448 337715 3451
rect 431678 3448 431684 3460
rect 337703 3420 431684 3448
rect 337703 3417 337715 3420
rect 337657 3411 337715 3417
rect 431678 3408 431684 3420
rect 431736 3408 431742 3460
rect 433518 3408 433524 3460
rect 433576 3448 433582 3460
rect 527177 3451 527235 3457
rect 527177 3448 527189 3451
rect 433576 3420 527189 3448
rect 433576 3408 433582 3420
rect 527177 3417 527189 3420
rect 527223 3448 527235 3451
rect 527542 3448 527548 3460
rect 527223 3420 527548 3448
rect 527223 3417 527235 3420
rect 527177 3411 527235 3417
rect 527542 3408 527548 3420
rect 527600 3408 527606 3460
rect 248414 3340 248420 3392
rect 248472 3380 248478 3392
rect 248693 3383 248751 3389
rect 248693 3380 248705 3383
rect 248472 3352 248705 3380
rect 248472 3340 248478 3352
rect 248693 3349 248705 3352
rect 248739 3349 248751 3383
rect 248693 3343 248751 3349
rect 336277 3383 336335 3389
rect 336277 3349 336289 3383
rect 336323 3380 336335 3383
rect 336458 3380 336464 3392
rect 336323 3352 336464 3380
rect 336323 3349 336335 3352
rect 336277 3343 336335 3349
rect 336458 3340 336464 3352
rect 336516 3340 336522 3392
rect 338206 3340 338212 3392
rect 338264 3380 338270 3392
rect 338853 3383 338911 3389
rect 338853 3380 338865 3383
rect 338264 3352 338865 3380
rect 338264 3340 338270 3352
rect 338853 3349 338865 3352
rect 338899 3349 338911 3383
rect 338853 3343 338911 3349
rect 339862 3340 339868 3392
rect 339920 3380 339926 3392
rect 426894 3380 426900 3392
rect 339920 3352 426900 3380
rect 339920 3340 339926 3352
rect 426894 3340 426900 3352
rect 426952 3340 426958 3392
rect 433334 3340 433340 3392
rect 433392 3340 433398 3392
rect 434441 3383 434499 3389
rect 434441 3349 434453 3383
rect 434487 3380 434499 3383
rect 434530 3380 434536 3392
rect 434487 3352 434536 3380
rect 434487 3349 434499 3352
rect 434441 3343 434499 3349
rect 434530 3340 434536 3352
rect 434588 3340 434594 3392
rect 1104 3290 682824 3312
rect 1104 3238 86825 3290
rect 86877 3238 86889 3290
rect 86941 3238 86953 3290
rect 87005 3238 87017 3290
rect 87069 3238 87081 3290
rect 87133 3238 257255 3290
rect 257307 3238 257319 3290
rect 257371 3238 257383 3290
rect 257435 3238 257447 3290
rect 257499 3238 257511 3290
rect 257563 3238 427685 3290
rect 427737 3238 427749 3290
rect 427801 3238 427813 3290
rect 427865 3238 427877 3290
rect 427929 3238 427941 3290
rect 427993 3238 598115 3290
rect 598167 3238 598179 3290
rect 598231 3238 598243 3290
rect 598295 3238 598307 3290
rect 598359 3238 598371 3290
rect 598423 3238 682824 3290
rect 1104 3216 682824 3238
rect 78858 3136 78864 3188
rect 78916 3136 78922 3188
rect 171594 3136 171600 3188
rect 171652 3136 171658 3188
rect 218054 3136 218060 3188
rect 218112 3136 218118 3188
rect 242158 3136 242164 3188
rect 242216 3176 242222 3188
rect 338393 3179 338451 3185
rect 338393 3176 338405 3179
rect 242216 3148 338405 3176
rect 242216 3136 242222 3148
rect 338393 3145 338405 3148
rect 338439 3145 338451 3179
rect 338393 3139 338451 3145
rect 247034 3068 247040 3120
rect 247092 3108 247098 3120
rect 278961 3111 279019 3117
rect 278961 3108 278973 3111
rect 247092 3080 278973 3108
rect 247092 3068 247098 3080
rect 278961 3077 278973 3080
rect 279007 3108 279019 3111
rect 295705 3111 295763 3117
rect 279007 3080 279648 3108
rect 279007 3077 279019 3080
rect 278961 3071 279019 3077
rect 248414 3000 248420 3052
rect 248472 3040 248478 3052
rect 248969 3043 249027 3049
rect 248969 3040 248981 3043
rect 248472 3012 248981 3040
rect 248472 3000 248478 3012
rect 248969 3009 248981 3012
rect 249015 3009 249027 3043
rect 248969 3003 249027 3009
rect 264330 3000 264336 3052
rect 264388 3000 264394 3052
rect 279620 3049 279648 3080
rect 279804 3080 287054 3108
rect 279605 3043 279663 3049
rect 279605 3009 279617 3043
rect 279651 3009 279663 3043
rect 279605 3003 279663 3009
rect 249702 2932 249708 2984
rect 249760 2972 249766 2984
rect 279804 2972 279832 3080
rect 279881 3043 279939 3049
rect 279881 3009 279893 3043
rect 279927 3040 279939 3043
rect 279927 3012 283420 3040
rect 279927 3009 279939 3012
rect 279881 3003 279939 3009
rect 249760 2944 279832 2972
rect 249760 2932 249766 2944
rect 283392 2904 283420 3012
rect 287026 2972 287054 3080
rect 295705 3077 295717 3111
rect 295751 3108 295763 3111
rect 295751 3080 338344 3108
rect 295751 3077 295763 3080
rect 295705 3071 295763 3077
rect 295153 3043 295211 3049
rect 295153 3040 295165 3043
rect 294432 3012 295165 3040
rect 294432 2981 294460 3012
rect 295153 3009 295165 3012
rect 295199 3009 295211 3043
rect 295153 3003 295211 3009
rect 310698 3000 310704 3052
rect 310756 3000 310762 3052
rect 337378 3000 337384 3052
rect 337436 3000 337442 3052
rect 294417 2975 294475 2981
rect 294417 2972 294429 2975
rect 287026 2944 294429 2972
rect 294417 2941 294429 2944
rect 294463 2941 294475 2975
rect 294417 2935 294475 2941
rect 336826 2932 336832 2984
rect 336884 2932 336890 2984
rect 338316 2972 338344 3080
rect 338408 3040 338436 3139
rect 357066 3136 357072 3188
rect 357124 3136 357130 3188
rect 403434 3136 403440 3188
rect 403492 3136 403498 3188
rect 426894 3136 426900 3188
rect 426952 3176 426958 3188
rect 426952 3148 431954 3176
rect 426952 3136 426958 3148
rect 387981 3111 388039 3117
rect 387981 3108 387993 3111
rect 339144 3080 387993 3108
rect 339037 3043 339095 3049
rect 339037 3040 339049 3043
rect 338408 3012 339049 3040
rect 339037 3009 339049 3012
rect 339083 3009 339095 3043
rect 339037 3003 339095 3009
rect 339144 2972 339172 3080
rect 387981 3077 387993 3080
rect 388027 3108 388039 3111
rect 388438 3108 388444 3120
rect 388027 3080 388444 3108
rect 388027 3077 388039 3080
rect 387981 3071 388039 3077
rect 388438 3068 388444 3080
rect 388496 3068 388502 3120
rect 431926 3108 431954 3148
rect 433334 3136 433340 3188
rect 433392 3176 433398 3188
rect 433392 3148 525656 3176
rect 433392 3136 433398 3148
rect 434257 3111 434315 3117
rect 434257 3108 434269 3111
rect 431926 3080 434269 3108
rect 434257 3077 434269 3080
rect 434303 3077 434315 3111
rect 434257 3071 434315 3077
rect 449894 3068 449900 3120
rect 449952 3068 449958 3120
rect 496170 3068 496176 3120
rect 496228 3068 496234 3120
rect 525628 3117 525656 3148
rect 588906 3136 588912 3188
rect 588964 3136 588970 3188
rect 681734 3136 681740 3188
rect 681792 3136 681798 3188
rect 525613 3111 525671 3117
rect 525613 3077 525625 3111
rect 525659 3077 525671 3111
rect 525613 3071 525671 3077
rect 525904 3080 528554 3108
rect 339586 3000 339592 3052
rect 339644 3000 339650 3052
rect 342073 3043 342131 3049
rect 342073 3009 342085 3043
rect 342119 3040 342131 3043
rect 342714 3040 342720 3052
rect 342119 3012 342720 3040
rect 342119 3009 342131 3012
rect 342073 3003 342131 3009
rect 342714 3000 342720 3012
rect 342772 3000 342778 3052
rect 430758 3000 430764 3052
rect 430816 3040 430822 3052
rect 431405 3043 431463 3049
rect 431405 3040 431417 3043
rect 430816 3012 431417 3040
rect 430816 3000 430822 3012
rect 431405 3009 431417 3012
rect 431451 3009 431463 3043
rect 431405 3003 431463 3009
rect 432966 3000 432972 3052
rect 433024 3000 433030 3052
rect 433518 3000 433524 3052
rect 433576 3000 433582 3052
rect 434809 3043 434867 3049
rect 434809 3009 434821 3043
rect 434855 3040 434867 3043
rect 435450 3040 435456 3052
rect 434855 3012 435456 3040
rect 434855 3009 434867 3012
rect 434809 3003 434867 3009
rect 435450 3000 435456 3012
rect 435508 3000 435514 3052
rect 463234 3000 463240 3052
rect 463292 3040 463298 3052
rect 463881 3043 463939 3049
rect 463881 3040 463893 3043
rect 463292 3012 463893 3040
rect 463292 3000 463298 3012
rect 463881 3009 463893 3012
rect 463927 3009 463939 3043
rect 463881 3003 463939 3009
rect 478690 3000 478696 3052
rect 478748 3040 478754 3052
rect 525904 3049 525932 3080
rect 479337 3043 479395 3049
rect 479337 3040 479349 3043
rect 478748 3012 479349 3040
rect 478748 3000 478754 3012
rect 479337 3009 479349 3012
rect 479383 3009 479395 3043
rect 479337 3003 479395 3009
rect 525889 3043 525947 3049
rect 525889 3009 525901 3043
rect 525935 3009 525947 3043
rect 527545 3043 527603 3049
rect 525889 3003 525947 3009
rect 525996 3012 527128 3040
rect 338316 2944 339172 2972
rect 341518 2932 341524 2984
rect 341576 2932 341582 2984
rect 431862 2932 431868 2984
rect 431920 2932 431926 2984
rect 464433 2975 464491 2981
rect 464433 2941 464445 2975
rect 464479 2972 464491 2975
rect 479889 2975 479947 2981
rect 464479 2944 470594 2972
rect 464479 2941 464491 2944
rect 464433 2935 464491 2941
rect 372617 2907 372675 2913
rect 372617 2904 372629 2907
rect 283392 2876 372629 2904
rect 372617 2873 372629 2876
rect 372663 2904 372675 2907
rect 372982 2904 372988 2916
rect 372663 2876 372988 2904
rect 372663 2873 372675 2876
rect 372617 2867 372675 2873
rect 372982 2864 372988 2876
rect 373040 2864 373046 2916
rect 470566 2904 470594 2944
rect 479889 2941 479901 2975
rect 479935 2972 479947 2975
rect 525996 2972 526024 3012
rect 479935 2944 526024 2972
rect 479935 2941 479947 2944
rect 479889 2935 479947 2941
rect 526990 2932 526996 2984
rect 527048 2932 527054 2984
rect 527100 2972 527128 3012
rect 527545 3009 527557 3043
rect 527591 3040 527603 3043
rect 528186 3040 528192 3052
rect 527591 3012 528192 3040
rect 527591 3009 527603 3012
rect 527545 3003 527603 3009
rect 528186 3000 528192 3012
rect 528244 3000 528250 3052
rect 528526 3040 528554 3080
rect 539502 3040 539508 3052
rect 528526 3012 539508 3040
rect 539502 3000 539508 3012
rect 539560 3000 539566 3052
rect 573453 2975 573511 2981
rect 573453 2972 573465 2975
rect 527100 2944 573465 2972
rect 573453 2941 573465 2944
rect 573499 2972 573511 2975
rect 573910 2972 573916 2984
rect 573499 2944 573916 2972
rect 573499 2941 573511 2944
rect 573453 2935 573511 2941
rect 573910 2932 573916 2944
rect 573968 2932 573974 2984
rect 470566 2876 547874 2904
rect 136453 2839 136511 2845
rect 136453 2805 136465 2839
rect 136499 2836 136511 2839
rect 136542 2836 136548 2848
rect 136499 2808 136548 2836
rect 136499 2805 136511 2808
rect 136453 2799 136511 2805
rect 136542 2796 136548 2808
rect 136600 2796 136606 2848
rect 187694 2796 187700 2848
rect 187752 2796 187758 2848
rect 202966 2796 202972 2848
rect 203024 2836 203030 2848
rect 203061 2839 203119 2845
rect 203061 2836 203073 2839
rect 203024 2808 203073 2836
rect 203024 2796 203030 2808
rect 203061 2805 203073 2808
rect 203107 2805 203119 2839
rect 203061 2799 203119 2805
rect 249242 2796 249248 2848
rect 249300 2796 249306 2848
rect 277210 2796 277216 2848
rect 277268 2796 277274 2848
rect 292669 2839 292727 2845
rect 292669 2805 292681 2839
rect 292715 2836 292727 2839
rect 292850 2836 292856 2848
rect 292715 2808 292856 2836
rect 292715 2805 292727 2808
rect 292669 2799 292727 2805
rect 292850 2796 292856 2808
rect 292908 2796 292914 2848
rect 323397 2839 323455 2845
rect 323397 2805 323409 2839
rect 323443 2836 323455 2839
rect 323578 2836 323584 2848
rect 323443 2808 323584 2836
rect 323443 2805 323455 2808
rect 323397 2799 323455 2805
rect 323578 2796 323584 2808
rect 323636 2796 323642 2848
rect 324498 2796 324504 2848
rect 324556 2796 324562 2848
rect 326154 2796 326160 2848
rect 326212 2796 326218 2848
rect 331582 2796 331588 2848
rect 331640 2836 331646 2848
rect 331677 2839 331735 2845
rect 331677 2836 331689 2839
rect 331640 2808 331689 2836
rect 331640 2796 331646 2808
rect 331677 2805 331689 2808
rect 331723 2805 331735 2839
rect 331677 2799 331735 2805
rect 333054 2796 333060 2848
rect 333112 2836 333118 2848
rect 333241 2839 333299 2845
rect 333241 2836 333253 2839
rect 333112 2808 333253 2836
rect 333112 2796 333118 2808
rect 333241 2805 333253 2808
rect 333287 2805 333299 2839
rect 333241 2799 333299 2805
rect 334618 2796 334624 2848
rect 334676 2836 334682 2848
rect 334805 2839 334863 2845
rect 334805 2836 334817 2839
rect 334676 2808 334817 2836
rect 334676 2796 334682 2808
rect 334805 2805 334817 2808
rect 334851 2805 334863 2839
rect 334805 2799 334863 2805
rect 335722 2796 335728 2848
rect 335780 2796 335786 2848
rect 340230 2796 340236 2848
rect 340288 2796 340294 2848
rect 342714 2796 342720 2848
rect 342772 2796 342778 2848
rect 367462 2796 367468 2848
rect 367520 2796 367526 2848
rect 370866 2796 370872 2848
rect 370924 2796 370930 2848
rect 382826 2796 382832 2848
rect 382884 2796 382890 2848
rect 386417 2839 386475 2845
rect 386417 2805 386429 2839
rect 386463 2836 386475 2839
rect 386598 2836 386604 2848
rect 386463 2808 386604 2836
rect 386463 2805 386475 2808
rect 386417 2799 386475 2805
rect 386598 2796 386604 2808
rect 386656 2796 386662 2848
rect 417329 2839 417387 2845
rect 417329 2805 417341 2839
rect 417375 2836 417387 2839
rect 417510 2836 417516 2848
rect 417375 2808 417516 2836
rect 417375 2805 417387 2808
rect 417329 2799 417387 2805
rect 417510 2796 417516 2808
rect 417568 2796 417574 2848
rect 418890 2796 418896 2848
rect 418948 2796 418954 2848
rect 430758 2796 430764 2848
rect 430816 2796 430822 2848
rect 435450 2796 435456 2848
rect 435508 2796 435514 2848
rect 463234 2796 463240 2848
rect 463292 2796 463298 2848
rect 465258 2796 465264 2848
rect 465316 2796 465322 2848
rect 478690 2796 478696 2848
rect 478748 2796 478754 2848
rect 480714 2796 480720 2848
rect 480772 2796 480778 2848
rect 511626 2796 511632 2848
rect 511684 2796 511690 2848
rect 528186 2796 528192 2848
rect 528244 2796 528250 2848
rect 528830 2796 528836 2848
rect 528888 2836 528894 2848
rect 529017 2839 529075 2845
rect 529017 2836 529029 2839
rect 528888 2808 529029 2836
rect 528888 2796 528894 2808
rect 529017 2805 529029 2808
rect 529063 2805 529075 2839
rect 547846 2836 547874 2876
rect 558086 2836 558092 2848
rect 547846 2808 558092 2836
rect 529017 2799 529075 2805
rect 558086 2796 558092 2808
rect 558144 2796 558150 2848
rect 604454 2796 604460 2848
rect 604512 2796 604518 2848
rect 619818 2796 619824 2848
rect 619876 2796 619882 2848
rect 650730 2796 650736 2848
rect 650788 2796 650794 2848
rect 666186 2796 666192 2848
rect 666244 2796 666250 2848
rect 1104 2746 682824 2768
rect 1104 2694 86165 2746
rect 86217 2694 86229 2746
rect 86281 2694 86293 2746
rect 86345 2694 86357 2746
rect 86409 2694 86421 2746
rect 86473 2694 256595 2746
rect 256647 2694 256659 2746
rect 256711 2694 256723 2746
rect 256775 2694 256787 2746
rect 256839 2694 256851 2746
rect 256903 2694 427025 2746
rect 427077 2694 427089 2746
rect 427141 2694 427153 2746
rect 427205 2694 427217 2746
rect 427269 2694 427281 2746
rect 427333 2694 597455 2746
rect 597507 2694 597519 2746
rect 597571 2694 597583 2746
rect 597635 2694 597647 2746
rect 597699 2694 597711 2746
rect 597763 2694 682824 2746
rect 1104 2672 682824 2694
rect 1854 2592 1860 2644
rect 1912 2592 1918 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 17313 2635 17371 2641
rect 17313 2632 17325 2635
rect 16632 2604 17325 2632
rect 16632 2592 16638 2604
rect 17313 2601 17325 2604
rect 17359 2601 17371 2635
rect 17313 2595 17371 2601
rect 46934 2592 46940 2644
rect 46992 2632 46998 2644
rect 48225 2635 48283 2641
rect 48225 2632 48237 2635
rect 46992 2604 48237 2632
rect 46992 2592 46998 2604
rect 48225 2601 48237 2604
rect 48271 2601 48283 2635
rect 48225 2595 48283 2601
rect 63678 2592 63684 2644
rect 63736 2592 63742 2644
rect 94590 2592 94596 2644
rect 94648 2592 94654 2644
rect 97350 2592 97356 2644
rect 97408 2632 97414 2644
rect 97997 2635 98055 2641
rect 97997 2632 98009 2635
rect 97408 2604 98009 2632
rect 97408 2592 97414 2604
rect 97997 2601 98009 2604
rect 98043 2632 98055 2635
rect 98043 2604 180794 2632
rect 98043 2601 98055 2604
rect 97997 2595 98055 2601
rect 32953 2567 33011 2573
rect 32953 2533 32965 2567
rect 32999 2564 33011 2567
rect 48961 2567 49019 2573
rect 48961 2564 48973 2567
rect 32999 2536 35894 2564
rect 32999 2533 33011 2536
rect 32953 2527 33011 2533
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 17497 2431 17555 2437
rect 2087 2400 2636 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2608 2304 2636 2400
rect 17497 2397 17509 2431
rect 17543 2428 17555 2431
rect 17543 2400 18092 2428
rect 17543 2397 17555 2400
rect 17497 2391 17555 2397
rect 18064 2304 18092 2400
rect 31754 2388 31760 2440
rect 31812 2428 31818 2440
rect 32769 2431 32827 2437
rect 32769 2428 32781 2431
rect 31812 2400 32781 2428
rect 31812 2388 31818 2400
rect 32769 2397 32781 2400
rect 32815 2428 32827 2431
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 32815 2400 33425 2428
rect 32815 2397 32827 2400
rect 32769 2391 32827 2397
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 35866 2428 35894 2536
rect 48424 2536 48973 2564
rect 41049 2499 41107 2505
rect 41049 2465 41061 2499
rect 41095 2496 41107 2499
rect 41095 2468 45554 2496
rect 41095 2465 41107 2468
rect 41049 2459 41107 2465
rect 40773 2431 40831 2437
rect 40773 2428 40785 2431
rect 35866 2400 40785 2428
rect 33413 2391 33471 2397
rect 40773 2397 40785 2400
rect 40819 2397 40831 2431
rect 40773 2391 40831 2397
rect 45526 2360 45554 2468
rect 48424 2437 48452 2536
rect 48961 2533 48973 2536
rect 49007 2564 49019 2567
rect 49007 2536 136956 2564
rect 49007 2533 49019 2536
rect 48961 2527 49019 2533
rect 134705 2499 134763 2505
rect 134705 2496 134717 2499
rect 55186 2468 134717 2496
rect 48409 2431 48467 2437
rect 48409 2397 48421 2431
rect 48455 2397 48467 2431
rect 48409 2391 48467 2397
rect 55186 2360 55214 2468
rect 134705 2465 134717 2468
rect 134751 2465 134763 2499
rect 134705 2459 134763 2465
rect 63865 2431 63923 2437
rect 63865 2397 63877 2431
rect 63911 2428 63923 2431
rect 63911 2400 64460 2428
rect 63911 2397 63923 2400
rect 63865 2391 63923 2397
rect 64432 2369 64460 2400
rect 78858 2388 78864 2440
rect 78916 2428 78922 2440
rect 79321 2431 79379 2437
rect 79321 2428 79333 2431
rect 78916 2400 79333 2428
rect 78916 2388 78922 2400
rect 79321 2397 79333 2400
rect 79367 2397 79379 2431
rect 79321 2391 79379 2397
rect 94777 2431 94835 2437
rect 94777 2397 94789 2431
rect 94823 2428 94835 2431
rect 95326 2428 95332 2440
rect 94823 2400 95332 2428
rect 94823 2397 94835 2400
rect 94777 2391 94835 2397
rect 95326 2388 95332 2400
rect 95384 2388 95390 2440
rect 96724 2400 96936 2428
rect 45526 2332 55214 2360
rect 64417 2363 64475 2369
rect 64417 2329 64429 2363
rect 64463 2360 64475 2363
rect 96724 2360 96752 2400
rect 64463 2332 96752 2360
rect 64463 2329 64475 2332
rect 64417 2323 64475 2329
rect 96798 2320 96804 2372
rect 96856 2320 96862 2372
rect 96908 2360 96936 2400
rect 97350 2388 97356 2440
rect 97408 2388 97414 2440
rect 110233 2431 110291 2437
rect 110233 2397 110245 2431
rect 110279 2428 110291 2431
rect 110690 2428 110696 2440
rect 110279 2400 110696 2428
rect 110279 2397 110291 2400
rect 110233 2391 110291 2397
rect 110690 2388 110696 2400
rect 110748 2388 110754 2440
rect 112809 2431 112867 2437
rect 112809 2397 112821 2431
rect 112855 2428 112867 2431
rect 113450 2428 113456 2440
rect 112855 2400 113456 2428
rect 112855 2397 112867 2400
rect 112809 2391 112867 2397
rect 113450 2388 113456 2400
rect 113508 2388 113514 2440
rect 125502 2388 125508 2440
rect 125560 2428 125566 2440
rect 126149 2431 126207 2437
rect 126149 2428 126161 2431
rect 125560 2400 126161 2428
rect 125560 2388 125566 2400
rect 126149 2397 126161 2400
rect 126195 2397 126207 2431
rect 134720 2428 134748 2459
rect 135441 2431 135499 2437
rect 135441 2428 135453 2431
rect 134720 2400 135453 2428
rect 126149 2391 126207 2397
rect 135441 2397 135453 2400
rect 135487 2397 135499 2431
rect 135441 2391 135499 2397
rect 136542 2388 136548 2440
rect 136600 2388 136606 2440
rect 96908 2332 110828 2360
rect 2590 2252 2596 2304
rect 2648 2252 2654 2304
rect 18046 2252 18052 2304
rect 18104 2252 18110 2304
rect 79134 2252 79140 2304
rect 79192 2252 79198 2304
rect 95326 2252 95332 2304
rect 95384 2252 95390 2304
rect 110046 2252 110052 2304
rect 110104 2252 110110 2304
rect 110690 2252 110696 2304
rect 110748 2252 110754 2304
rect 110800 2292 110828 2332
rect 112254 2320 112260 2372
rect 112312 2320 112318 2372
rect 113146 2332 128354 2360
rect 113146 2292 113174 2332
rect 110800 2264 113174 2292
rect 113450 2252 113456 2304
rect 113508 2252 113514 2304
rect 125686 2252 125692 2304
rect 125744 2252 125750 2304
rect 128326 2292 128354 2332
rect 135990 2320 135996 2372
rect 136048 2320 136054 2372
rect 136818 2320 136824 2372
rect 136876 2320 136882 2372
rect 136928 2360 136956 2536
rect 137986 2536 138336 2564
rect 137986 2360 138014 2536
rect 138106 2388 138112 2440
rect 138164 2388 138170 2440
rect 136928 2332 138014 2360
rect 138308 2360 138336 2536
rect 140682 2524 140688 2576
rect 140740 2564 140746 2576
rect 140961 2567 141019 2573
rect 140961 2564 140973 2567
rect 140740 2536 140973 2564
rect 140740 2524 140746 2536
rect 140961 2533 140973 2536
rect 141007 2533 141019 2567
rect 140961 2527 141019 2533
rect 155862 2524 155868 2576
rect 155920 2564 155926 2576
rect 156417 2567 156475 2573
rect 156417 2564 156429 2567
rect 155920 2536 156429 2564
rect 155920 2524 155926 2536
rect 156417 2533 156429 2536
rect 156463 2533 156475 2567
rect 156417 2527 156475 2533
rect 138382 2456 138388 2508
rect 138440 2496 138446 2508
rect 180766 2496 180794 2604
rect 187326 2592 187332 2644
rect 187384 2592 187390 2644
rect 202782 2592 202788 2644
rect 202840 2592 202846 2644
rect 233050 2592 233056 2644
rect 233108 2632 233114 2644
rect 233697 2635 233755 2641
rect 233697 2632 233709 2635
rect 233108 2604 233709 2632
rect 233108 2592 233114 2604
rect 233697 2601 233709 2604
rect 233743 2601 233755 2635
rect 233697 2595 233755 2601
rect 244274 2592 244280 2644
rect 244332 2632 244338 2644
rect 248046 2632 248052 2644
rect 244332 2604 248052 2632
rect 244332 2592 244338 2604
rect 248046 2592 248052 2604
rect 248104 2592 248110 2644
rect 249150 2592 249156 2644
rect 249208 2592 249214 2644
rect 273346 2592 273352 2644
rect 273404 2632 273410 2644
rect 273404 2604 294368 2632
rect 273404 2592 273410 2604
rect 218238 2524 218244 2576
rect 218296 2524 218302 2576
rect 238018 2524 238024 2576
rect 238076 2564 238082 2576
rect 247034 2564 247040 2576
rect 238076 2536 247040 2564
rect 238076 2524 238082 2536
rect 247034 2524 247040 2536
rect 247092 2524 247098 2576
rect 249242 2524 249248 2576
rect 249300 2564 249306 2576
rect 294340 2564 294368 2604
rect 295518 2592 295524 2644
rect 295576 2592 295582 2644
rect 367462 2632 367468 2644
rect 295628 2604 367468 2632
rect 295628 2564 295656 2604
rect 367462 2592 367468 2604
rect 367520 2592 367526 2644
rect 465258 2632 465264 2644
rect 371712 2604 465264 2632
rect 249300 2536 292574 2564
rect 294340 2536 295656 2564
rect 295720 2536 342116 2564
rect 249300 2524 249306 2536
rect 190549 2499 190607 2505
rect 190549 2496 190561 2499
rect 138440 2468 151814 2496
rect 180766 2468 190561 2496
rect 138440 2456 138446 2468
rect 141145 2431 141203 2437
rect 141145 2397 141157 2431
rect 141191 2428 141203 2431
rect 141694 2428 141700 2440
rect 141191 2400 141700 2428
rect 141191 2397 141203 2400
rect 141145 2391 141203 2397
rect 141694 2388 141700 2400
rect 141752 2388 141758 2440
rect 143721 2431 143779 2437
rect 143721 2397 143733 2431
rect 143767 2428 143779 2431
rect 143767 2400 144408 2428
rect 143767 2397 143779 2400
rect 143721 2391 143779 2397
rect 143169 2363 143227 2369
rect 143169 2360 143181 2363
rect 138308 2332 143181 2360
rect 143169 2329 143181 2332
rect 143215 2329 143227 2363
rect 143169 2323 143227 2329
rect 144380 2304 144408 2400
rect 151786 2360 151814 2468
rect 190549 2465 190561 2468
rect 190595 2465 190607 2499
rect 206741 2499 206799 2505
rect 190549 2459 190607 2465
rect 200086 2468 206048 2496
rect 156601 2431 156659 2437
rect 156601 2397 156613 2431
rect 156647 2428 156659 2431
rect 157150 2428 157156 2440
rect 156647 2400 157156 2428
rect 156647 2397 156659 2400
rect 156601 2391 156659 2397
rect 157150 2388 157156 2400
rect 157208 2388 157214 2440
rect 159177 2431 159235 2437
rect 159177 2397 159189 2431
rect 159223 2428 159235 2431
rect 159223 2400 159864 2428
rect 159223 2397 159235 2400
rect 159177 2391 159235 2397
rect 158625 2363 158683 2369
rect 158625 2360 158637 2363
rect 151786 2332 158637 2360
rect 158625 2329 158637 2332
rect 158671 2329 158683 2363
rect 158625 2323 158683 2329
rect 159836 2304 159864 2400
rect 171594 2388 171600 2440
rect 171652 2428 171658 2440
rect 172057 2431 172115 2437
rect 172057 2428 172069 2431
rect 171652 2400 172069 2428
rect 171652 2388 171658 2400
rect 172057 2397 172069 2400
rect 172103 2397 172115 2431
rect 172057 2391 172115 2397
rect 187513 2431 187571 2437
rect 187513 2397 187525 2431
rect 187559 2397 187571 2431
rect 187513 2391 187571 2397
rect 188893 2431 188951 2437
rect 188893 2397 188905 2431
rect 188939 2428 188951 2431
rect 189534 2428 189540 2440
rect 188939 2400 189540 2428
rect 188939 2397 188951 2400
rect 188893 2391 188951 2397
rect 138198 2292 138204 2304
rect 128326 2264 138204 2292
rect 138198 2252 138204 2264
rect 138256 2252 138262 2304
rect 138290 2252 138296 2304
rect 138348 2252 138354 2304
rect 141694 2252 141700 2304
rect 141752 2252 141758 2304
rect 144362 2252 144368 2304
rect 144420 2252 144426 2304
rect 157150 2252 157156 2304
rect 157208 2252 157214 2304
rect 159818 2252 159824 2304
rect 159876 2252 159882 2304
rect 171870 2252 171876 2304
rect 171928 2252 171934 2304
rect 187528 2292 187556 2391
rect 189534 2388 189540 2400
rect 189592 2388 189598 2440
rect 190825 2431 190883 2437
rect 190825 2397 190837 2431
rect 190871 2428 190883 2431
rect 191374 2428 191380 2440
rect 190871 2400 191380 2428
rect 190871 2397 190883 2400
rect 190825 2391 190883 2397
rect 191374 2388 191380 2400
rect 191432 2388 191438 2440
rect 188614 2320 188620 2372
rect 188672 2320 188678 2372
rect 200086 2360 200114 2468
rect 202966 2388 202972 2440
rect 203024 2388 203030 2440
rect 204165 2431 204223 2437
rect 204165 2397 204177 2431
rect 204211 2428 204223 2431
rect 204211 2400 205036 2428
rect 204211 2397 204223 2400
rect 204165 2391 204223 2397
rect 190840 2332 200114 2360
rect 187694 2292 187700 2304
rect 187528 2264 187700 2292
rect 187694 2252 187700 2264
rect 187752 2292 187758 2304
rect 190840 2292 190868 2332
rect 203886 2320 203892 2372
rect 203944 2320 203950 2372
rect 187752 2264 190868 2292
rect 187752 2252 187758 2264
rect 191374 2252 191380 2304
rect 191432 2252 191438 2304
rect 205008 2301 205036 2400
rect 205910 2320 205916 2372
rect 205968 2320 205974 2372
rect 206020 2360 206048 2468
rect 206741 2465 206753 2499
rect 206787 2496 206799 2499
rect 228174 2496 228180 2508
rect 206787 2468 228180 2496
rect 206787 2465 206799 2468
rect 206741 2459 206799 2465
rect 206189 2431 206247 2437
rect 206189 2397 206201 2431
rect 206235 2428 206247 2431
rect 206756 2428 206784 2459
rect 228174 2456 228180 2468
rect 228232 2456 228238 2508
rect 240134 2456 240140 2508
rect 240192 2496 240198 2508
rect 292546 2496 292574 2536
rect 295720 2496 295748 2536
rect 240192 2468 253934 2496
rect 240192 2456 240198 2468
rect 206235 2400 206784 2428
rect 206235 2397 206247 2400
rect 206189 2391 206247 2397
rect 218054 2388 218060 2440
rect 218112 2428 218118 2440
rect 218425 2431 218483 2437
rect 218425 2428 218437 2431
rect 218112 2400 218437 2428
rect 218112 2388 218118 2400
rect 218425 2397 218437 2400
rect 218471 2397 218483 2431
rect 218425 2391 218483 2397
rect 233881 2431 233939 2437
rect 233881 2397 233893 2431
rect 233927 2428 233939 2431
rect 246761 2431 246819 2437
rect 246761 2428 246773 2431
rect 233927 2400 234384 2428
rect 233927 2397 233939 2400
rect 233881 2391 233939 2397
rect 232682 2360 232688 2372
rect 206020 2332 232688 2360
rect 232682 2320 232688 2332
rect 232740 2320 232746 2372
rect 234356 2304 234384 2400
rect 246224 2400 246773 2428
rect 204993 2295 205051 2301
rect 204993 2261 205005 2295
rect 205039 2292 205051 2295
rect 230658 2292 230664 2304
rect 205039 2264 230664 2292
rect 205039 2261 205051 2264
rect 204993 2255 205051 2261
rect 230658 2252 230664 2264
rect 230716 2252 230722 2304
rect 234338 2252 234344 2304
rect 234396 2252 234402 2304
rect 239582 2252 239588 2304
rect 239640 2292 239646 2304
rect 246224 2301 246252 2400
rect 246761 2397 246773 2400
rect 246807 2397 246819 2431
rect 246761 2391 246819 2397
rect 248046 2388 248052 2440
rect 248104 2428 248110 2440
rect 249337 2431 249395 2437
rect 249337 2428 249349 2431
rect 248104 2400 249349 2428
rect 248104 2388 248110 2400
rect 249337 2397 249349 2400
rect 249383 2397 249395 2431
rect 249337 2391 249395 2397
rect 247037 2363 247095 2369
rect 247037 2329 247049 2363
rect 247083 2360 247095 2363
rect 250438 2360 250444 2372
rect 247083 2332 250444 2360
rect 247083 2329 247095 2332
rect 247037 2323 247095 2329
rect 250438 2320 250444 2332
rect 250496 2320 250502 2372
rect 253906 2360 253934 2468
rect 258046 2468 291148 2496
rect 292546 2468 295748 2496
rect 258046 2360 258074 2468
rect 264330 2388 264336 2440
rect 264388 2428 264394 2440
rect 264793 2431 264851 2437
rect 264793 2428 264805 2431
rect 264388 2400 264805 2428
rect 264388 2388 264394 2400
rect 264793 2397 264805 2400
rect 264839 2397 264851 2431
rect 273073 2431 273131 2437
rect 273073 2428 273085 2431
rect 264793 2391 264851 2397
rect 272536 2400 273085 2428
rect 253906 2332 258074 2360
rect 272536 2304 272564 2400
rect 273073 2397 273085 2400
rect 273119 2397 273131 2431
rect 273073 2391 273131 2397
rect 273346 2388 273352 2440
rect 273404 2388 273410 2440
rect 275281 2431 275339 2437
rect 275281 2428 275293 2431
rect 274744 2400 275293 2428
rect 274744 2304 274772 2400
rect 275281 2397 275293 2400
rect 275327 2397 275339 2431
rect 275281 2391 275339 2397
rect 276014 2388 276020 2440
rect 276072 2428 276078 2440
rect 277210 2428 277216 2440
rect 276072 2400 277216 2428
rect 276072 2388 276078 2400
rect 277210 2388 277216 2400
rect 277268 2428 277274 2440
rect 277397 2431 277455 2437
rect 277397 2428 277409 2431
rect 277268 2400 277409 2428
rect 277268 2388 277274 2400
rect 277397 2397 277409 2400
rect 277443 2397 277455 2431
rect 280249 2431 280307 2437
rect 280249 2428 280261 2431
rect 277397 2391 277455 2397
rect 278976 2400 280261 2428
rect 275554 2320 275560 2372
rect 275612 2320 275618 2372
rect 277670 2320 277676 2372
rect 277728 2320 277734 2372
rect 278976 2304 279004 2400
rect 280249 2397 280261 2400
rect 280295 2397 280307 2431
rect 288529 2431 288587 2437
rect 288529 2428 288541 2431
rect 280249 2391 280307 2397
rect 287992 2400 288541 2428
rect 287992 2304 288020 2400
rect 288529 2397 288541 2400
rect 288575 2397 288587 2431
rect 290645 2431 290703 2437
rect 290645 2428 290657 2431
rect 288529 2391 288587 2397
rect 290200 2400 290657 2428
rect 290200 2372 290228 2400
rect 290645 2397 290657 2400
rect 290691 2397 290703 2431
rect 290645 2391 290703 2397
rect 288805 2363 288863 2369
rect 288805 2329 288817 2363
rect 288851 2329 288863 2363
rect 288805 2323 288863 2329
rect 246209 2295 246267 2301
rect 246209 2292 246221 2295
rect 239640 2264 246221 2292
rect 239640 2252 239646 2264
rect 246209 2261 246221 2264
rect 246255 2261 246267 2295
rect 246209 2255 246267 2261
rect 264606 2252 264612 2304
rect 264664 2252 264670 2304
rect 272518 2252 272524 2304
rect 272576 2252 272582 2304
rect 274726 2252 274732 2304
rect 274784 2252 274790 2304
rect 278958 2252 278964 2304
rect 279016 2252 279022 2304
rect 280062 2252 280068 2304
rect 280120 2252 280126 2304
rect 287974 2252 287980 2304
rect 288032 2252 288038 2304
rect 288820 2292 288848 2323
rect 290182 2320 290188 2372
rect 290240 2320 290246 2372
rect 290918 2320 290924 2372
rect 290976 2320 290982 2372
rect 291120 2360 291148 2468
rect 295794 2456 295800 2508
rect 295852 2496 295858 2508
rect 295852 2468 340920 2496
rect 295852 2456 295858 2468
rect 292850 2388 292856 2440
rect 292908 2388 292914 2440
rect 293328 2400 293540 2428
rect 293328 2360 293356 2400
rect 291120 2332 293356 2360
rect 293402 2320 293408 2372
rect 293460 2320 293466 2372
rect 293512 2360 293540 2400
rect 294414 2388 294420 2440
rect 294472 2428 294478 2440
rect 295705 2431 295763 2437
rect 295705 2428 295717 2431
rect 294472 2400 295717 2428
rect 294472 2388 294478 2400
rect 295705 2397 295717 2400
rect 295751 2397 295763 2431
rect 295705 2391 295763 2397
rect 310698 2388 310704 2440
rect 310756 2428 310762 2440
rect 311161 2431 311219 2437
rect 311161 2428 311173 2431
rect 310756 2400 311173 2428
rect 310756 2388 310762 2400
rect 311161 2397 311173 2400
rect 311207 2397 311219 2431
rect 311161 2391 311219 2397
rect 320910 2388 320916 2440
rect 320968 2428 320974 2440
rect 321557 2431 321615 2437
rect 321557 2428 321569 2431
rect 320968 2400 321569 2428
rect 320968 2388 320974 2400
rect 321557 2397 321569 2400
rect 321603 2397 321615 2431
rect 321557 2391 321615 2397
rect 323578 2388 323584 2440
rect 323636 2388 323642 2440
rect 324498 2428 324504 2440
rect 323688 2400 324504 2428
rect 293512 2332 295748 2360
rect 295610 2292 295616 2304
rect 288820 2264 295616 2292
rect 295610 2252 295616 2264
rect 295668 2252 295674 2304
rect 295720 2292 295748 2332
rect 302206 2332 322060 2360
rect 302206 2292 302234 2332
rect 295720 2264 302234 2292
rect 310974 2252 310980 2304
rect 311032 2252 311038 2304
rect 320910 2252 320916 2304
rect 320968 2252 320974 2304
rect 322032 2292 322060 2332
rect 322106 2320 322112 2372
rect 322164 2320 322170 2372
rect 323688 2292 323716 2400
rect 324498 2388 324504 2400
rect 324556 2428 324562 2440
rect 324777 2431 324835 2437
rect 324777 2428 324789 2431
rect 324556 2400 324789 2428
rect 324556 2388 324562 2400
rect 324777 2397 324789 2400
rect 324823 2397 324835 2431
rect 324777 2391 324835 2397
rect 326154 2388 326160 2440
rect 326212 2428 326218 2440
rect 326617 2431 326675 2437
rect 326617 2428 326629 2431
rect 326212 2400 326629 2428
rect 326212 2388 326218 2400
rect 326617 2397 326629 2400
rect 326663 2397 326675 2431
rect 326617 2391 326675 2397
rect 331582 2388 331588 2440
rect 331640 2388 331646 2440
rect 333054 2388 333060 2440
rect 333112 2388 333118 2440
rect 334618 2388 334624 2440
rect 334676 2388 334682 2440
rect 335722 2388 335728 2440
rect 335780 2388 335786 2440
rect 336458 2388 336464 2440
rect 336516 2388 336522 2440
rect 338206 2388 338212 2440
rect 338264 2388 338270 2440
rect 339589 2431 339647 2437
rect 339589 2397 339601 2431
rect 339635 2428 339647 2431
rect 339862 2428 339868 2440
rect 339635 2400 339868 2428
rect 339635 2397 339647 2400
rect 339589 2391 339647 2397
rect 339862 2388 339868 2400
rect 339920 2388 339926 2440
rect 340230 2388 340236 2440
rect 340288 2388 340294 2440
rect 324130 2320 324136 2372
rect 324188 2320 324194 2372
rect 325326 2320 325332 2372
rect 325384 2320 325390 2372
rect 331306 2320 331312 2372
rect 331364 2320 331370 2372
rect 332594 2320 332600 2372
rect 332652 2320 332658 2372
rect 334066 2320 334072 2372
rect 334124 2320 334130 2372
rect 335446 2320 335452 2372
rect 335504 2320 335510 2372
rect 337010 2320 337016 2372
rect 337068 2320 337074 2372
rect 337654 2320 337660 2372
rect 337712 2320 337718 2372
rect 339034 2320 339040 2372
rect 339092 2320 339098 2372
rect 340782 2320 340788 2372
rect 340840 2320 340846 2372
rect 340892 2360 340920 2468
rect 342088 2437 342116 2536
rect 344986 2468 371280 2496
rect 342073 2431 342131 2437
rect 342073 2397 342085 2431
rect 342119 2428 342131 2431
rect 342533 2431 342591 2437
rect 342533 2428 342545 2431
rect 342119 2400 342545 2428
rect 342119 2397 342131 2400
rect 342073 2391 342131 2397
rect 342533 2397 342545 2400
rect 342579 2397 342591 2431
rect 342533 2391 342591 2397
rect 344986 2360 345014 2468
rect 357066 2388 357072 2440
rect 357124 2428 357130 2440
rect 357437 2431 357495 2437
rect 357437 2428 357449 2431
rect 357124 2400 357449 2428
rect 357124 2388 357130 2400
rect 357437 2397 357449 2400
rect 357483 2397 357495 2431
rect 357437 2391 357495 2397
rect 367462 2388 367468 2440
rect 367520 2428 367526 2440
rect 367741 2431 367799 2437
rect 367741 2428 367753 2431
rect 367520 2400 367753 2428
rect 367520 2388 367526 2400
rect 367741 2397 367753 2400
rect 367787 2397 367799 2431
rect 369857 2431 369915 2437
rect 369857 2428 369869 2431
rect 367741 2391 367799 2397
rect 369136 2400 369869 2428
rect 340892 2332 345014 2360
rect 368290 2320 368296 2372
rect 368348 2320 368354 2372
rect 369136 2304 369164 2400
rect 369857 2397 369869 2400
rect 369903 2397 369915 2431
rect 369857 2391 369915 2397
rect 370314 2388 370320 2440
rect 370372 2428 370378 2440
rect 370866 2428 370872 2440
rect 370372 2400 370872 2428
rect 370372 2388 370378 2400
rect 370866 2388 370872 2400
rect 370924 2428 370930 2440
rect 371145 2431 371203 2437
rect 371145 2428 371157 2431
rect 370924 2400 371157 2428
rect 370924 2388 370930 2400
rect 371145 2397 371157 2400
rect 371191 2397 371203 2431
rect 371145 2391 371203 2397
rect 370406 2320 370412 2372
rect 370464 2320 370470 2372
rect 371252 2360 371280 2468
rect 371712 2437 371740 2604
rect 465258 2592 465264 2604
rect 465316 2592 465322 2644
rect 478874 2592 478880 2644
rect 478932 2632 478938 2644
rect 480993 2635 481051 2641
rect 480993 2632 481005 2635
rect 478932 2604 481005 2632
rect 478932 2592 478938 2604
rect 480993 2601 481005 2604
rect 481039 2601 481051 2635
rect 480993 2595 481051 2601
rect 510522 2592 510528 2644
rect 510580 2632 510586 2644
rect 511905 2635 511963 2641
rect 511905 2632 511917 2635
rect 510580 2604 511917 2632
rect 510580 2592 510586 2604
rect 511905 2601 511917 2604
rect 511951 2601 511963 2635
rect 604454 2632 604460 2644
rect 511905 2595 511963 2601
rect 518866 2604 604460 2632
rect 372798 2524 372804 2576
rect 372856 2524 372862 2576
rect 388254 2524 388260 2576
rect 388312 2524 388318 2576
rect 478690 2564 478696 2576
rect 393286 2536 478696 2564
rect 385865 2499 385923 2505
rect 385865 2465 385877 2499
rect 385911 2496 385923 2499
rect 393286 2496 393314 2536
rect 478690 2524 478696 2536
rect 478748 2524 478754 2576
rect 385911 2468 393314 2496
rect 418065 2499 418123 2505
rect 385911 2465 385923 2468
rect 385865 2459 385923 2465
rect 418065 2465 418077 2499
rect 418111 2496 418123 2499
rect 478785 2499 478843 2505
rect 418111 2468 441614 2496
rect 418111 2465 418123 2468
rect 418065 2459 418123 2465
rect 371697 2431 371755 2437
rect 371697 2397 371709 2431
rect 371743 2397 371755 2431
rect 371697 2391 371755 2397
rect 372982 2388 372988 2440
rect 373040 2388 373046 2440
rect 383105 2431 383163 2437
rect 383105 2397 383117 2431
rect 383151 2397 383163 2431
rect 385313 2431 385371 2437
rect 385313 2428 385325 2431
rect 383105 2391 383163 2397
rect 384592 2400 385325 2428
rect 382826 2360 382832 2372
rect 371252 2332 382832 2360
rect 382826 2320 382832 2332
rect 382884 2360 382890 2372
rect 383120 2360 383148 2391
rect 382884 2332 383148 2360
rect 382884 2320 382890 2332
rect 383654 2320 383660 2372
rect 383712 2320 383718 2372
rect 384592 2304 384620 2400
rect 385313 2397 385325 2400
rect 385359 2397 385371 2431
rect 385313 2391 385371 2397
rect 386598 2388 386604 2440
rect 386656 2388 386662 2440
rect 388438 2388 388444 2440
rect 388496 2388 388502 2440
rect 403434 2388 403440 2440
rect 403492 2428 403498 2440
rect 403897 2431 403955 2437
rect 403897 2428 403909 2431
rect 403492 2400 403909 2428
rect 403492 2388 403498 2400
rect 403897 2397 403909 2400
rect 403943 2397 403955 2431
rect 416225 2431 416283 2437
rect 416225 2428 416237 2431
rect 403897 2391 403955 2397
rect 415504 2400 416237 2428
rect 387150 2320 387156 2372
rect 387208 2320 387214 2372
rect 415504 2304 415532 2400
rect 416225 2397 416237 2400
rect 416271 2397 416283 2431
rect 416225 2391 416283 2397
rect 417510 2388 417516 2440
rect 417568 2388 417574 2440
rect 418890 2388 418896 2440
rect 418948 2428 418954 2440
rect 419353 2431 419411 2437
rect 419353 2428 419365 2431
rect 418948 2400 419365 2428
rect 418948 2388 418954 2400
rect 419353 2397 419365 2400
rect 419399 2397 419411 2431
rect 419353 2391 419411 2397
rect 428461 2431 428519 2437
rect 428461 2397 428473 2431
rect 428507 2428 428519 2431
rect 430301 2431 430359 2437
rect 428507 2400 429148 2428
rect 428507 2397 428519 2400
rect 428461 2391 428519 2397
rect 416774 2320 416780 2372
rect 416832 2320 416838 2372
rect 428182 2320 428188 2372
rect 428240 2320 428246 2372
rect 429120 2304 429148 2400
rect 430301 2397 430313 2431
rect 430347 2428 430359 2431
rect 430347 2400 430988 2428
rect 430347 2397 430359 2400
rect 430301 2391 430359 2397
rect 429746 2320 429752 2372
rect 429804 2320 429810 2372
rect 430960 2304 430988 2400
rect 431678 2388 431684 2440
rect 431736 2388 431742 2440
rect 432233 2431 432291 2437
rect 432233 2397 432245 2431
rect 432279 2428 432291 2431
rect 433334 2428 433340 2440
rect 432279 2400 433340 2428
rect 432279 2397 432291 2400
rect 432233 2391 432291 2397
rect 433334 2388 433340 2400
rect 433392 2388 433398 2440
rect 433426 2388 433432 2440
rect 433484 2388 433490 2440
rect 434530 2388 434536 2440
rect 434588 2428 434594 2440
rect 434809 2431 434867 2437
rect 434809 2428 434821 2431
rect 434588 2400 434821 2428
rect 434588 2388 434594 2400
rect 434809 2397 434821 2400
rect 434855 2397 434867 2431
rect 434809 2391 434867 2397
rect 435913 2431 435971 2437
rect 435913 2397 435925 2431
rect 435959 2428 435971 2431
rect 441586 2428 441614 2468
rect 478785 2465 478797 2499
rect 478831 2496 478843 2499
rect 510801 2499 510859 2505
rect 478831 2468 510384 2496
rect 478831 2465 478843 2468
rect 478785 2459 478843 2465
rect 435959 2400 436876 2428
rect 441586 2400 451274 2428
rect 435959 2397 435971 2400
rect 435913 2391 435971 2397
rect 432874 2320 432880 2372
rect 432932 2320 432938 2372
rect 435358 2320 435364 2372
rect 435416 2320 435422 2372
rect 436848 2304 436876 2400
rect 449894 2320 449900 2372
rect 449952 2360 449958 2372
rect 450173 2363 450231 2369
rect 450173 2360 450185 2363
rect 449952 2332 450185 2360
rect 449952 2320 449958 2332
rect 450173 2329 450185 2332
rect 450219 2329 450231 2363
rect 451246 2360 451274 2400
rect 461854 2388 461860 2440
rect 461912 2428 461918 2440
rect 462501 2431 462559 2437
rect 462501 2428 462513 2431
rect 461912 2400 462513 2428
rect 461912 2388 461918 2400
rect 462501 2397 462513 2400
rect 462547 2397 462559 2431
rect 462501 2391 462559 2397
rect 463252 2400 463464 2428
rect 463252 2360 463280 2400
rect 451246 2332 463280 2360
rect 450173 2323 450231 2329
rect 463326 2320 463332 2372
rect 463384 2320 463390 2372
rect 463436 2360 463464 2400
rect 465258 2388 465264 2440
rect 465316 2428 465322 2440
rect 465721 2431 465779 2437
rect 465721 2428 465733 2431
rect 465316 2400 465733 2428
rect 465316 2388 465322 2400
rect 465721 2397 465733 2400
rect 465767 2397 465779 2431
rect 465721 2391 465779 2397
rect 477310 2388 477316 2440
rect 477368 2428 477374 2440
rect 477957 2431 478015 2437
rect 477957 2428 477969 2431
rect 477368 2400 477969 2428
rect 477368 2388 477374 2400
rect 477957 2397 477969 2400
rect 478003 2397 478015 2431
rect 477957 2391 478015 2397
rect 480714 2388 480720 2440
rect 480772 2428 480778 2440
rect 481177 2431 481235 2437
rect 481177 2428 481189 2431
rect 480772 2400 481189 2428
rect 480772 2388 480778 2400
rect 481177 2397 481189 2400
rect 481223 2397 481235 2431
rect 481177 2391 481235 2397
rect 496170 2388 496176 2440
rect 496228 2428 496234 2440
rect 496633 2431 496691 2437
rect 496633 2428 496645 2431
rect 496228 2400 496645 2428
rect 496228 2388 496234 2400
rect 496633 2397 496645 2400
rect 496679 2397 496691 2431
rect 496633 2391 496691 2397
rect 509694 2388 509700 2440
rect 509752 2428 509758 2440
rect 510249 2431 510307 2437
rect 510249 2428 510261 2431
rect 509752 2400 510261 2428
rect 509752 2388 509758 2400
rect 510249 2397 510261 2400
rect 510295 2397 510307 2431
rect 510249 2391 510307 2397
rect 510356 2360 510384 2468
rect 510801 2465 510813 2499
rect 510847 2496 510859 2499
rect 518866 2496 518894 2604
rect 604454 2592 604460 2604
rect 604512 2592 604518 2644
rect 604638 2592 604644 2644
rect 604696 2592 604702 2644
rect 620094 2592 620100 2644
rect 620152 2592 620158 2644
rect 625430 2592 625436 2644
rect 625488 2632 625494 2644
rect 626077 2635 626135 2641
rect 626077 2632 626089 2635
rect 625488 2604 626089 2632
rect 625488 2592 625494 2604
rect 626077 2601 626089 2604
rect 626123 2632 626135 2635
rect 681921 2635 681979 2641
rect 681921 2632 681933 2635
rect 626123 2604 681933 2632
rect 626123 2601 626135 2604
rect 626077 2595 626135 2601
rect 681921 2601 681933 2604
rect 681967 2601 681979 2635
rect 681921 2595 681979 2601
rect 525058 2524 525064 2576
rect 525116 2524 525122 2576
rect 619818 2564 619824 2576
rect 526272 2536 619824 2564
rect 510847 2468 518894 2496
rect 510847 2465 510859 2468
rect 510801 2459 510859 2465
rect 511626 2388 511632 2440
rect 511684 2428 511690 2440
rect 512089 2431 512147 2437
rect 512089 2428 512101 2431
rect 511684 2400 512101 2428
rect 511684 2388 511690 2400
rect 512089 2397 512101 2400
rect 512135 2397 512147 2431
rect 512089 2391 512147 2397
rect 525058 2388 525064 2440
rect 525116 2428 525122 2440
rect 526272 2437 526300 2536
rect 619818 2524 619824 2536
rect 619876 2524 619882 2576
rect 635737 2567 635795 2573
rect 635737 2564 635749 2567
rect 623240 2536 635749 2564
rect 570785 2499 570843 2505
rect 570785 2496 570797 2499
rect 526364 2468 570797 2496
rect 525705 2431 525763 2437
rect 525705 2428 525717 2431
rect 525116 2400 525717 2428
rect 525116 2388 525122 2400
rect 525705 2397 525717 2400
rect 525751 2397 525763 2431
rect 525705 2391 525763 2397
rect 526257 2431 526315 2437
rect 526257 2397 526269 2431
rect 526303 2397 526315 2431
rect 526257 2391 526315 2397
rect 526364 2360 526392 2468
rect 570785 2465 570797 2468
rect 570831 2496 570843 2499
rect 572533 2499 572591 2505
rect 570831 2468 571380 2496
rect 570831 2465 570843 2468
rect 570785 2459 570843 2465
rect 527542 2388 527548 2440
rect 527600 2388 527606 2440
rect 528830 2388 528836 2440
rect 528888 2388 528894 2440
rect 530305 2431 530363 2437
rect 530305 2397 530317 2431
rect 530351 2428 530363 2431
rect 530351 2400 530992 2428
rect 530351 2397 530363 2400
rect 530305 2391 530363 2397
rect 463436 2332 477448 2360
rect 322032 2264 323716 2292
rect 326430 2252 326436 2304
rect 326488 2252 326494 2304
rect 341886 2252 341892 2304
rect 341944 2252 341950 2304
rect 357342 2252 357348 2304
rect 357400 2252 357406 2304
rect 369118 2252 369124 2304
rect 369176 2252 369182 2304
rect 384574 2252 384580 2304
rect 384632 2252 384638 2304
rect 403710 2252 403716 2304
rect 403768 2252 403774 2304
rect 415486 2252 415492 2304
rect 415544 2252 415550 2304
rect 419166 2252 419172 2304
rect 419224 2252 419230 2304
rect 429102 2252 429108 2304
rect 429160 2252 429166 2304
rect 430942 2252 430948 2304
rect 431000 2252 431006 2304
rect 434622 2252 434628 2304
rect 434680 2252 434686 2304
rect 436830 2252 436836 2304
rect 436888 2252 436894 2304
rect 450078 2252 450084 2304
rect 450136 2252 450142 2304
rect 461854 2252 461860 2304
rect 461912 2252 461918 2304
rect 464982 2252 464988 2304
rect 465040 2292 465046 2304
rect 465537 2295 465595 2301
rect 465537 2292 465549 2295
rect 465040 2264 465549 2292
rect 465040 2252 465046 2264
rect 465537 2261 465549 2264
rect 465583 2261 465595 2295
rect 465537 2255 465595 2261
rect 477310 2252 477316 2304
rect 477368 2252 477374 2304
rect 477420 2292 477448 2332
rect 480226 2332 509234 2360
rect 510356 2332 526392 2360
rect 480226 2292 480254 2332
rect 477420 2264 480254 2292
rect 496446 2252 496452 2304
rect 496504 2252 496510 2304
rect 509206 2292 509234 2332
rect 528278 2320 528284 2372
rect 528336 2320 528342 2372
rect 529750 2320 529756 2372
rect 529808 2320 529814 2372
rect 530964 2304 530992 2400
rect 542262 2388 542268 2440
rect 542320 2428 542326 2440
rect 542817 2431 542875 2437
rect 542817 2428 542829 2431
rect 542320 2400 542829 2428
rect 542320 2388 542326 2400
rect 542817 2397 542829 2400
rect 542863 2428 542875 2431
rect 543461 2431 543519 2437
rect 543461 2428 543473 2431
rect 542863 2400 543473 2428
rect 542863 2397 542875 2400
rect 542817 2391 542875 2397
rect 543461 2397 543473 2400
rect 543507 2397 543519 2431
rect 555881 2431 555939 2437
rect 555881 2428 555893 2431
rect 543461 2391 543519 2397
rect 555344 2400 555893 2428
rect 555344 2304 555372 2400
rect 555881 2397 555893 2400
rect 555927 2397 555939 2431
rect 555881 2391 555939 2397
rect 558086 2388 558092 2440
rect 558144 2428 558150 2440
rect 571352 2437 571380 2468
rect 572533 2465 572545 2499
rect 572579 2496 572591 2499
rect 572579 2468 623176 2496
rect 572579 2465 572591 2468
rect 572533 2459 572591 2465
rect 558457 2431 558515 2437
rect 558457 2428 558469 2431
rect 558144 2400 558469 2428
rect 558144 2388 558150 2400
rect 558457 2397 558469 2400
rect 558503 2397 558515 2431
rect 558457 2391 558515 2397
rect 571337 2431 571395 2437
rect 571337 2397 571349 2431
rect 571383 2397 571395 2431
rect 571337 2391 571395 2397
rect 571996 2400 572392 2428
rect 557077 2363 557135 2369
rect 557077 2329 557089 2363
rect 557123 2360 557135 2363
rect 571996 2360 572024 2400
rect 557123 2332 572024 2360
rect 572364 2360 572392 2400
rect 573910 2388 573916 2440
rect 573968 2388 573974 2440
rect 588906 2388 588912 2440
rect 588964 2428 588970 2440
rect 589369 2431 589427 2437
rect 589369 2428 589381 2431
rect 588964 2400 589381 2428
rect 588964 2388 588970 2400
rect 589369 2397 589381 2400
rect 589415 2397 589427 2431
rect 589369 2391 589427 2397
rect 604454 2388 604460 2440
rect 604512 2428 604518 2440
rect 604825 2431 604883 2437
rect 604825 2428 604837 2431
rect 604512 2400 604837 2428
rect 604512 2388 604518 2400
rect 604825 2397 604837 2400
rect 604871 2397 604883 2431
rect 604825 2391 604883 2397
rect 619818 2388 619824 2440
rect 619876 2428 619882 2440
rect 620281 2431 620339 2437
rect 620281 2428 620293 2431
rect 619876 2400 620293 2428
rect 619876 2388 619882 2400
rect 620281 2397 620293 2400
rect 620327 2397 620339 2431
rect 620281 2391 620339 2397
rect 572364 2332 620324 2360
rect 557123 2329 557135 2332
rect 557077 2323 557135 2329
rect 511626 2292 511632 2304
rect 509206 2264 511632 2292
rect 511626 2252 511632 2264
rect 511684 2252 511690 2304
rect 527082 2252 527088 2304
rect 527140 2292 527146 2304
rect 527361 2295 527419 2301
rect 527361 2292 527373 2295
rect 527140 2264 527373 2292
rect 527140 2252 527146 2264
rect 527361 2261 527373 2264
rect 527407 2261 527419 2295
rect 527361 2255 527419 2261
rect 530946 2252 530952 2304
rect 531004 2252 531010 2304
rect 539502 2252 539508 2304
rect 539560 2292 539566 2304
rect 543001 2295 543059 2301
rect 543001 2292 543013 2295
rect 539560 2264 543013 2292
rect 539560 2252 539566 2264
rect 543001 2261 543013 2264
rect 543047 2261 543059 2295
rect 543001 2255 543059 2261
rect 555326 2252 555332 2304
rect 555384 2252 555390 2304
rect 556154 2252 556160 2304
rect 556212 2292 556218 2304
rect 558273 2295 558331 2301
rect 558273 2292 558285 2295
rect 556212 2264 558285 2292
rect 556212 2252 556218 2264
rect 558273 2261 558285 2264
rect 558319 2261 558331 2295
rect 558273 2255 558331 2261
rect 572622 2252 572628 2304
rect 572680 2292 572686 2304
rect 573729 2295 573787 2301
rect 573729 2292 573741 2295
rect 572680 2264 573741 2292
rect 572680 2252 572686 2264
rect 573729 2261 573741 2264
rect 573775 2261 573787 2295
rect 573729 2255 573787 2261
rect 589182 2252 589188 2304
rect 589240 2252 589246 2304
rect 620296 2292 620324 2332
rect 623038 2320 623044 2372
rect 623096 2320 623102 2372
rect 623148 2360 623176 2468
rect 623240 2428 623268 2536
rect 635737 2533 635749 2536
rect 635783 2533 635795 2567
rect 635737 2527 635795 2533
rect 651006 2524 651012 2576
rect 651064 2524 651070 2576
rect 666462 2524 666468 2576
rect 666520 2524 666526 2576
rect 666186 2496 666192 2508
rect 625126 2468 666192 2496
rect 623317 2431 623375 2437
rect 623317 2428 623329 2431
rect 623240 2400 623329 2428
rect 623317 2397 623329 2400
rect 623363 2397 623375 2431
rect 625126 2428 625154 2468
rect 666186 2456 666192 2468
rect 666244 2496 666250 2508
rect 666244 2468 666692 2496
rect 666244 2456 666250 2468
rect 623317 2391 623375 2397
rect 623424 2400 625154 2428
rect 623424 2360 623452 2400
rect 625430 2388 625436 2440
rect 625488 2388 625494 2440
rect 635550 2388 635556 2440
rect 635608 2428 635614 2440
rect 666664 2437 666692 2468
rect 636197 2431 636255 2437
rect 636197 2428 636209 2431
rect 635608 2400 636209 2428
rect 635608 2388 635614 2400
rect 636197 2397 636209 2400
rect 636243 2397 636255 2431
rect 636197 2391 636255 2397
rect 651193 2431 651251 2437
rect 651193 2397 651205 2431
rect 651239 2397 651251 2431
rect 651193 2391 651251 2397
rect 666649 2431 666707 2437
rect 666649 2397 666661 2431
rect 666695 2397 666707 2431
rect 666649 2391 666707 2397
rect 623148 2332 623452 2360
rect 624878 2320 624884 2372
rect 624936 2320 624942 2372
rect 650730 2360 650736 2372
rect 625126 2332 650736 2360
rect 625126 2292 625154 2332
rect 650730 2320 650736 2332
rect 650788 2360 650794 2372
rect 651208 2360 651236 2391
rect 681734 2388 681740 2440
rect 681792 2428 681798 2440
rect 682105 2431 682163 2437
rect 682105 2428 682117 2431
rect 681792 2400 682117 2428
rect 681792 2388 681798 2400
rect 682105 2397 682117 2400
rect 682151 2397 682163 2431
rect 682105 2391 682163 2397
rect 650788 2332 651236 2360
rect 650788 2320 650794 2332
rect 620296 2264 625154 2292
rect 1104 2202 682824 2224
rect 1104 2150 86825 2202
rect 86877 2150 86889 2202
rect 86941 2150 86953 2202
rect 87005 2150 87017 2202
rect 87069 2150 87081 2202
rect 87133 2150 257255 2202
rect 257307 2150 257319 2202
rect 257371 2150 257383 2202
rect 257435 2150 257447 2202
rect 257499 2150 257511 2202
rect 257563 2150 427685 2202
rect 427737 2150 427749 2202
rect 427801 2150 427813 2202
rect 427865 2150 427877 2202
rect 427929 2150 427941 2202
rect 427993 2150 598115 2202
rect 598167 2150 598179 2202
rect 598231 2150 598243 2202
rect 598295 2150 598307 2202
rect 598359 2150 598371 2202
rect 598423 2150 682824 2202
rect 1104 2128 682824 2150
rect 2590 2048 2596 2100
rect 2648 2088 2654 2100
rect 96798 2088 96804 2100
rect 2648 2060 96804 2088
rect 2648 2048 2654 2060
rect 96798 2048 96804 2060
rect 96856 2048 96862 2100
rect 110690 2048 110696 2100
rect 110748 2088 110754 2100
rect 203886 2088 203892 2100
rect 110748 2060 203892 2088
rect 110748 2048 110754 2060
rect 203886 2048 203892 2060
rect 203944 2048 203950 2100
rect 218238 2048 218244 2100
rect 218296 2088 218302 2100
rect 231762 2088 231768 2100
rect 218296 2060 231768 2088
rect 218296 2048 218302 2060
rect 231762 2048 231768 2060
rect 231820 2048 231826 2100
rect 243262 2048 243268 2100
rect 243320 2088 243326 2100
rect 274726 2088 274732 2100
rect 243320 2060 274732 2088
rect 243320 2048 243326 2060
rect 274726 2048 274732 2060
rect 274784 2048 274790 2100
rect 290918 2048 290924 2100
rect 290976 2088 290982 2100
rect 384574 2088 384580 2100
rect 290976 2060 384580 2088
rect 290976 2048 290982 2060
rect 384574 2048 384580 2060
rect 384632 2048 384638 2100
rect 416774 2048 416780 2100
rect 416832 2088 416838 2100
rect 509694 2088 509700 2100
rect 416832 2060 509700 2088
rect 416832 2048 416838 2060
rect 509694 2048 509700 2060
rect 509752 2048 509758 2100
rect 528186 2048 528192 2100
rect 528244 2088 528250 2100
rect 589182 2088 589188 2100
rect 528244 2060 589188 2088
rect 528244 2048 528250 2060
rect 589182 2048 589188 2060
rect 589240 2048 589246 2100
rect 79134 1980 79140 2032
rect 79192 2020 79198 2032
rect 136542 2020 136548 2032
rect 79192 1992 136548 2020
rect 79192 1980 79198 1992
rect 136542 1980 136548 1992
rect 136600 1980 136606 2032
rect 235534 1980 235540 2032
rect 235592 2020 235598 2032
rect 278958 2020 278964 2032
rect 235592 1992 278964 2020
rect 235592 1980 235598 1992
rect 278958 1980 278964 1992
rect 279016 1980 279022 2032
rect 322106 1980 322112 2032
rect 322164 2020 322170 2032
rect 415486 2020 415492 2032
rect 322164 1992 415492 2020
rect 322164 1980 322170 1992
rect 415486 1980 415492 1992
rect 415544 1980 415550 2032
rect 429102 1980 429108 2032
rect 429160 2020 429166 2032
rect 450078 2020 450084 2032
rect 429160 1992 450084 2020
rect 429160 1980 429166 1992
rect 450078 1980 450084 1992
rect 450136 1980 450142 2032
rect 463326 1980 463332 2032
rect 463384 2020 463390 2032
rect 555326 2020 555332 2032
rect 463384 1992 555332 2020
rect 463384 1980 463390 1992
rect 555326 1980 555332 1992
rect 555384 1980 555390 2032
rect 18046 1912 18052 1964
rect 18104 1952 18110 1964
rect 112254 1952 112260 1964
rect 18104 1924 112260 1952
rect 18104 1912 18110 1924
rect 112254 1912 112260 1924
rect 112312 1912 112318 1964
rect 125686 1912 125692 1964
rect 125744 1952 125750 1964
rect 138106 1952 138112 1964
rect 125744 1924 138112 1952
rect 125744 1912 125750 1924
rect 138106 1912 138112 1924
rect 138164 1912 138170 1964
rect 235994 1912 236000 1964
rect 236052 1952 236058 1964
rect 244182 1952 244188 1964
rect 236052 1924 244188 1952
rect 236052 1912 236058 1924
rect 244182 1912 244188 1924
rect 244240 1912 244246 1964
rect 244366 1912 244372 1964
rect 244424 1952 244430 1964
rect 290182 1952 290188 1964
rect 244424 1924 290188 1952
rect 244424 1912 244430 1924
rect 290182 1912 290188 1924
rect 290240 1912 290246 1964
rect 293402 1912 293408 1964
rect 293460 1952 293466 1964
rect 386598 1952 386604 1964
rect 293460 1924 386604 1952
rect 293460 1912 293466 1924
rect 386598 1912 386604 1924
rect 386656 1912 386662 1964
rect 530946 1912 530952 1964
rect 531004 1952 531010 1964
rect 624878 1952 624884 1964
rect 531004 1924 624884 1952
rect 531004 1912 531010 1924
rect 624878 1912 624884 1924
rect 624936 1912 624942 1964
rect 238478 1844 238484 1896
rect 238536 1884 238542 1896
rect 249702 1884 249708 1896
rect 238536 1856 249708 1884
rect 238536 1844 238542 1856
rect 249702 1844 249708 1856
rect 249760 1844 249766 1896
rect 277670 1844 277676 1896
rect 277728 1884 277734 1896
rect 370314 1884 370320 1896
rect 277728 1856 370320 1884
rect 277728 1844 277734 1856
rect 370314 1844 370320 1856
rect 370372 1844 370378 1896
rect 370406 1844 370412 1896
rect 370464 1884 370470 1896
rect 463234 1884 463240 1896
rect 370464 1856 463240 1884
rect 370464 1844 370470 1856
rect 463234 1844 463240 1856
rect 463292 1844 463298 1896
rect 528830 1844 528836 1896
rect 528888 1884 528894 1896
rect 623038 1884 623044 1896
rect 528888 1856 623044 1884
rect 528888 1844 528894 1856
rect 623038 1844 623044 1856
rect 623096 1844 623102 1896
rect 95326 1776 95332 1828
rect 95384 1816 95390 1828
rect 188614 1816 188620 1828
rect 95384 1788 188620 1816
rect 95384 1776 95390 1788
rect 188614 1776 188620 1788
rect 188672 1776 188678 1828
rect 244090 1776 244096 1828
rect 244148 1816 244154 1828
rect 320910 1816 320916 1828
rect 244148 1788 320916 1816
rect 244148 1776 244154 1788
rect 320910 1776 320916 1788
rect 320968 1776 320974 1828
rect 342714 1776 342720 1828
rect 342772 1816 342778 1828
rect 435358 1816 435364 1828
rect 342772 1788 435364 1816
rect 342772 1776 342778 1788
rect 435358 1776 435364 1788
rect 435416 1776 435422 1828
rect 436830 1776 436836 1828
rect 436888 1816 436894 1828
rect 529750 1816 529756 1828
rect 436888 1788 529756 1816
rect 436888 1776 436894 1788
rect 529750 1776 529756 1788
rect 529808 1776 529814 1828
rect 113450 1708 113456 1760
rect 113508 1748 113514 1760
rect 205910 1748 205916 1760
rect 113508 1720 205916 1748
rect 113508 1708 113514 1720
rect 205910 1708 205916 1720
rect 205968 1708 205974 1760
rect 244182 1708 244188 1760
rect 244240 1748 244246 1760
rect 294414 1748 294420 1760
rect 244240 1720 294420 1748
rect 244240 1708 244246 1720
rect 294414 1708 294420 1720
rect 294472 1708 294478 1760
rect 331582 1708 331588 1760
rect 331640 1748 331646 1760
rect 357342 1748 357348 1760
rect 331640 1720 357348 1748
rect 331640 1708 331646 1720
rect 357342 1708 357348 1720
rect 357400 1708 357406 1760
rect 430942 1708 430948 1760
rect 431000 1748 431006 1760
rect 496446 1748 496452 1760
rect 431000 1720 496452 1748
rect 431000 1708 431006 1720
rect 496446 1708 496452 1720
rect 496504 1708 496510 1760
rect 241514 1640 241520 1692
rect 241572 1680 241578 1692
rect 241572 1652 246436 1680
rect 241572 1640 241578 1652
rect 246298 1612 246304 1624
rect 241486 1584 246304 1612
rect 232222 1476 232228 1488
rect 227548 1448 232228 1476
rect 189534 1300 189540 1352
rect 189592 1340 189598 1352
rect 227254 1340 227260 1352
rect 189592 1312 227260 1340
rect 189592 1300 189598 1312
rect 227254 1300 227260 1312
rect 227312 1300 227318 1352
rect 227548 1340 227576 1448
rect 232222 1436 232228 1448
rect 232280 1436 232286 1488
rect 235258 1436 235264 1488
rect 235316 1476 235322 1488
rect 241486 1476 241514 1584
rect 246298 1572 246304 1584
rect 246356 1572 246362 1624
rect 246408 1612 246436 1652
rect 246482 1640 246488 1692
rect 246540 1680 246546 1692
rect 276014 1680 276020 1692
rect 246540 1652 276020 1680
rect 246540 1640 246546 1652
rect 276014 1640 276020 1652
rect 276072 1640 276078 1692
rect 324130 1640 324136 1692
rect 324188 1680 324194 1692
rect 417510 1680 417516 1692
rect 324188 1652 417516 1680
rect 324188 1640 324194 1652
rect 417510 1640 417516 1652
rect 417568 1640 417574 1692
rect 435450 1640 435456 1692
rect 435508 1680 435514 1692
rect 528278 1680 528284 1692
rect 435508 1652 528284 1680
rect 435508 1640 435514 1652
rect 528278 1640 528284 1652
rect 528336 1640 528342 1692
rect 246408 1584 253934 1612
rect 243538 1504 243544 1556
rect 243596 1544 243602 1556
rect 244274 1544 244280 1556
rect 243596 1516 244280 1544
rect 243596 1504 243602 1516
rect 244274 1504 244280 1516
rect 244332 1504 244338 1556
rect 253906 1544 253934 1584
rect 275554 1572 275560 1624
rect 275612 1612 275618 1624
rect 369118 1612 369124 1624
rect 275612 1584 369124 1612
rect 275612 1572 275618 1584
rect 369118 1572 369124 1584
rect 369176 1572 369182 1624
rect 383654 1572 383660 1624
rect 383712 1612 383718 1624
rect 477310 1612 477316 1624
rect 383712 1584 477316 1612
rect 383712 1572 383718 1584
rect 477310 1572 477316 1584
rect 477368 1572 477374 1624
rect 292850 1544 292856 1556
rect 253906 1516 292856 1544
rect 292850 1504 292856 1516
rect 292908 1504 292914 1556
rect 325326 1504 325332 1556
rect 325384 1544 325390 1556
rect 418890 1544 418896 1556
rect 325384 1516 418896 1544
rect 325384 1504 325390 1516
rect 418890 1504 418896 1516
rect 418948 1504 418954 1556
rect 235316 1448 241514 1476
rect 235316 1436 235322 1448
rect 241882 1436 241888 1488
rect 241940 1476 241946 1488
rect 246482 1476 246488 1488
rect 241940 1448 246488 1476
rect 241940 1436 241946 1448
rect 246482 1436 246488 1448
rect 246540 1436 246546 1488
rect 250438 1436 250444 1488
rect 250496 1476 250502 1488
rect 340230 1476 340236 1488
rect 250496 1448 340236 1476
rect 250496 1436 250502 1448
rect 340230 1436 340236 1448
rect 340288 1436 340294 1488
rect 387150 1436 387156 1488
rect 387208 1476 387214 1488
rect 480714 1476 480720 1488
rect 387208 1448 480720 1476
rect 387208 1436 387214 1448
rect 480714 1436 480720 1448
rect 480772 1436 480778 1488
rect 231762 1368 231768 1420
rect 231820 1408 231826 1420
rect 231820 1380 233464 1408
rect 231820 1368 231826 1380
rect 227456 1312 227576 1340
rect 171870 1232 171876 1284
rect 171928 1272 171934 1284
rect 227456 1272 227484 1312
rect 227806 1300 227812 1352
rect 227864 1340 227870 1352
rect 227864 1312 233356 1340
rect 227864 1300 227870 1312
rect 229370 1272 229376 1284
rect 171928 1244 227484 1272
rect 227548 1244 229376 1272
rect 171928 1232 171934 1244
rect 159818 1164 159824 1216
rect 159876 1204 159882 1216
rect 227548 1204 227576 1244
rect 229370 1232 229376 1244
rect 229428 1232 229434 1284
rect 229462 1232 229468 1284
rect 229520 1272 229526 1284
rect 231946 1272 231952 1284
rect 229520 1244 231952 1272
rect 229520 1232 229526 1244
rect 231946 1232 231952 1244
rect 232004 1232 232010 1284
rect 159876 1176 227576 1204
rect 159876 1164 159882 1176
rect 227622 1164 227628 1216
rect 227680 1204 227686 1216
rect 227680 1176 231716 1204
rect 227680 1164 227686 1176
rect 157150 1096 157156 1148
rect 157208 1136 157214 1148
rect 227438 1136 227444 1148
rect 157208 1108 227444 1136
rect 157208 1096 157214 1108
rect 227438 1096 227444 1108
rect 227496 1096 227502 1148
rect 227714 1096 227720 1148
rect 227772 1136 227778 1148
rect 227772 1108 231302 1136
rect 227772 1096 227778 1108
rect 144362 1028 144368 1080
rect 144420 1068 144426 1080
rect 144420 1040 224080 1068
rect 144420 1028 144426 1040
rect 141694 960 141700 1012
rect 141752 1000 141758 1012
rect 141752 972 223988 1000
rect 141752 960 141758 972
rect 135990 892 135996 944
rect 136048 932 136054 944
rect 136048 904 223804 932
rect 136048 892 136054 904
rect 138290 824 138296 876
rect 138348 864 138354 876
rect 138348 836 219434 864
rect 138348 824 138354 836
rect 219406 660 219434 836
rect 223776 728 223804 904
rect 223960 796 223988 972
rect 224052 864 224080 1040
rect 224218 1028 224224 1080
rect 224276 1068 224282 1080
rect 228634 1068 228640 1080
rect 224276 1040 228640 1068
rect 224276 1028 224282 1040
rect 228634 1028 228640 1040
rect 228692 1028 228698 1080
rect 228726 1028 228732 1080
rect 228784 1068 228790 1080
rect 228784 1040 230500 1068
rect 228784 1028 228790 1040
rect 224310 960 224316 1012
rect 224368 1000 224374 1012
rect 224368 972 230106 1000
rect 224368 960 224374 972
rect 224236 904 228956 932
rect 224236 864 224264 904
rect 224052 836 224264 864
rect 227254 824 227260 876
rect 227312 864 227318 876
rect 228726 864 228732 876
rect 227312 836 228732 864
rect 227312 824 227318 836
rect 228726 824 228732 836
rect 228784 824 228790 876
rect 227622 796 227628 808
rect 223960 768 227628 796
rect 227622 756 227628 768
rect 227680 756 227686 808
rect 224126 728 224132 740
rect 223776 700 224132 728
rect 224126 688 224132 700
rect 224184 688 224190 740
rect 227714 660 227720 672
rect 219406 632 227720 660
rect 227714 620 227720 632
rect 227772 620 227778 672
rect 136818 212 136824 264
rect 136876 252 136882 264
rect 224126 252 224132 264
rect 136876 224 224132 252
rect 136876 212 136882 224
rect 224126 212 224132 224
rect 224184 212 224190 264
rect 202966 144 202972 196
rect 203024 184 203030 196
rect 227714 184 227720 196
rect 203024 156 227720 184
rect 203024 144 203030 156
rect 227714 144 227720 156
rect 227772 144 227778 196
rect 191374 8 191380 60
rect 191432 48 191438 60
rect 228010 48 228066 800
rect 228174 756 228180 808
rect 228232 796 228238 808
rect 228418 796 228474 800
rect 228232 768 228474 796
rect 228232 756 228238 768
rect 191432 20 228066 48
rect 191432 8 191438 20
rect 228010 0 228066 20
rect 228418 0 228474 768
rect 228634 756 228640 808
rect 228692 796 228698 808
rect 228826 796 228882 800
rect 228692 768 228882 796
rect 228692 756 228698 768
rect 228826 0 228882 768
rect 228928 728 228956 904
rect 230078 864 230106 972
rect 230472 864 230500 1040
rect 230032 836 230106 864
rect 230400 836 230500 864
rect 231274 864 231302 1108
rect 231688 864 231716 1176
rect 232222 1096 232228 1148
rect 232280 1136 232286 1148
rect 232280 1108 232544 1136
rect 232280 1096 232286 1108
rect 232516 864 232544 1108
rect 233328 864 233356 1312
rect 233436 1204 233464 1380
rect 241624 1380 242940 1408
rect 237190 1300 237196 1352
rect 237248 1340 237254 1352
rect 241624 1340 241652 1380
rect 237248 1312 241652 1340
rect 242912 1340 242940 1380
rect 243998 1368 244004 1420
rect 244056 1368 244062 1420
rect 244826 1368 244832 1420
rect 244884 1408 244890 1420
rect 323578 1408 323584 1420
rect 244884 1380 323584 1408
rect 244884 1368 244890 1380
rect 323578 1368 323584 1380
rect 323636 1368 323642 1420
rect 340782 1368 340788 1420
rect 340840 1408 340846 1420
rect 434530 1408 434536 1420
rect 340840 1380 434536 1408
rect 340840 1368 340846 1380
rect 434530 1368 434536 1380
rect 434588 1368 434594 1420
rect 244016 1340 244044 1368
rect 244550 1340 244556 1352
rect 242912 1312 243676 1340
rect 244016 1312 244556 1340
rect 237248 1300 237254 1312
rect 243538 1272 243544 1284
rect 235460 1244 243544 1272
rect 235460 1204 235488 1244
rect 243538 1232 243544 1244
rect 243596 1232 243602 1284
rect 243648 1272 243676 1312
rect 244550 1300 244556 1312
rect 244608 1300 244614 1352
rect 249426 1300 249432 1352
rect 249484 1340 249490 1352
rect 249484 1312 253934 1340
rect 249484 1300 249490 1312
rect 243648 1244 243860 1272
rect 239950 1204 239956 1216
rect 233436 1176 233764 1204
rect 233736 864 233764 1176
rect 231274 836 231348 864
rect 229234 728 229290 800
rect 229370 756 229376 808
rect 229428 796 229434 808
rect 230032 800 230060 836
rect 229642 796 229698 800
rect 229428 768 229698 796
rect 230032 768 230106 800
rect 230400 796 230428 836
rect 230458 796 230514 800
rect 230400 768 230514 796
rect 229428 756 229434 768
rect 228928 700 229290 728
rect 229234 0 229290 700
rect 229642 0 229698 768
rect 230050 0 230106 768
rect 230458 0 230514 768
rect 230658 756 230664 808
rect 230716 796 230722 808
rect 231320 800 231348 836
rect 230866 796 230922 800
rect 230716 768 230922 796
rect 230716 756 230722 768
rect 230866 0 230922 768
rect 231274 768 231348 800
rect 231596 836 231716 864
rect 232424 836 232544 864
rect 233252 836 233356 864
rect 233620 836 233764 864
rect 234540 1176 235488 1204
rect 236196 1176 239956 1204
rect 234540 864 234568 1176
rect 236196 864 236224 1176
rect 239950 1164 239956 1176
rect 240008 1164 240014 1216
rect 240042 1164 240048 1216
rect 240100 1204 240106 1216
rect 243630 1204 243636 1216
rect 240100 1176 243636 1204
rect 240100 1164 240106 1176
rect 243630 1164 243636 1176
rect 243688 1164 243694 1216
rect 243832 1204 243860 1244
rect 243906 1232 243912 1284
rect 243964 1272 243970 1284
rect 243964 1244 244412 1272
rect 243964 1232 243970 1244
rect 244274 1204 244280 1216
rect 243832 1176 244280 1204
rect 244274 1164 244280 1176
rect 244332 1164 244338 1216
rect 242066 1136 242072 1148
rect 237408 1108 242072 1136
rect 237408 864 237436 1108
rect 242066 1096 242072 1108
rect 242124 1096 242130 1148
rect 242526 1096 242532 1148
rect 242584 1136 242590 1148
rect 243998 1136 244004 1148
rect 242584 1108 244004 1136
rect 242584 1096 242590 1108
rect 243998 1096 244004 1108
rect 244056 1096 244062 1148
rect 244384 1136 244412 1244
rect 244826 1232 244832 1284
rect 244884 1272 244890 1284
rect 253906 1272 253934 1312
rect 338206 1300 338212 1352
rect 338264 1340 338270 1352
rect 432874 1340 432880 1352
rect 338264 1312 432880 1340
rect 338264 1300 338270 1312
rect 432874 1300 432880 1312
rect 432932 1300 432938 1352
rect 331306 1272 331312 1284
rect 244884 1244 251174 1272
rect 253906 1244 331312 1272
rect 244884 1232 244890 1244
rect 244734 1164 244740 1216
rect 244792 1204 244798 1216
rect 249150 1204 249156 1216
rect 244792 1176 249156 1204
rect 244792 1164 244798 1176
rect 249150 1164 249156 1176
rect 249208 1164 249214 1216
rect 251146 1204 251174 1244
rect 331306 1232 331312 1244
rect 331364 1232 331370 1284
rect 335722 1232 335728 1284
rect 335780 1272 335786 1284
rect 429746 1272 429752 1284
rect 335780 1244 429752 1272
rect 335780 1232 335786 1244
rect 429746 1232 429752 1244
rect 429804 1232 429810 1284
rect 251146 1176 253934 1204
rect 244826 1136 244832 1148
rect 244384 1108 244832 1136
rect 244826 1096 244832 1108
rect 244884 1096 244890 1148
rect 244918 1096 244924 1148
rect 244976 1136 244982 1148
rect 249334 1136 249340 1148
rect 244976 1108 249340 1136
rect 244976 1096 244982 1108
rect 249334 1096 249340 1108
rect 249392 1096 249398 1148
rect 253906 1136 253934 1176
rect 334618 1164 334624 1216
rect 334676 1204 334682 1216
rect 428182 1204 428188 1216
rect 334676 1176 428188 1204
rect 334676 1164 334682 1176
rect 428182 1164 428188 1176
rect 428240 1164 428246 1216
rect 337654 1136 337660 1148
rect 253906 1108 337660 1136
rect 337654 1096 337660 1108
rect 337712 1096 337718 1148
rect 368290 1096 368296 1148
rect 368348 1136 368354 1148
rect 461854 1136 461860 1148
rect 368348 1108 461860 1136
rect 368348 1096 368354 1108
rect 461854 1096 461860 1108
rect 461912 1096 461918 1148
rect 332594 1068 332600 1080
rect 238634 1040 242020 1068
rect 238634 864 238662 1040
rect 241882 1000 241888 1012
rect 240264 972 241888 1000
rect 240134 932 240140 944
rect 239324 904 240140 932
rect 234540 836 234614 864
rect 236196 836 236316 864
rect 237408 836 237512 864
rect 238634 836 238800 864
rect 231596 796 231624 836
rect 231682 796 231738 800
rect 231596 768 231738 796
rect 231274 0 231330 768
rect 231682 0 231738 768
rect 231946 620 231952 672
rect 232004 660 232010 672
rect 232090 660 232146 800
rect 232424 796 232452 836
rect 232498 796 232554 800
rect 232424 768 232554 796
rect 232004 632 232146 660
rect 232004 620 232010 632
rect 232090 0 232146 632
rect 232498 0 232554 768
rect 232682 756 232688 808
rect 232740 796 232746 808
rect 232906 796 232962 800
rect 232740 768 232962 796
rect 233252 796 233280 836
rect 233314 796 233370 800
rect 233252 768 233370 796
rect 233620 796 233648 836
rect 233722 796 233778 800
rect 233620 768 233778 796
rect 232740 756 232746 768
rect 232906 0 232962 768
rect 233314 0 233370 768
rect 233722 0 233778 768
rect 234130 796 234186 800
rect 234338 796 234344 808
rect 234130 768 234344 796
rect 234130 0 234186 768
rect 234338 756 234344 768
rect 234396 756 234402 808
rect 234586 800 234614 836
rect 234538 768 234614 800
rect 234946 796 235002 800
rect 235258 796 235264 808
rect 234946 768 235264 796
rect 234538 0 234594 768
rect 234946 0 235002 768
rect 235258 756 235264 768
rect 235316 756 235322 808
rect 235354 796 235410 800
rect 235534 796 235540 808
rect 235354 768 235540 796
rect 235354 0 235410 768
rect 235534 756 235540 768
rect 235592 756 235598 808
rect 235762 796 235818 800
rect 235994 796 236000 808
rect 235762 768 236000 796
rect 235762 0 235818 768
rect 235994 756 236000 768
rect 236052 756 236058 808
rect 236170 796 236226 800
rect 236288 796 236316 836
rect 236170 768 236316 796
rect 236578 796 236634 800
rect 236822 796 236828 808
rect 236578 768 236828 796
rect 236170 0 236226 768
rect 236578 0 236634 768
rect 236822 756 236828 768
rect 236880 756 236886 808
rect 236986 796 237042 800
rect 237190 796 237196 808
rect 236986 768 237196 796
rect 236986 0 237042 768
rect 237190 756 237196 768
rect 237248 756 237254 808
rect 237394 796 237450 800
rect 237484 796 237512 836
rect 237394 768 237512 796
rect 237802 796 237858 800
rect 238018 796 238024 808
rect 237802 768 238024 796
rect 237394 0 237450 768
rect 237802 0 237858 768
rect 238018 756 238024 768
rect 238076 756 238082 808
rect 238210 796 238266 800
rect 238478 796 238484 808
rect 238210 768 238484 796
rect 238210 0 238266 768
rect 238478 756 238484 768
rect 238536 756 238542 808
rect 238618 660 238674 800
rect 238772 660 238800 836
rect 238618 632 238800 660
rect 239026 796 239082 800
rect 239324 796 239352 904
rect 240134 892 240140 904
rect 240192 892 240198 944
rect 240264 864 240292 972
rect 241882 960 241888 972
rect 241940 960 241946 1012
rect 241992 1000 242020 1040
rect 244200 1040 332600 1068
rect 244200 1000 244228 1040
rect 332594 1028 332600 1040
rect 332652 1028 332658 1080
rect 333054 1028 333060 1080
rect 333112 1068 333118 1080
rect 403710 1068 403716 1080
rect 333112 1040 403716 1068
rect 333112 1028 333118 1040
rect 403710 1028 403716 1040
rect 403768 1028 403774 1080
rect 241992 972 244228 1000
rect 244642 960 244648 1012
rect 244700 1000 244706 1012
rect 336826 1000 336832 1012
rect 244700 972 336832 1000
rect 244700 960 244706 972
rect 336826 960 336832 972
rect 336884 960 336890 1012
rect 335446 932 335452 944
rect 241348 904 335452 932
rect 241238 864 241244 876
rect 240264 836 240364 864
rect 239026 768 239352 796
rect 239434 796 239490 800
rect 239582 796 239588 808
rect 239434 768 239588 796
rect 238618 0 238674 632
rect 239026 0 239082 768
rect 239434 0 239490 768
rect 239582 756 239588 768
rect 239640 756 239646 808
rect 239842 796 239898 800
rect 240042 796 240048 808
rect 239842 768 240048 796
rect 239842 0 239898 768
rect 240042 756 240048 768
rect 240100 756 240106 808
rect 240250 796 240306 800
rect 240336 796 240364 836
rect 240980 836 241244 864
rect 240250 768 240364 796
rect 240658 796 240714 800
rect 240980 796 241008 836
rect 241238 824 241244 836
rect 241296 824 241302 876
rect 240658 768 241008 796
rect 241066 796 241122 800
rect 241348 796 241376 904
rect 335446 892 335452 904
rect 335504 892 335510 944
rect 243262 864 243268 876
rect 243004 836 243268 864
rect 241066 768 241376 796
rect 241474 796 241530 800
rect 241790 796 241796 808
rect 241474 768 241796 796
rect 240250 0 240306 768
rect 240658 0 240714 768
rect 241066 0 241122 768
rect 241474 0 241530 768
rect 241790 756 241796 768
rect 241848 756 241854 808
rect 241882 796 241938 800
rect 242158 796 242164 808
rect 241882 768 242164 796
rect 241882 0 241938 768
rect 242158 756 242164 768
rect 242216 756 242222 808
rect 242290 796 242346 800
rect 242526 796 242532 808
rect 242290 768 242532 796
rect 242290 0 242346 768
rect 242526 756 242532 768
rect 242584 756 242590 808
rect 242698 796 242754 800
rect 243004 796 243032 836
rect 243262 824 243268 836
rect 243320 824 243326 876
rect 244182 864 244188 876
rect 243372 836 244188 864
rect 242698 768 243032 796
rect 243106 796 243162 800
rect 243372 796 243400 836
rect 244182 824 244188 836
rect 244240 824 244246 876
rect 244458 824 244464 876
rect 244516 864 244522 876
rect 334066 864 334072 876
rect 244516 836 334072 864
rect 244516 824 244522 836
rect 334066 824 334072 836
rect 334124 824 334130 876
rect 243106 768 243400 796
rect 243514 796 243570 800
rect 243814 796 243820 808
rect 243514 768 243820 796
rect 242698 0 242754 768
rect 243106 0 243162 768
rect 243514 0 243570 768
rect 243814 756 243820 768
rect 243872 756 243878 808
rect 243922 796 243978 800
rect 244090 796 244096 808
rect 243922 768 244096 796
rect 243922 0 243978 768
rect 244090 756 244096 768
rect 244148 756 244154 808
rect 244330 796 244386 800
rect 244550 796 244556 808
rect 244330 768 244556 796
rect 244330 0 244386 768
rect 244550 756 244556 768
rect 244608 756 244614 808
rect 244738 796 244794 800
rect 244918 796 244924 808
rect 244738 768 244924 796
rect 244738 0 244794 768
rect 244918 756 244924 768
rect 244976 756 244982 808
rect 245146 388 245202 800
rect 245378 388 245384 400
rect 245146 360 245384 388
rect 245146 0 245202 360
rect 245378 348 245384 360
rect 245436 348 245442 400
rect 245554 252 245610 800
rect 245838 252 245844 264
rect 245554 224 245844 252
rect 245554 0 245610 224
rect 245838 212 245844 224
rect 245896 212 245902 264
rect 245962 48 246018 800
rect 249150 552 249156 604
rect 249208 592 249214 604
rect 336458 592 336464 604
rect 249208 564 336464 592
rect 249208 552 249214 564
rect 336458 552 336464 564
rect 336516 552 336522 604
rect 249334 416 249340 468
rect 249392 456 249398 468
rect 339034 456 339040 468
rect 249392 428 339040 456
rect 249392 416 249398 428
rect 339034 416 339040 428
rect 339092 416 339098 468
rect 246114 280 246120 332
rect 246172 320 246178 332
rect 272518 320 272524 332
rect 246172 292 272524 320
rect 246172 280 246178 292
rect 272518 280 272524 292
rect 272576 280 272582 332
rect 246298 212 246304 264
rect 246356 252 246362 264
rect 264606 252 264612 264
rect 246356 224 264612 252
rect 246356 212 246362 224
rect 264606 212 264612 224
rect 264664 212 264670 264
rect 246114 144 246120 196
rect 246172 184 246178 196
rect 287974 184 287980 196
rect 246172 156 287980 184
rect 246172 144 246178 156
rect 287974 144 287980 156
rect 288032 144 288038 196
rect 246390 76 246396 128
rect 246448 116 246454 128
rect 310974 116 310980 128
rect 246448 88 310980 116
rect 246448 76 246454 88
rect 310974 76 310980 88
rect 311032 76 311038 128
rect 341518 48 341524 60
rect 245962 20 341524 48
rect 245962 0 246018 20
rect 341518 8 341524 20
rect 341576 8 341582 60
<< via1 >>
rect 1860 9188 1912 9240
rect 16580 9188 16632 9240
rect 31760 9188 31812 9240
rect 62028 9188 62080 9240
rect 76932 9188 76984 9240
rect 107568 9188 107620 9240
rect 122748 9188 122800 9240
rect 169668 9188 169720 9240
rect 184848 9188 184900 9240
rect 215208 9188 215260 9240
rect 230388 9188 230440 9240
rect 260472 9188 260524 9240
rect 275928 9188 275980 9240
rect 321468 9188 321520 9240
rect 336832 9188 336884 9240
rect 368388 9188 368440 9240
rect 383568 9188 383620 9240
rect 46940 8916 46992 8968
rect 92388 8916 92440 8968
rect 137928 8916 137980 8968
rect 153108 8916 153160 8968
rect 200028 8916 200080 8968
rect 245568 8916 245620 8968
rect 291108 8916 291160 8968
rect 413928 9188 413980 9240
rect 429108 9188 429160 9240
rect 459468 9188 459520 9240
rect 474648 9188 474700 9240
rect 520924 9188 520976 9240
rect 536748 9188 536800 9240
rect 306288 8916 306340 8968
rect 353208 8848 353260 8900
rect 567108 9188 567160 9240
rect 582288 9188 582340 9240
rect 612648 9188 612700 9240
rect 627644 9188 627696 9240
rect 444104 8916 444156 8968
rect 489828 8916 489880 8968
rect 505008 8916 505060 8968
rect 398748 8848 398800 8900
rect 673368 9188 673420 9240
rect 597284 8916 597336 8968
rect 643008 8916 643060 8968
rect 658188 8916 658240 8968
rect 551928 8848 551980 8900
rect 86825 7590 86877 7642
rect 86889 7590 86941 7642
rect 86953 7590 87005 7642
rect 87017 7590 87069 7642
rect 87081 7590 87133 7642
rect 257255 7590 257307 7642
rect 257319 7590 257371 7642
rect 257383 7590 257435 7642
rect 257447 7590 257499 7642
rect 257511 7590 257563 7642
rect 427685 7590 427737 7642
rect 427749 7590 427801 7642
rect 427813 7590 427865 7642
rect 427877 7590 427929 7642
rect 427941 7590 427993 7642
rect 598115 7590 598167 7642
rect 598179 7590 598231 7642
rect 598243 7590 598295 7642
rect 598307 7590 598359 7642
rect 598371 7590 598423 7642
rect 86165 7046 86217 7098
rect 86229 7046 86281 7098
rect 86293 7046 86345 7098
rect 86357 7046 86409 7098
rect 86421 7046 86473 7098
rect 256595 7046 256647 7098
rect 256659 7046 256711 7098
rect 256723 7046 256775 7098
rect 256787 7046 256839 7098
rect 256851 7046 256903 7098
rect 427025 7046 427077 7098
rect 427089 7046 427141 7098
rect 427153 7046 427205 7098
rect 427217 7046 427269 7098
rect 427281 7046 427333 7098
rect 597455 7046 597507 7098
rect 597519 7046 597571 7098
rect 597583 7046 597635 7098
rect 597647 7046 597699 7098
rect 597711 7046 597763 7098
rect 62028 6808 62080 6860
rect 63684 6808 63736 6860
rect 76932 6808 76984 6860
rect 78864 6808 78916 6860
rect 92388 6808 92440 6860
rect 94596 6808 94648 6860
rect 107568 6808 107620 6860
rect 110052 6808 110104 6860
rect 122748 6808 122800 6860
rect 125508 6808 125560 6860
rect 137928 6808 137980 6860
rect 140688 6808 140740 6860
rect 153108 6808 153160 6860
rect 155868 6808 155920 6860
rect 169668 6808 169720 6860
rect 171600 6808 171652 6860
rect 184848 6808 184900 6860
rect 187332 6808 187384 6860
rect 200028 6808 200080 6860
rect 202788 6808 202840 6860
rect 215208 6808 215260 6860
rect 218060 6808 218112 6860
rect 230388 6808 230440 6860
rect 233056 6808 233108 6860
rect 245568 6808 245620 6860
rect 249156 6808 249208 6860
rect 260472 6808 260524 6860
rect 264336 6808 264388 6860
rect 275928 6808 275980 6860
rect 280068 6808 280120 6860
rect 291108 6808 291160 6860
rect 295524 6808 295576 6860
rect 321468 6808 321520 6860
rect 326436 6808 326488 6860
rect 336832 6808 336884 6860
rect 341892 6808 341944 6860
rect 353208 6808 353260 6860
rect 357072 6808 357124 6860
rect 368388 6808 368440 6860
rect 372804 6808 372856 6860
rect 398748 6808 398800 6860
rect 403440 6808 403492 6860
rect 413928 6808 413980 6860
rect 419172 6808 419224 6860
rect 429108 6808 429160 6860
rect 434628 6808 434680 6860
rect 444104 6808 444156 6860
rect 449900 6808 449952 6860
rect 474648 6808 474700 6860
rect 478880 6808 478932 6860
rect 505008 6808 505060 6860
rect 510528 6808 510580 6860
rect 520924 6808 520976 6860
rect 527088 6808 527140 6860
rect 551928 6808 551980 6860
rect 556160 6808 556212 6860
rect 582288 6808 582340 6860
rect 588912 6808 588964 6860
rect 597284 6808 597336 6860
rect 604644 6808 604696 6860
rect 658188 6808 658240 6860
rect 666468 6808 666520 6860
rect 86825 6502 86877 6554
rect 86889 6502 86941 6554
rect 86953 6502 87005 6554
rect 87017 6502 87069 6554
rect 87081 6502 87133 6554
rect 257255 6502 257307 6554
rect 257319 6502 257371 6554
rect 257383 6502 257435 6554
rect 257447 6502 257499 6554
rect 257511 6502 257563 6554
rect 427685 6502 427737 6554
rect 427749 6502 427801 6554
rect 427813 6502 427865 6554
rect 427877 6502 427929 6554
rect 427941 6502 427993 6554
rect 598115 6502 598167 6554
rect 598179 6502 598231 6554
rect 598243 6502 598295 6554
rect 598307 6502 598359 6554
rect 598371 6502 598423 6554
rect 306288 6128 306340 6180
rect 310704 6128 310756 6180
rect 383568 6128 383620 6180
rect 388260 6128 388312 6180
rect 459468 6128 459520 6180
rect 464988 6128 465040 6180
rect 489828 6128 489880 6180
rect 496176 6128 496228 6180
rect 536748 6128 536800 6180
rect 542268 6128 542320 6180
rect 567108 6128 567160 6180
rect 572628 6128 572680 6180
rect 612648 6128 612700 6180
rect 620100 6128 620152 6180
rect 627644 6128 627696 6180
rect 635556 6128 635608 6180
rect 643008 6128 643060 6180
rect 651012 6128 651064 6180
rect 673368 6128 673420 6180
rect 681740 6128 681792 6180
rect 86165 5958 86217 6010
rect 86229 5958 86281 6010
rect 86293 5958 86345 6010
rect 86357 5958 86409 6010
rect 86421 5958 86473 6010
rect 256595 5958 256647 6010
rect 256659 5958 256711 6010
rect 256723 5958 256775 6010
rect 256787 5958 256839 6010
rect 256851 5958 256903 6010
rect 427025 5958 427077 6010
rect 427089 5958 427141 6010
rect 427153 5958 427205 6010
rect 427217 5958 427269 6010
rect 427281 5958 427333 6010
rect 597455 5958 597507 6010
rect 597519 5958 597571 6010
rect 597583 5958 597635 6010
rect 597647 5958 597699 6010
rect 597711 5958 597763 6010
rect 86825 5414 86877 5466
rect 86889 5414 86941 5466
rect 86953 5414 87005 5466
rect 87017 5414 87069 5466
rect 87081 5414 87133 5466
rect 257255 5414 257307 5466
rect 257319 5414 257371 5466
rect 257383 5414 257435 5466
rect 257447 5414 257499 5466
rect 257511 5414 257563 5466
rect 427685 5414 427737 5466
rect 427749 5414 427801 5466
rect 427813 5414 427865 5466
rect 427877 5414 427929 5466
rect 427941 5414 427993 5466
rect 598115 5414 598167 5466
rect 598179 5414 598231 5466
rect 598243 5414 598295 5466
rect 598307 5414 598359 5466
rect 598371 5414 598423 5466
rect 86165 4870 86217 4922
rect 86229 4870 86281 4922
rect 86293 4870 86345 4922
rect 86357 4870 86409 4922
rect 86421 4870 86473 4922
rect 256595 4870 256647 4922
rect 256659 4870 256711 4922
rect 256723 4870 256775 4922
rect 256787 4870 256839 4922
rect 256851 4870 256903 4922
rect 427025 4870 427077 4922
rect 427089 4870 427141 4922
rect 427153 4870 427205 4922
rect 427217 4870 427269 4922
rect 427281 4870 427333 4922
rect 597455 4870 597507 4922
rect 597519 4870 597571 4922
rect 597583 4870 597635 4922
rect 597647 4870 597699 4922
rect 597711 4870 597763 4922
rect 86825 4326 86877 4378
rect 86889 4326 86941 4378
rect 86953 4326 87005 4378
rect 87017 4326 87069 4378
rect 87081 4326 87133 4378
rect 257255 4326 257307 4378
rect 257319 4326 257371 4378
rect 257383 4326 257435 4378
rect 257447 4326 257499 4378
rect 257511 4326 257563 4378
rect 427685 4326 427737 4378
rect 427749 4326 427801 4378
rect 427813 4326 427865 4378
rect 427877 4326 427929 4378
rect 427941 4326 427993 4378
rect 598115 4326 598167 4378
rect 598179 4326 598231 4378
rect 598243 4326 598295 4378
rect 598307 4326 598359 4378
rect 598371 4326 598423 4378
rect 86165 3782 86217 3834
rect 86229 3782 86281 3834
rect 86293 3782 86345 3834
rect 86357 3782 86409 3834
rect 86421 3782 86473 3834
rect 256595 3782 256647 3834
rect 256659 3782 256711 3834
rect 256723 3782 256775 3834
rect 256787 3782 256839 3834
rect 256851 3782 256903 3834
rect 427025 3782 427077 3834
rect 427089 3782 427141 3834
rect 427153 3782 427205 3834
rect 427217 3782 427269 3834
rect 427281 3782 427333 3834
rect 597455 3782 597507 3834
rect 597519 3782 597571 3834
rect 597583 3782 597635 3834
rect 597647 3782 597699 3834
rect 597711 3782 597763 3834
rect 339592 3476 339644 3528
rect 432972 3476 433024 3528
rect 433432 3476 433484 3528
rect 526996 3476 527048 3528
rect 337384 3408 337436 3460
rect 431684 3408 431736 3460
rect 433524 3408 433576 3460
rect 527548 3408 527600 3460
rect 248420 3340 248472 3392
rect 336464 3340 336516 3392
rect 338212 3340 338264 3392
rect 339868 3383 339920 3392
rect 339868 3349 339877 3383
rect 339877 3349 339911 3383
rect 339911 3349 339920 3383
rect 339868 3340 339920 3349
rect 426900 3340 426952 3392
rect 433340 3383 433392 3392
rect 433340 3349 433349 3383
rect 433349 3349 433383 3383
rect 433383 3349 433392 3383
rect 433340 3340 433392 3349
rect 434536 3340 434588 3392
rect 86825 3238 86877 3290
rect 86889 3238 86941 3290
rect 86953 3238 87005 3290
rect 87017 3238 87069 3290
rect 87081 3238 87133 3290
rect 257255 3238 257307 3290
rect 257319 3238 257371 3290
rect 257383 3238 257435 3290
rect 257447 3238 257499 3290
rect 257511 3238 257563 3290
rect 427685 3238 427737 3290
rect 427749 3238 427801 3290
rect 427813 3238 427865 3290
rect 427877 3238 427929 3290
rect 427941 3238 427993 3290
rect 598115 3238 598167 3290
rect 598179 3238 598231 3290
rect 598243 3238 598295 3290
rect 598307 3238 598359 3290
rect 598371 3238 598423 3290
rect 78864 3179 78916 3188
rect 78864 3145 78873 3179
rect 78873 3145 78907 3179
rect 78907 3145 78916 3179
rect 78864 3136 78916 3145
rect 171600 3179 171652 3188
rect 171600 3145 171609 3179
rect 171609 3145 171643 3179
rect 171643 3145 171652 3179
rect 171600 3136 171652 3145
rect 218060 3179 218112 3188
rect 218060 3145 218069 3179
rect 218069 3145 218103 3179
rect 218103 3145 218112 3179
rect 218060 3136 218112 3145
rect 242164 3136 242216 3188
rect 247040 3068 247092 3120
rect 248420 3000 248472 3052
rect 264336 3043 264388 3052
rect 264336 3009 264345 3043
rect 264345 3009 264379 3043
rect 264379 3009 264388 3043
rect 264336 3000 264388 3009
rect 249708 2932 249760 2984
rect 310704 3043 310756 3052
rect 310704 3009 310713 3043
rect 310713 3009 310747 3043
rect 310747 3009 310756 3043
rect 310704 3000 310756 3009
rect 337384 3043 337436 3052
rect 337384 3009 337393 3043
rect 337393 3009 337427 3043
rect 337427 3009 337436 3043
rect 337384 3000 337436 3009
rect 336832 2975 336884 2984
rect 336832 2941 336841 2975
rect 336841 2941 336875 2975
rect 336875 2941 336884 2975
rect 336832 2932 336884 2941
rect 357072 3179 357124 3188
rect 357072 3145 357081 3179
rect 357081 3145 357115 3179
rect 357115 3145 357124 3179
rect 357072 3136 357124 3145
rect 403440 3179 403492 3188
rect 403440 3145 403449 3179
rect 403449 3145 403483 3179
rect 403483 3145 403492 3179
rect 403440 3136 403492 3145
rect 426900 3136 426952 3188
rect 388444 3068 388496 3120
rect 433340 3136 433392 3188
rect 449900 3111 449952 3120
rect 449900 3077 449909 3111
rect 449909 3077 449943 3111
rect 449943 3077 449952 3111
rect 449900 3068 449952 3077
rect 496176 3111 496228 3120
rect 496176 3077 496185 3111
rect 496185 3077 496219 3111
rect 496219 3077 496228 3111
rect 496176 3068 496228 3077
rect 588912 3179 588964 3188
rect 588912 3145 588921 3179
rect 588921 3145 588955 3179
rect 588955 3145 588964 3179
rect 588912 3136 588964 3145
rect 681740 3179 681792 3188
rect 681740 3145 681749 3179
rect 681749 3145 681783 3179
rect 681783 3145 681792 3179
rect 681740 3136 681792 3145
rect 339592 3043 339644 3052
rect 339592 3009 339601 3043
rect 339601 3009 339635 3043
rect 339635 3009 339644 3043
rect 339592 3000 339644 3009
rect 342720 3000 342772 3052
rect 430764 3000 430816 3052
rect 432972 3043 433024 3052
rect 432972 3009 432981 3043
rect 432981 3009 433015 3043
rect 433015 3009 433024 3043
rect 432972 3000 433024 3009
rect 433524 3043 433576 3052
rect 433524 3009 433533 3043
rect 433533 3009 433567 3043
rect 433567 3009 433576 3043
rect 433524 3000 433576 3009
rect 435456 3000 435508 3052
rect 463240 3000 463292 3052
rect 478696 3000 478748 3052
rect 341524 2975 341576 2984
rect 341524 2941 341533 2975
rect 341533 2941 341567 2975
rect 341567 2941 341576 2975
rect 341524 2932 341576 2941
rect 431868 2975 431920 2984
rect 431868 2941 431877 2975
rect 431877 2941 431911 2975
rect 431911 2941 431920 2975
rect 431868 2932 431920 2941
rect 372988 2864 373040 2916
rect 526996 2975 527048 2984
rect 526996 2941 527005 2975
rect 527005 2941 527039 2975
rect 527039 2941 527048 2975
rect 526996 2932 527048 2941
rect 528192 3000 528244 3052
rect 539508 3000 539560 3052
rect 573916 2932 573968 2984
rect 136548 2796 136600 2848
rect 187700 2839 187752 2848
rect 187700 2805 187709 2839
rect 187709 2805 187743 2839
rect 187743 2805 187752 2839
rect 187700 2796 187752 2805
rect 202972 2796 203024 2848
rect 249248 2839 249300 2848
rect 249248 2805 249257 2839
rect 249257 2805 249291 2839
rect 249291 2805 249300 2839
rect 249248 2796 249300 2805
rect 277216 2839 277268 2848
rect 277216 2805 277225 2839
rect 277225 2805 277259 2839
rect 277259 2805 277268 2839
rect 277216 2796 277268 2805
rect 292856 2796 292908 2848
rect 323584 2796 323636 2848
rect 324504 2839 324556 2848
rect 324504 2805 324513 2839
rect 324513 2805 324547 2839
rect 324547 2805 324556 2839
rect 324504 2796 324556 2805
rect 326160 2839 326212 2848
rect 326160 2805 326169 2839
rect 326169 2805 326203 2839
rect 326203 2805 326212 2839
rect 326160 2796 326212 2805
rect 331588 2796 331640 2848
rect 333060 2796 333112 2848
rect 334624 2796 334676 2848
rect 335728 2839 335780 2848
rect 335728 2805 335737 2839
rect 335737 2805 335771 2839
rect 335771 2805 335780 2839
rect 335728 2796 335780 2805
rect 340236 2839 340288 2848
rect 340236 2805 340245 2839
rect 340245 2805 340279 2839
rect 340279 2805 340288 2839
rect 340236 2796 340288 2805
rect 342720 2839 342772 2848
rect 342720 2805 342729 2839
rect 342729 2805 342763 2839
rect 342763 2805 342772 2839
rect 342720 2796 342772 2805
rect 367468 2839 367520 2848
rect 367468 2805 367477 2839
rect 367477 2805 367511 2839
rect 367511 2805 367520 2839
rect 367468 2796 367520 2805
rect 370872 2839 370924 2848
rect 370872 2805 370881 2839
rect 370881 2805 370915 2839
rect 370915 2805 370924 2839
rect 370872 2796 370924 2805
rect 382832 2839 382884 2848
rect 382832 2805 382841 2839
rect 382841 2805 382875 2839
rect 382875 2805 382884 2839
rect 382832 2796 382884 2805
rect 386604 2796 386656 2848
rect 417516 2796 417568 2848
rect 418896 2839 418948 2848
rect 418896 2805 418905 2839
rect 418905 2805 418939 2839
rect 418939 2805 418948 2839
rect 418896 2796 418948 2805
rect 430764 2839 430816 2848
rect 430764 2805 430773 2839
rect 430773 2805 430807 2839
rect 430807 2805 430816 2839
rect 430764 2796 430816 2805
rect 435456 2839 435508 2848
rect 435456 2805 435465 2839
rect 435465 2805 435499 2839
rect 435499 2805 435508 2839
rect 435456 2796 435508 2805
rect 463240 2839 463292 2848
rect 463240 2805 463249 2839
rect 463249 2805 463283 2839
rect 463283 2805 463292 2839
rect 463240 2796 463292 2805
rect 465264 2839 465316 2848
rect 465264 2805 465273 2839
rect 465273 2805 465307 2839
rect 465307 2805 465316 2839
rect 465264 2796 465316 2805
rect 478696 2839 478748 2848
rect 478696 2805 478705 2839
rect 478705 2805 478739 2839
rect 478739 2805 478748 2839
rect 478696 2796 478748 2805
rect 480720 2839 480772 2848
rect 480720 2805 480729 2839
rect 480729 2805 480763 2839
rect 480763 2805 480772 2839
rect 480720 2796 480772 2805
rect 511632 2839 511684 2848
rect 511632 2805 511641 2839
rect 511641 2805 511675 2839
rect 511675 2805 511684 2839
rect 511632 2796 511684 2805
rect 528192 2839 528244 2848
rect 528192 2805 528201 2839
rect 528201 2805 528235 2839
rect 528235 2805 528244 2839
rect 528192 2796 528244 2805
rect 528836 2796 528888 2848
rect 558092 2839 558144 2848
rect 558092 2805 558101 2839
rect 558101 2805 558135 2839
rect 558135 2805 558144 2839
rect 558092 2796 558144 2805
rect 604460 2839 604512 2848
rect 604460 2805 604469 2839
rect 604469 2805 604503 2839
rect 604503 2805 604512 2839
rect 604460 2796 604512 2805
rect 619824 2839 619876 2848
rect 619824 2805 619833 2839
rect 619833 2805 619867 2839
rect 619867 2805 619876 2839
rect 619824 2796 619876 2805
rect 650736 2839 650788 2848
rect 650736 2805 650745 2839
rect 650745 2805 650779 2839
rect 650779 2805 650788 2839
rect 650736 2796 650788 2805
rect 666192 2839 666244 2848
rect 666192 2805 666201 2839
rect 666201 2805 666235 2839
rect 666235 2805 666244 2839
rect 666192 2796 666244 2805
rect 86165 2694 86217 2746
rect 86229 2694 86281 2746
rect 86293 2694 86345 2746
rect 86357 2694 86409 2746
rect 86421 2694 86473 2746
rect 256595 2694 256647 2746
rect 256659 2694 256711 2746
rect 256723 2694 256775 2746
rect 256787 2694 256839 2746
rect 256851 2694 256903 2746
rect 427025 2694 427077 2746
rect 427089 2694 427141 2746
rect 427153 2694 427205 2746
rect 427217 2694 427269 2746
rect 427281 2694 427333 2746
rect 597455 2694 597507 2746
rect 597519 2694 597571 2746
rect 597583 2694 597635 2746
rect 597647 2694 597699 2746
rect 597711 2694 597763 2746
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 16580 2592 16632 2644
rect 46940 2592 46992 2644
rect 63684 2635 63736 2644
rect 63684 2601 63693 2635
rect 63693 2601 63727 2635
rect 63727 2601 63736 2635
rect 63684 2592 63736 2601
rect 94596 2635 94648 2644
rect 94596 2601 94605 2635
rect 94605 2601 94639 2635
rect 94639 2601 94648 2635
rect 94596 2592 94648 2601
rect 97356 2592 97408 2644
rect 31760 2388 31812 2440
rect 78864 2388 78916 2440
rect 95332 2388 95384 2440
rect 96804 2363 96856 2372
rect 96804 2329 96813 2363
rect 96813 2329 96847 2363
rect 96847 2329 96856 2363
rect 96804 2320 96856 2329
rect 97356 2431 97408 2440
rect 97356 2397 97365 2431
rect 97365 2397 97399 2431
rect 97399 2397 97408 2431
rect 97356 2388 97408 2397
rect 110696 2388 110748 2440
rect 113456 2388 113508 2440
rect 125508 2431 125560 2440
rect 125508 2397 125517 2431
rect 125517 2397 125551 2431
rect 125551 2397 125560 2431
rect 125508 2388 125560 2397
rect 136548 2431 136600 2440
rect 136548 2397 136557 2431
rect 136557 2397 136591 2431
rect 136591 2397 136600 2431
rect 136548 2388 136600 2397
rect 2596 2295 2648 2304
rect 2596 2261 2605 2295
rect 2605 2261 2639 2295
rect 2639 2261 2648 2295
rect 2596 2252 2648 2261
rect 18052 2295 18104 2304
rect 18052 2261 18061 2295
rect 18061 2261 18095 2295
rect 18095 2261 18104 2295
rect 18052 2252 18104 2261
rect 79140 2295 79192 2304
rect 79140 2261 79149 2295
rect 79149 2261 79183 2295
rect 79183 2261 79192 2295
rect 79140 2252 79192 2261
rect 95332 2295 95384 2304
rect 95332 2261 95341 2295
rect 95341 2261 95375 2295
rect 95375 2261 95384 2295
rect 95332 2252 95384 2261
rect 110052 2295 110104 2304
rect 110052 2261 110061 2295
rect 110061 2261 110095 2295
rect 110095 2261 110104 2295
rect 110052 2252 110104 2261
rect 110696 2295 110748 2304
rect 110696 2261 110705 2295
rect 110705 2261 110739 2295
rect 110739 2261 110748 2295
rect 110696 2252 110748 2261
rect 112260 2363 112312 2372
rect 112260 2329 112269 2363
rect 112269 2329 112303 2363
rect 112303 2329 112312 2363
rect 112260 2320 112312 2329
rect 113456 2295 113508 2304
rect 113456 2261 113465 2295
rect 113465 2261 113499 2295
rect 113499 2261 113508 2295
rect 113456 2252 113508 2261
rect 125692 2295 125744 2304
rect 125692 2261 125701 2295
rect 125701 2261 125735 2295
rect 125735 2261 125744 2295
rect 125692 2252 125744 2261
rect 135996 2363 136048 2372
rect 135996 2329 136005 2363
rect 136005 2329 136039 2363
rect 136039 2329 136048 2363
rect 135996 2320 136048 2329
rect 136824 2363 136876 2372
rect 136824 2329 136833 2363
rect 136833 2329 136867 2363
rect 136867 2329 136876 2363
rect 136824 2320 136876 2329
rect 138112 2431 138164 2440
rect 138112 2397 138121 2431
rect 138121 2397 138155 2431
rect 138155 2397 138164 2431
rect 138112 2388 138164 2397
rect 140688 2524 140740 2576
rect 155868 2524 155920 2576
rect 138388 2456 138440 2508
rect 187332 2635 187384 2644
rect 187332 2601 187341 2635
rect 187341 2601 187375 2635
rect 187375 2601 187384 2635
rect 187332 2592 187384 2601
rect 202788 2635 202840 2644
rect 202788 2601 202797 2635
rect 202797 2601 202831 2635
rect 202831 2601 202840 2635
rect 202788 2592 202840 2601
rect 233056 2592 233108 2644
rect 244280 2592 244332 2644
rect 248052 2635 248104 2644
rect 248052 2601 248061 2635
rect 248061 2601 248095 2635
rect 248095 2601 248104 2635
rect 248052 2592 248104 2601
rect 249156 2635 249208 2644
rect 249156 2601 249165 2635
rect 249165 2601 249199 2635
rect 249199 2601 249208 2635
rect 249156 2592 249208 2601
rect 273352 2592 273404 2644
rect 218244 2567 218296 2576
rect 218244 2533 218253 2567
rect 218253 2533 218287 2567
rect 218287 2533 218296 2567
rect 218244 2524 218296 2533
rect 238024 2524 238076 2576
rect 247040 2524 247092 2576
rect 249248 2524 249300 2576
rect 295524 2635 295576 2644
rect 295524 2601 295533 2635
rect 295533 2601 295567 2635
rect 295567 2601 295576 2635
rect 295524 2592 295576 2601
rect 367468 2592 367520 2644
rect 141700 2388 141752 2440
rect 157156 2388 157208 2440
rect 171600 2388 171652 2440
rect 189540 2431 189592 2440
rect 138204 2252 138256 2304
rect 138296 2295 138348 2304
rect 138296 2261 138305 2295
rect 138305 2261 138339 2295
rect 138339 2261 138348 2295
rect 138296 2252 138348 2261
rect 141700 2295 141752 2304
rect 141700 2261 141709 2295
rect 141709 2261 141743 2295
rect 141743 2261 141752 2295
rect 141700 2252 141752 2261
rect 144368 2295 144420 2304
rect 144368 2261 144377 2295
rect 144377 2261 144411 2295
rect 144411 2261 144420 2295
rect 144368 2252 144420 2261
rect 157156 2295 157208 2304
rect 157156 2261 157165 2295
rect 157165 2261 157199 2295
rect 157199 2261 157208 2295
rect 157156 2252 157208 2261
rect 159824 2295 159876 2304
rect 159824 2261 159833 2295
rect 159833 2261 159867 2295
rect 159867 2261 159876 2295
rect 159824 2252 159876 2261
rect 171876 2295 171928 2304
rect 171876 2261 171885 2295
rect 171885 2261 171919 2295
rect 171919 2261 171928 2295
rect 171876 2252 171928 2261
rect 189540 2397 189549 2431
rect 189549 2397 189583 2431
rect 189583 2397 189592 2431
rect 189540 2388 189592 2397
rect 191380 2388 191432 2440
rect 188620 2363 188672 2372
rect 188620 2329 188629 2363
rect 188629 2329 188663 2363
rect 188663 2329 188672 2363
rect 188620 2320 188672 2329
rect 202972 2431 203024 2440
rect 202972 2397 202981 2431
rect 202981 2397 203015 2431
rect 203015 2397 203024 2431
rect 202972 2388 203024 2397
rect 187700 2252 187752 2304
rect 203892 2363 203944 2372
rect 203892 2329 203901 2363
rect 203901 2329 203935 2363
rect 203935 2329 203944 2363
rect 203892 2320 203944 2329
rect 191380 2295 191432 2304
rect 191380 2261 191389 2295
rect 191389 2261 191423 2295
rect 191423 2261 191432 2295
rect 191380 2252 191432 2261
rect 205916 2363 205968 2372
rect 205916 2329 205925 2363
rect 205925 2329 205959 2363
rect 205959 2329 205968 2363
rect 205916 2320 205968 2329
rect 228180 2456 228232 2508
rect 240140 2456 240192 2508
rect 218060 2388 218112 2440
rect 232688 2320 232740 2372
rect 230664 2252 230716 2304
rect 234344 2295 234396 2304
rect 234344 2261 234353 2295
rect 234353 2261 234387 2295
rect 234387 2261 234396 2295
rect 234344 2252 234396 2261
rect 239588 2252 239640 2304
rect 248052 2388 248104 2440
rect 250444 2320 250496 2372
rect 264336 2388 264388 2440
rect 273352 2431 273404 2440
rect 273352 2397 273361 2431
rect 273361 2397 273395 2431
rect 273395 2397 273404 2431
rect 273352 2388 273404 2397
rect 276020 2388 276072 2440
rect 277216 2388 277268 2440
rect 275560 2363 275612 2372
rect 275560 2329 275569 2363
rect 275569 2329 275603 2363
rect 275603 2329 275612 2363
rect 275560 2320 275612 2329
rect 277676 2363 277728 2372
rect 277676 2329 277685 2363
rect 277685 2329 277719 2363
rect 277719 2329 277728 2363
rect 277676 2320 277728 2329
rect 264612 2295 264664 2304
rect 264612 2261 264621 2295
rect 264621 2261 264655 2295
rect 264655 2261 264664 2295
rect 264612 2252 264664 2261
rect 272524 2295 272576 2304
rect 272524 2261 272533 2295
rect 272533 2261 272567 2295
rect 272567 2261 272576 2295
rect 272524 2252 272576 2261
rect 274732 2295 274784 2304
rect 274732 2261 274741 2295
rect 274741 2261 274775 2295
rect 274775 2261 274784 2295
rect 274732 2252 274784 2261
rect 278964 2295 279016 2304
rect 278964 2261 278973 2295
rect 278973 2261 279007 2295
rect 279007 2261 279016 2295
rect 278964 2252 279016 2261
rect 280068 2295 280120 2304
rect 280068 2261 280077 2295
rect 280077 2261 280111 2295
rect 280111 2261 280120 2295
rect 280068 2252 280120 2261
rect 287980 2295 288032 2304
rect 287980 2261 287989 2295
rect 287989 2261 288023 2295
rect 288023 2261 288032 2295
rect 287980 2252 288032 2261
rect 290188 2363 290240 2372
rect 290188 2329 290197 2363
rect 290197 2329 290231 2363
rect 290231 2329 290240 2363
rect 290188 2320 290240 2329
rect 290924 2363 290976 2372
rect 290924 2329 290933 2363
rect 290933 2329 290967 2363
rect 290967 2329 290976 2363
rect 290924 2320 290976 2329
rect 295800 2456 295852 2508
rect 292856 2431 292908 2440
rect 292856 2397 292865 2431
rect 292865 2397 292899 2431
rect 292899 2397 292908 2431
rect 292856 2388 292908 2397
rect 293408 2363 293460 2372
rect 293408 2329 293417 2363
rect 293417 2329 293451 2363
rect 293451 2329 293460 2363
rect 293408 2320 293460 2329
rect 294420 2431 294472 2440
rect 294420 2397 294429 2431
rect 294429 2397 294463 2431
rect 294463 2397 294472 2431
rect 294420 2388 294472 2397
rect 310704 2388 310756 2440
rect 320916 2388 320968 2440
rect 323584 2431 323636 2440
rect 323584 2397 323593 2431
rect 323593 2397 323627 2431
rect 323627 2397 323636 2431
rect 323584 2388 323636 2397
rect 295616 2252 295668 2304
rect 310980 2295 311032 2304
rect 310980 2261 310989 2295
rect 310989 2261 311023 2295
rect 311023 2261 311032 2295
rect 310980 2252 311032 2261
rect 320916 2295 320968 2304
rect 320916 2261 320925 2295
rect 320925 2261 320959 2295
rect 320959 2261 320968 2295
rect 320916 2252 320968 2261
rect 322112 2363 322164 2372
rect 322112 2329 322121 2363
rect 322121 2329 322155 2363
rect 322155 2329 322164 2363
rect 322112 2320 322164 2329
rect 324504 2388 324556 2440
rect 326160 2388 326212 2440
rect 331588 2431 331640 2440
rect 331588 2397 331597 2431
rect 331597 2397 331631 2431
rect 331631 2397 331640 2431
rect 331588 2388 331640 2397
rect 333060 2431 333112 2440
rect 333060 2397 333069 2431
rect 333069 2397 333103 2431
rect 333103 2397 333112 2431
rect 333060 2388 333112 2397
rect 334624 2431 334676 2440
rect 334624 2397 334633 2431
rect 334633 2397 334667 2431
rect 334667 2397 334676 2431
rect 334624 2388 334676 2397
rect 335728 2431 335780 2440
rect 335728 2397 335737 2431
rect 335737 2397 335771 2431
rect 335771 2397 335780 2431
rect 335728 2388 335780 2397
rect 336464 2431 336516 2440
rect 336464 2397 336473 2431
rect 336473 2397 336507 2431
rect 336507 2397 336516 2431
rect 336464 2388 336516 2397
rect 338212 2431 338264 2440
rect 338212 2397 338221 2431
rect 338221 2397 338255 2431
rect 338255 2397 338264 2431
rect 338212 2388 338264 2397
rect 339868 2388 339920 2440
rect 340236 2431 340288 2440
rect 340236 2397 340245 2431
rect 340245 2397 340279 2431
rect 340279 2397 340288 2431
rect 340236 2388 340288 2397
rect 324136 2363 324188 2372
rect 324136 2329 324145 2363
rect 324145 2329 324179 2363
rect 324179 2329 324188 2363
rect 324136 2320 324188 2329
rect 325332 2363 325384 2372
rect 325332 2329 325341 2363
rect 325341 2329 325375 2363
rect 325375 2329 325384 2363
rect 325332 2320 325384 2329
rect 331312 2363 331364 2372
rect 331312 2329 331321 2363
rect 331321 2329 331355 2363
rect 331355 2329 331364 2363
rect 331312 2320 331364 2329
rect 332600 2363 332652 2372
rect 332600 2329 332609 2363
rect 332609 2329 332643 2363
rect 332643 2329 332652 2363
rect 332600 2320 332652 2329
rect 334072 2363 334124 2372
rect 334072 2329 334081 2363
rect 334081 2329 334115 2363
rect 334115 2329 334124 2363
rect 334072 2320 334124 2329
rect 335452 2363 335504 2372
rect 335452 2329 335461 2363
rect 335461 2329 335495 2363
rect 335495 2329 335504 2363
rect 335452 2320 335504 2329
rect 337016 2363 337068 2372
rect 337016 2329 337025 2363
rect 337025 2329 337059 2363
rect 337059 2329 337068 2363
rect 337016 2320 337068 2329
rect 337660 2363 337712 2372
rect 337660 2329 337669 2363
rect 337669 2329 337703 2363
rect 337703 2329 337712 2363
rect 337660 2320 337712 2329
rect 339040 2363 339092 2372
rect 339040 2329 339049 2363
rect 339049 2329 339083 2363
rect 339083 2329 339092 2363
rect 339040 2320 339092 2329
rect 340788 2363 340840 2372
rect 340788 2329 340797 2363
rect 340797 2329 340831 2363
rect 340831 2329 340840 2363
rect 340788 2320 340840 2329
rect 357072 2388 357124 2440
rect 367468 2388 367520 2440
rect 368296 2363 368348 2372
rect 368296 2329 368305 2363
rect 368305 2329 368339 2363
rect 368339 2329 368348 2363
rect 368296 2320 368348 2329
rect 370320 2388 370372 2440
rect 370872 2388 370924 2440
rect 370412 2363 370464 2372
rect 370412 2329 370421 2363
rect 370421 2329 370455 2363
rect 370455 2329 370464 2363
rect 370412 2320 370464 2329
rect 465264 2592 465316 2644
rect 478880 2592 478932 2644
rect 510528 2592 510580 2644
rect 372804 2567 372856 2576
rect 372804 2533 372813 2567
rect 372813 2533 372847 2567
rect 372847 2533 372856 2567
rect 372804 2524 372856 2533
rect 388260 2567 388312 2576
rect 388260 2533 388269 2567
rect 388269 2533 388303 2567
rect 388303 2533 388312 2567
rect 388260 2524 388312 2533
rect 478696 2524 478748 2576
rect 372988 2431 373040 2440
rect 372988 2397 372997 2431
rect 372997 2397 373031 2431
rect 373031 2397 373040 2431
rect 372988 2388 373040 2397
rect 382832 2320 382884 2372
rect 383660 2363 383712 2372
rect 383660 2329 383669 2363
rect 383669 2329 383703 2363
rect 383703 2329 383712 2363
rect 383660 2320 383712 2329
rect 386604 2431 386656 2440
rect 386604 2397 386613 2431
rect 386613 2397 386647 2431
rect 386647 2397 386656 2431
rect 386604 2388 386656 2397
rect 388444 2431 388496 2440
rect 388444 2397 388453 2431
rect 388453 2397 388487 2431
rect 388487 2397 388496 2431
rect 388444 2388 388496 2397
rect 403440 2388 403492 2440
rect 387156 2363 387208 2372
rect 387156 2329 387165 2363
rect 387165 2329 387199 2363
rect 387199 2329 387208 2363
rect 387156 2320 387208 2329
rect 417516 2431 417568 2440
rect 417516 2397 417525 2431
rect 417525 2397 417559 2431
rect 417559 2397 417568 2431
rect 417516 2388 417568 2397
rect 418896 2388 418948 2440
rect 416780 2363 416832 2372
rect 416780 2329 416789 2363
rect 416789 2329 416823 2363
rect 416823 2329 416832 2363
rect 416780 2320 416832 2329
rect 428188 2363 428240 2372
rect 428188 2329 428197 2363
rect 428197 2329 428231 2363
rect 428231 2329 428240 2363
rect 428188 2320 428240 2329
rect 429752 2363 429804 2372
rect 429752 2329 429761 2363
rect 429761 2329 429795 2363
rect 429795 2329 429804 2363
rect 429752 2320 429804 2329
rect 431684 2431 431736 2440
rect 431684 2397 431693 2431
rect 431693 2397 431727 2431
rect 431727 2397 431736 2431
rect 431684 2388 431736 2397
rect 433340 2388 433392 2440
rect 433432 2431 433484 2440
rect 433432 2397 433441 2431
rect 433441 2397 433475 2431
rect 433475 2397 433484 2431
rect 433432 2388 433484 2397
rect 434536 2388 434588 2440
rect 432880 2363 432932 2372
rect 432880 2329 432889 2363
rect 432889 2329 432923 2363
rect 432923 2329 432932 2363
rect 432880 2320 432932 2329
rect 435364 2363 435416 2372
rect 435364 2329 435373 2363
rect 435373 2329 435407 2363
rect 435407 2329 435416 2363
rect 435364 2320 435416 2329
rect 449900 2320 449952 2372
rect 461860 2388 461912 2440
rect 463332 2363 463384 2372
rect 463332 2329 463341 2363
rect 463341 2329 463375 2363
rect 463375 2329 463384 2363
rect 463332 2320 463384 2329
rect 465264 2388 465316 2440
rect 477316 2388 477368 2440
rect 480720 2388 480772 2440
rect 496176 2388 496228 2440
rect 509700 2431 509752 2440
rect 509700 2397 509709 2431
rect 509709 2397 509743 2431
rect 509743 2397 509752 2431
rect 509700 2388 509752 2397
rect 604460 2592 604512 2644
rect 604644 2635 604696 2644
rect 604644 2601 604653 2635
rect 604653 2601 604687 2635
rect 604687 2601 604696 2635
rect 604644 2592 604696 2601
rect 620100 2635 620152 2644
rect 620100 2601 620109 2635
rect 620109 2601 620143 2635
rect 620143 2601 620152 2635
rect 620100 2592 620152 2601
rect 625436 2592 625488 2644
rect 525064 2567 525116 2576
rect 525064 2533 525073 2567
rect 525073 2533 525107 2567
rect 525107 2533 525116 2567
rect 525064 2524 525116 2533
rect 511632 2388 511684 2440
rect 525064 2388 525116 2440
rect 619824 2524 619876 2576
rect 527548 2431 527600 2440
rect 527548 2397 527557 2431
rect 527557 2397 527591 2431
rect 527591 2397 527600 2431
rect 527548 2388 527600 2397
rect 528836 2431 528888 2440
rect 528836 2397 528845 2431
rect 528845 2397 528879 2431
rect 528879 2397 528888 2431
rect 528836 2388 528888 2397
rect 326436 2295 326488 2304
rect 326436 2261 326445 2295
rect 326445 2261 326479 2295
rect 326479 2261 326488 2295
rect 326436 2252 326488 2261
rect 341892 2295 341944 2304
rect 341892 2261 341901 2295
rect 341901 2261 341935 2295
rect 341935 2261 341944 2295
rect 341892 2252 341944 2261
rect 357348 2295 357400 2304
rect 357348 2261 357357 2295
rect 357357 2261 357391 2295
rect 357391 2261 357400 2295
rect 357348 2252 357400 2261
rect 369124 2295 369176 2304
rect 369124 2261 369133 2295
rect 369133 2261 369167 2295
rect 369167 2261 369176 2295
rect 369124 2252 369176 2261
rect 384580 2295 384632 2304
rect 384580 2261 384589 2295
rect 384589 2261 384623 2295
rect 384623 2261 384632 2295
rect 384580 2252 384632 2261
rect 403716 2295 403768 2304
rect 403716 2261 403725 2295
rect 403725 2261 403759 2295
rect 403759 2261 403768 2295
rect 403716 2252 403768 2261
rect 415492 2295 415544 2304
rect 415492 2261 415501 2295
rect 415501 2261 415535 2295
rect 415535 2261 415544 2295
rect 415492 2252 415544 2261
rect 419172 2295 419224 2304
rect 419172 2261 419181 2295
rect 419181 2261 419215 2295
rect 419215 2261 419224 2295
rect 419172 2252 419224 2261
rect 429108 2295 429160 2304
rect 429108 2261 429117 2295
rect 429117 2261 429151 2295
rect 429151 2261 429160 2295
rect 429108 2252 429160 2261
rect 430948 2295 431000 2304
rect 430948 2261 430957 2295
rect 430957 2261 430991 2295
rect 430991 2261 431000 2295
rect 430948 2252 431000 2261
rect 434628 2295 434680 2304
rect 434628 2261 434637 2295
rect 434637 2261 434671 2295
rect 434671 2261 434680 2295
rect 434628 2252 434680 2261
rect 436836 2295 436888 2304
rect 436836 2261 436845 2295
rect 436845 2261 436879 2295
rect 436879 2261 436888 2295
rect 436836 2252 436888 2261
rect 450084 2295 450136 2304
rect 450084 2261 450093 2295
rect 450093 2261 450127 2295
rect 450127 2261 450136 2295
rect 450084 2252 450136 2261
rect 461860 2295 461912 2304
rect 461860 2261 461869 2295
rect 461869 2261 461903 2295
rect 461903 2261 461912 2295
rect 461860 2252 461912 2261
rect 464988 2252 465040 2304
rect 477316 2295 477368 2304
rect 477316 2261 477325 2295
rect 477325 2261 477359 2295
rect 477359 2261 477368 2295
rect 477316 2252 477368 2261
rect 496452 2295 496504 2304
rect 496452 2261 496461 2295
rect 496461 2261 496495 2295
rect 496495 2261 496504 2295
rect 496452 2252 496504 2261
rect 528284 2363 528336 2372
rect 528284 2329 528293 2363
rect 528293 2329 528327 2363
rect 528327 2329 528336 2363
rect 528284 2320 528336 2329
rect 529756 2363 529808 2372
rect 529756 2329 529765 2363
rect 529765 2329 529799 2363
rect 529799 2329 529808 2363
rect 529756 2320 529808 2329
rect 542268 2388 542320 2440
rect 558092 2388 558144 2440
rect 573916 2431 573968 2440
rect 573916 2397 573925 2431
rect 573925 2397 573959 2431
rect 573959 2397 573968 2431
rect 573916 2388 573968 2397
rect 588912 2388 588964 2440
rect 604460 2388 604512 2440
rect 619824 2388 619876 2440
rect 511632 2252 511684 2304
rect 527088 2252 527140 2304
rect 530952 2295 531004 2304
rect 530952 2261 530961 2295
rect 530961 2261 530995 2295
rect 530995 2261 531004 2295
rect 530952 2252 531004 2261
rect 539508 2252 539560 2304
rect 555332 2295 555384 2304
rect 555332 2261 555341 2295
rect 555341 2261 555375 2295
rect 555375 2261 555384 2295
rect 555332 2252 555384 2261
rect 556160 2252 556212 2304
rect 572628 2252 572680 2304
rect 589188 2295 589240 2304
rect 589188 2261 589197 2295
rect 589197 2261 589231 2295
rect 589231 2261 589240 2295
rect 589188 2252 589240 2261
rect 623044 2363 623096 2372
rect 623044 2329 623053 2363
rect 623053 2329 623087 2363
rect 623087 2329 623096 2363
rect 623044 2320 623096 2329
rect 651012 2567 651064 2576
rect 651012 2533 651021 2567
rect 651021 2533 651055 2567
rect 651055 2533 651064 2567
rect 651012 2524 651064 2533
rect 666468 2567 666520 2576
rect 666468 2533 666477 2567
rect 666477 2533 666511 2567
rect 666511 2533 666520 2567
rect 666468 2524 666520 2533
rect 666192 2456 666244 2508
rect 625436 2431 625488 2440
rect 625436 2397 625445 2431
rect 625445 2397 625479 2431
rect 625479 2397 625488 2431
rect 625436 2388 625488 2397
rect 635556 2431 635608 2440
rect 635556 2397 635565 2431
rect 635565 2397 635599 2431
rect 635599 2397 635608 2431
rect 635556 2388 635608 2397
rect 624884 2363 624936 2372
rect 624884 2329 624893 2363
rect 624893 2329 624927 2363
rect 624927 2329 624936 2363
rect 624884 2320 624936 2329
rect 650736 2320 650788 2372
rect 681740 2388 681792 2440
rect 86825 2150 86877 2202
rect 86889 2150 86941 2202
rect 86953 2150 87005 2202
rect 87017 2150 87069 2202
rect 87081 2150 87133 2202
rect 257255 2150 257307 2202
rect 257319 2150 257371 2202
rect 257383 2150 257435 2202
rect 257447 2150 257499 2202
rect 257511 2150 257563 2202
rect 427685 2150 427737 2202
rect 427749 2150 427801 2202
rect 427813 2150 427865 2202
rect 427877 2150 427929 2202
rect 427941 2150 427993 2202
rect 598115 2150 598167 2202
rect 598179 2150 598231 2202
rect 598243 2150 598295 2202
rect 598307 2150 598359 2202
rect 598371 2150 598423 2202
rect 2596 2048 2648 2100
rect 96804 2048 96856 2100
rect 110696 2048 110748 2100
rect 203892 2048 203944 2100
rect 218244 2048 218296 2100
rect 231768 2048 231820 2100
rect 243268 2048 243320 2100
rect 274732 2048 274784 2100
rect 290924 2048 290976 2100
rect 384580 2048 384632 2100
rect 416780 2048 416832 2100
rect 509700 2048 509752 2100
rect 528192 2048 528244 2100
rect 589188 2048 589240 2100
rect 79140 1980 79192 2032
rect 136548 1980 136600 2032
rect 235540 1980 235592 2032
rect 278964 1980 279016 2032
rect 322112 1980 322164 2032
rect 415492 1980 415544 2032
rect 429108 1980 429160 2032
rect 450084 1980 450136 2032
rect 463332 1980 463384 2032
rect 555332 1980 555384 2032
rect 18052 1912 18104 1964
rect 112260 1912 112312 1964
rect 125692 1912 125744 1964
rect 138112 1912 138164 1964
rect 236000 1912 236052 1964
rect 244188 1912 244240 1964
rect 244372 1912 244424 1964
rect 290188 1912 290240 1964
rect 293408 1912 293460 1964
rect 386604 1912 386656 1964
rect 530952 1912 531004 1964
rect 624884 1912 624936 1964
rect 238484 1844 238536 1896
rect 249708 1844 249760 1896
rect 277676 1844 277728 1896
rect 370320 1844 370372 1896
rect 370412 1844 370464 1896
rect 463240 1844 463292 1896
rect 528836 1844 528888 1896
rect 623044 1844 623096 1896
rect 95332 1776 95384 1828
rect 188620 1776 188672 1828
rect 244096 1776 244148 1828
rect 320916 1776 320968 1828
rect 342720 1776 342772 1828
rect 435364 1776 435416 1828
rect 436836 1776 436888 1828
rect 529756 1776 529808 1828
rect 113456 1708 113508 1760
rect 205916 1708 205968 1760
rect 244188 1708 244240 1760
rect 294420 1708 294472 1760
rect 331588 1708 331640 1760
rect 357348 1708 357400 1760
rect 430948 1708 431000 1760
rect 496452 1708 496504 1760
rect 241520 1640 241572 1692
rect 189540 1300 189592 1352
rect 227260 1300 227312 1352
rect 232228 1436 232280 1488
rect 235264 1436 235316 1488
rect 246304 1572 246356 1624
rect 246488 1640 246540 1692
rect 276020 1640 276072 1692
rect 324136 1640 324188 1692
rect 417516 1640 417568 1692
rect 435456 1640 435508 1692
rect 528284 1640 528336 1692
rect 243544 1504 243596 1556
rect 244280 1504 244332 1556
rect 275560 1572 275612 1624
rect 369124 1572 369176 1624
rect 383660 1572 383712 1624
rect 477316 1572 477368 1624
rect 292856 1504 292908 1556
rect 325332 1504 325384 1556
rect 418896 1504 418948 1556
rect 241888 1436 241940 1488
rect 246488 1436 246540 1488
rect 250444 1436 250496 1488
rect 340236 1436 340288 1488
rect 387156 1436 387208 1488
rect 480720 1436 480772 1488
rect 231768 1368 231820 1420
rect 171876 1232 171928 1284
rect 227812 1300 227864 1352
rect 159824 1164 159876 1216
rect 229376 1232 229428 1284
rect 229468 1232 229520 1284
rect 231952 1232 232004 1284
rect 227628 1164 227680 1216
rect 157156 1096 157208 1148
rect 227444 1096 227496 1148
rect 227720 1096 227772 1148
rect 144368 1028 144420 1080
rect 141700 960 141752 1012
rect 135996 892 136048 944
rect 138296 824 138348 876
rect 224224 1028 224276 1080
rect 228640 1028 228692 1080
rect 228732 1028 228784 1080
rect 224316 960 224368 1012
rect 227260 824 227312 876
rect 228732 824 228784 876
rect 227628 756 227680 808
rect 224132 688 224184 740
rect 227720 620 227772 672
rect 136824 212 136876 264
rect 224132 212 224184 264
rect 202972 144 203024 196
rect 227720 144 227772 196
rect 191380 8 191432 60
rect 228180 756 228232 808
rect 228640 756 228692 808
rect 232228 1096 232280 1148
rect 237196 1300 237248 1352
rect 244004 1368 244056 1420
rect 244832 1368 244884 1420
rect 323584 1368 323636 1420
rect 340788 1368 340840 1420
rect 434536 1368 434588 1420
rect 243544 1232 243596 1284
rect 244556 1300 244608 1352
rect 249432 1300 249484 1352
rect 229376 756 229428 808
rect 230664 756 230716 808
rect 239956 1164 240008 1216
rect 240048 1164 240100 1216
rect 243636 1164 243688 1216
rect 243912 1232 243964 1284
rect 244280 1164 244332 1216
rect 242072 1096 242124 1148
rect 242532 1096 242584 1148
rect 244004 1096 244056 1148
rect 244832 1232 244884 1284
rect 338212 1300 338264 1352
rect 432880 1300 432932 1352
rect 244740 1164 244792 1216
rect 249156 1164 249208 1216
rect 331312 1232 331364 1284
rect 335728 1232 335780 1284
rect 429752 1232 429804 1284
rect 244832 1096 244884 1148
rect 244924 1096 244976 1148
rect 249340 1096 249392 1148
rect 334624 1164 334676 1216
rect 428188 1164 428240 1216
rect 337660 1096 337712 1148
rect 368296 1096 368348 1148
rect 461860 1096 461912 1148
rect 231952 620 232004 672
rect 232688 756 232740 808
rect 234344 756 234396 808
rect 235264 756 235316 808
rect 235540 756 235592 808
rect 236000 756 236052 808
rect 236828 756 236880 808
rect 237196 756 237248 808
rect 238024 756 238076 808
rect 238484 756 238536 808
rect 240140 892 240192 944
rect 241888 960 241940 1012
rect 332600 1028 332652 1080
rect 333060 1028 333112 1080
rect 403716 1028 403768 1080
rect 244648 960 244700 1012
rect 336832 960 336884 1012
rect 239588 756 239640 808
rect 240048 756 240100 808
rect 241244 824 241296 876
rect 335452 892 335504 944
rect 241796 756 241848 808
rect 242164 756 242216 808
rect 242532 756 242584 808
rect 243268 824 243320 876
rect 244188 824 244240 876
rect 244464 824 244516 876
rect 334072 824 334124 876
rect 243820 756 243872 808
rect 244096 756 244148 808
rect 244556 756 244608 808
rect 244924 756 244976 808
rect 245384 348 245436 400
rect 245844 212 245896 264
rect 249156 552 249208 604
rect 336464 552 336516 604
rect 249340 416 249392 468
rect 339040 416 339092 468
rect 246120 280 246172 332
rect 272524 280 272576 332
rect 246304 212 246356 264
rect 264612 212 264664 264
rect 246120 144 246172 196
rect 287980 144 288032 196
rect 246396 76 246448 128
rect 310980 76 311032 128
rect 341524 8 341576 60
<< metal2 >>
rect -1076 9784 -756 9796
rect -1076 9728 -1064 9784
rect -1008 9728 -984 9784
rect -928 9728 -904 9784
rect -848 9728 -824 9784
rect -768 9728 -756 9784
rect -1076 9704 -756 9728
rect -1076 9648 -1064 9704
rect -1008 9648 -984 9704
rect -928 9648 -904 9704
rect -848 9648 -824 9704
rect -768 9648 -756 9704
rect -1076 9624 -756 9648
rect -1076 9568 -1064 9624
rect -1008 9568 -984 9624
rect -928 9568 -904 9624
rect -848 9568 -824 9624
rect -768 9568 -756 9624
rect -1076 9544 -756 9568
rect -1076 9488 -1064 9544
rect -1008 9488 -984 9544
rect -928 9488 -904 9544
rect -848 9488 -824 9544
rect -768 9488 -756 9544
rect -1076 7740 -756 9488
rect 1860 9240 1912 9246
rect 1860 9182 1912 9188
rect 16580 9240 16632 9246
rect 16580 9182 16632 9188
rect 31760 9240 31812 9246
rect 31760 9182 31812 9188
rect 62028 9240 62080 9246
rect 62028 9182 62080 9188
rect 76932 9240 76984 9246
rect 76932 9182 76984 9188
rect -1076 7684 -1064 7740
rect -1008 7684 -984 7740
rect -928 7684 -904 7740
rect -848 7684 -824 7740
rect -768 7684 -756 7740
rect -1076 7660 -756 7684
rect -1076 7604 -1064 7660
rect -1008 7604 -984 7660
rect -928 7604 -904 7660
rect -848 7604 -824 7660
rect -768 7604 -756 7660
rect -1076 7580 -756 7604
rect -1076 7524 -1064 7580
rect -1008 7524 -984 7580
rect -928 7524 -904 7580
rect -848 7524 -824 7580
rect -768 7524 -756 7580
rect -1076 7500 -756 7524
rect -1076 7444 -1064 7500
rect -1008 7444 -984 7500
rect -928 7444 -904 7500
rect -848 7444 -824 7500
rect -768 7444 -756 7500
rect -1076 6381 -756 7444
rect -1076 6325 -1064 6381
rect -1008 6325 -984 6381
rect -928 6325 -904 6381
rect -848 6325 -824 6381
rect -768 6325 -756 6381
rect -1076 6301 -756 6325
rect -1076 6245 -1064 6301
rect -1008 6245 -984 6301
rect -928 6245 -904 6301
rect -848 6245 -824 6301
rect -768 6245 -756 6301
rect -1076 6221 -756 6245
rect -1076 6165 -1064 6221
rect -1008 6165 -984 6221
rect -928 6165 -904 6221
rect -848 6165 -824 6221
rect -768 6165 -756 6221
rect -1076 6141 -756 6165
rect -1076 6085 -1064 6141
rect -1008 6085 -984 6141
rect -928 6085 -904 6141
rect -848 6085 -824 6141
rect -768 6085 -756 6141
rect -1076 5022 -756 6085
rect -1076 4966 -1064 5022
rect -1008 4966 -984 5022
rect -928 4966 -904 5022
rect -848 4966 -824 5022
rect -768 4966 -756 5022
rect -1076 4942 -756 4966
rect -1076 4886 -1064 4942
rect -1008 4886 -984 4942
rect -928 4886 -904 4942
rect -848 4886 -824 4942
rect -768 4886 -756 4942
rect -1076 4862 -756 4886
rect -1076 4806 -1064 4862
rect -1008 4806 -984 4862
rect -928 4806 -904 4862
rect -848 4806 -824 4862
rect -768 4806 -756 4862
rect -1076 4782 -756 4806
rect -1076 4726 -1064 4782
rect -1008 4726 -984 4782
rect -928 4726 -904 4782
rect -848 4726 -824 4782
rect -768 4726 -756 4782
rect -1076 3663 -756 4726
rect -1076 3607 -1064 3663
rect -1008 3607 -984 3663
rect -928 3607 -904 3663
rect -848 3607 -824 3663
rect -768 3607 -756 3663
rect -1076 3583 -756 3607
rect -1076 3527 -1064 3583
rect -1008 3527 -984 3583
rect -928 3527 -904 3583
rect -848 3527 -824 3583
rect -768 3527 -756 3583
rect -1076 3503 -756 3527
rect -1076 3447 -1064 3503
rect -1008 3447 -984 3503
rect -928 3447 -904 3503
rect -848 3447 -824 3503
rect -768 3447 -756 3503
rect -1076 3423 -756 3447
rect -1076 3367 -1064 3423
rect -1008 3367 -984 3423
rect -928 3367 -904 3423
rect -848 3367 -824 3423
rect -768 3367 -756 3423
rect -1076 304 -756 3367
rect -416 9124 -96 9136
rect -416 9068 -404 9124
rect -348 9068 -324 9124
rect -268 9068 -244 9124
rect -188 9068 -164 9124
rect -108 9068 -96 9124
rect -416 9044 -96 9068
rect -416 8988 -404 9044
rect -348 8988 -324 9044
rect -268 8988 -244 9044
rect -188 8988 -164 9044
rect -108 8988 -96 9044
rect -416 8964 -96 8988
rect -416 8908 -404 8964
rect -348 8908 -324 8964
rect -268 8908 -244 8964
rect -188 8908 -164 8964
rect -108 8908 -96 8964
rect -416 8884 -96 8908
rect -416 8828 -404 8884
rect -348 8828 -324 8884
rect -268 8828 -244 8884
rect -188 8828 -164 8884
rect -108 8828 -96 8884
rect -416 7080 -96 8828
rect -416 7024 -404 7080
rect -348 7024 -324 7080
rect -268 7024 -244 7080
rect -188 7024 -164 7080
rect -108 7024 -96 7080
rect -416 7000 -96 7024
rect -416 6944 -404 7000
rect -348 6944 -324 7000
rect -268 6944 -244 7000
rect -188 6944 -164 7000
rect -108 6944 -96 7000
rect -416 6920 -96 6944
rect -416 6864 -404 6920
rect -348 6864 -324 6920
rect -268 6864 -244 6920
rect -188 6864 -164 6920
rect -108 6864 -96 6920
rect -416 6840 -96 6864
rect -416 6784 -404 6840
rect -348 6784 -324 6840
rect -268 6784 -244 6840
rect -188 6784 -164 6840
rect -108 6784 -96 6840
rect -416 5721 -96 6784
rect -416 5665 -404 5721
rect -348 5665 -324 5721
rect -268 5665 -244 5721
rect -188 5665 -164 5721
rect -108 5665 -96 5721
rect -416 5641 -96 5665
rect -416 5585 -404 5641
rect -348 5585 -324 5641
rect -268 5585 -244 5641
rect -188 5585 -164 5641
rect -108 5585 -96 5641
rect -416 5561 -96 5585
rect -416 5505 -404 5561
rect -348 5505 -324 5561
rect -268 5505 -244 5561
rect -188 5505 -164 5561
rect -108 5505 -96 5561
rect -416 5481 -96 5505
rect -416 5425 -404 5481
rect -348 5425 -324 5481
rect -268 5425 -244 5481
rect -188 5425 -164 5481
rect -108 5425 -96 5481
rect -416 4362 -96 5425
rect -416 4306 -404 4362
rect -348 4306 -324 4362
rect -268 4306 -244 4362
rect -188 4306 -164 4362
rect -108 4306 -96 4362
rect -416 4282 -96 4306
rect -416 4226 -404 4282
rect -348 4226 -324 4282
rect -268 4226 -244 4282
rect -188 4226 -164 4282
rect -108 4226 -96 4282
rect -416 4202 -96 4226
rect -416 4146 -404 4202
rect -348 4146 -324 4202
rect -268 4146 -244 4202
rect -188 4146 -164 4202
rect -108 4146 -96 4202
rect -416 4122 -96 4146
rect -416 4066 -404 4122
rect -348 4066 -324 4122
rect -268 4066 -244 4122
rect -188 4066 -164 4122
rect -108 4066 -96 4122
rect -416 3003 -96 4066
rect -416 2947 -404 3003
rect -348 2947 -324 3003
rect -268 2947 -244 3003
rect -188 2947 -164 3003
rect -108 2947 -96 3003
rect -416 2923 -96 2947
rect -416 2867 -404 2923
rect -348 2867 -324 2923
rect -268 2867 -244 2923
rect -188 2867 -164 2923
rect -108 2867 -96 2923
rect -416 2843 -96 2867
rect -416 2787 -404 2843
rect -348 2787 -324 2843
rect -268 2787 -244 2843
rect -188 2787 -164 2843
rect -108 2787 -96 2843
rect -416 2763 -96 2787
rect -416 2707 -404 2763
rect -348 2707 -324 2763
rect -268 2707 -244 2763
rect -188 2707 -164 2763
rect -108 2707 -96 2763
rect -416 964 -96 2707
rect 1872 2650 1900 9182
rect 16592 2650 16620 9182
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 31772 2446 31800 9182
rect 46940 8968 46992 8974
rect 46940 8910 46992 8916
rect 46952 2650 46980 8910
rect 62040 6866 62068 9182
rect 76944 6866 76972 9182
rect 86159 9124 86479 9796
rect 86159 9068 86171 9124
rect 86227 9068 86251 9124
rect 86307 9068 86331 9124
rect 86387 9068 86411 9124
rect 86467 9068 86479 9124
rect 86159 9044 86479 9068
rect 86159 8988 86171 9044
rect 86227 8988 86251 9044
rect 86307 8988 86331 9044
rect 86387 8988 86411 9044
rect 86467 8988 86479 9044
rect 86159 8964 86479 8988
rect 86159 8908 86171 8964
rect 86227 8908 86251 8964
rect 86307 8908 86331 8964
rect 86387 8908 86411 8964
rect 86467 8908 86479 8964
rect 86159 8884 86479 8908
rect 86159 8828 86171 8884
rect 86227 8828 86251 8884
rect 86307 8828 86331 8884
rect 86387 8828 86411 8884
rect 86467 8828 86479 8884
rect 86159 7098 86479 8828
rect 86159 7046 86165 7098
rect 86217 7080 86229 7098
rect 86281 7080 86293 7098
rect 86345 7080 86357 7098
rect 86409 7080 86421 7098
rect 86227 7046 86229 7080
rect 86409 7046 86411 7080
rect 86473 7046 86479 7098
rect 86159 7024 86171 7046
rect 86227 7024 86251 7046
rect 86307 7024 86331 7046
rect 86387 7024 86411 7046
rect 86467 7024 86479 7046
rect 86159 7000 86479 7024
rect 86159 6944 86171 7000
rect 86227 6944 86251 7000
rect 86307 6944 86331 7000
rect 86387 6944 86411 7000
rect 86467 6944 86479 7000
rect 86159 6920 86479 6944
rect 62028 6860 62080 6866
rect 62028 6802 62080 6808
rect 63684 6860 63736 6866
rect 63684 6802 63736 6808
rect 76932 6860 76984 6866
rect 76932 6802 76984 6808
rect 78864 6860 78916 6866
rect 78864 6802 78916 6808
rect 86159 6864 86171 6920
rect 86227 6864 86251 6920
rect 86307 6864 86331 6920
rect 86387 6864 86411 6920
rect 86467 6864 86479 6920
rect 86159 6840 86479 6864
rect 63696 2650 63724 6802
rect 78876 3194 78904 6802
rect 86159 6784 86171 6840
rect 86227 6784 86251 6840
rect 86307 6784 86331 6840
rect 86387 6784 86411 6840
rect 86467 6784 86479 6840
rect 86159 6010 86479 6784
rect 86159 5958 86165 6010
rect 86217 5958 86229 6010
rect 86281 5958 86293 6010
rect 86345 5958 86357 6010
rect 86409 5958 86421 6010
rect 86473 5958 86479 6010
rect 86159 5721 86479 5958
rect 86159 5665 86171 5721
rect 86227 5665 86251 5721
rect 86307 5665 86331 5721
rect 86387 5665 86411 5721
rect 86467 5665 86479 5721
rect 86159 5641 86479 5665
rect 86159 5585 86171 5641
rect 86227 5585 86251 5641
rect 86307 5585 86331 5641
rect 86387 5585 86411 5641
rect 86467 5585 86479 5641
rect 86159 5561 86479 5585
rect 86159 5505 86171 5561
rect 86227 5505 86251 5561
rect 86307 5505 86331 5561
rect 86387 5505 86411 5561
rect 86467 5505 86479 5561
rect 86159 5481 86479 5505
rect 86159 5425 86171 5481
rect 86227 5425 86251 5481
rect 86307 5425 86331 5481
rect 86387 5425 86411 5481
rect 86467 5425 86479 5481
rect 86159 4922 86479 5425
rect 86159 4870 86165 4922
rect 86217 4870 86229 4922
rect 86281 4870 86293 4922
rect 86345 4870 86357 4922
rect 86409 4870 86421 4922
rect 86473 4870 86479 4922
rect 86159 4362 86479 4870
rect 86159 4306 86171 4362
rect 86227 4306 86251 4362
rect 86307 4306 86331 4362
rect 86387 4306 86411 4362
rect 86467 4306 86479 4362
rect 86159 4282 86479 4306
rect 86159 4226 86171 4282
rect 86227 4226 86251 4282
rect 86307 4226 86331 4282
rect 86387 4226 86411 4282
rect 86467 4226 86479 4282
rect 86159 4202 86479 4226
rect 86159 4146 86171 4202
rect 86227 4146 86251 4202
rect 86307 4146 86331 4202
rect 86387 4146 86411 4202
rect 86467 4146 86479 4202
rect 86159 4122 86479 4146
rect 86159 4066 86171 4122
rect 86227 4066 86251 4122
rect 86307 4066 86331 4122
rect 86387 4066 86411 4122
rect 86467 4066 86479 4122
rect 86159 3834 86479 4066
rect 86159 3782 86165 3834
rect 86217 3782 86229 3834
rect 86281 3782 86293 3834
rect 86345 3782 86357 3834
rect 86409 3782 86421 3834
rect 86473 3782 86479 3834
rect 78864 3188 78916 3194
rect 78864 3130 78916 3136
rect 46940 2644 46992 2650
rect 46940 2586 46992 2592
rect 63684 2644 63736 2650
rect 63684 2586 63736 2592
rect 78876 2446 78904 3130
rect 86159 3003 86479 3782
rect 86159 2947 86171 3003
rect 86227 2947 86251 3003
rect 86307 2947 86331 3003
rect 86387 2947 86411 3003
rect 86467 2947 86479 3003
rect 86159 2923 86479 2947
rect 86159 2867 86171 2923
rect 86227 2867 86251 2923
rect 86307 2867 86331 2923
rect 86387 2867 86411 2923
rect 86467 2867 86479 2923
rect 86159 2843 86479 2867
rect 86159 2787 86171 2843
rect 86227 2787 86251 2843
rect 86307 2787 86331 2843
rect 86387 2787 86411 2843
rect 86467 2787 86479 2843
rect 86159 2763 86479 2787
rect 86159 2746 86171 2763
rect 86227 2746 86251 2763
rect 86307 2746 86331 2763
rect 86387 2746 86411 2763
rect 86467 2746 86479 2763
rect 86159 2694 86165 2746
rect 86227 2707 86229 2746
rect 86409 2707 86411 2746
rect 86217 2694 86229 2707
rect 86281 2694 86293 2707
rect 86345 2694 86357 2707
rect 86409 2694 86421 2707
rect 86473 2694 86479 2746
rect 31760 2440 31812 2446
rect 31760 2382 31812 2388
rect 78864 2440 78916 2446
rect 78864 2382 78916 2388
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 79140 2304 79192 2310
rect 79140 2246 79192 2252
rect 2608 2106 2636 2246
rect 2596 2100 2648 2106
rect 2596 2042 2648 2048
rect 18064 1970 18092 2246
rect 79152 2038 79180 2246
rect 79140 2032 79192 2038
rect 79140 1974 79192 1980
rect 18052 1964 18104 1970
rect 18052 1906 18104 1912
rect -416 908 -404 964
rect -348 908 -324 964
rect -268 908 -244 964
rect -188 908 -164 964
rect -108 908 -96 964
rect -416 884 -96 908
rect -416 828 -404 884
rect -348 828 -324 884
rect -268 828 -244 884
rect -188 828 -164 884
rect -108 828 -96 884
rect -416 804 -96 828
rect -416 748 -404 804
rect -348 748 -324 804
rect -268 748 -244 804
rect -188 748 -164 804
rect -108 748 -96 804
rect -416 724 -96 748
rect -416 668 -404 724
rect -348 668 -324 724
rect -268 668 -244 724
rect -188 668 -164 724
rect -108 668 -96 724
rect -416 656 -96 668
rect 86159 964 86479 2694
rect 86159 908 86171 964
rect 86227 908 86251 964
rect 86307 908 86331 964
rect 86387 908 86411 964
rect 86467 908 86479 964
rect 86159 884 86479 908
rect 86159 828 86171 884
rect 86227 828 86251 884
rect 86307 828 86331 884
rect 86387 828 86411 884
rect 86467 828 86479 884
rect 86159 804 86479 828
rect 86159 748 86171 804
rect 86227 748 86251 804
rect 86307 748 86331 804
rect 86387 748 86411 804
rect 86467 748 86479 804
rect 86159 724 86479 748
rect 86159 668 86171 724
rect 86227 668 86251 724
rect 86307 668 86331 724
rect 86387 668 86411 724
rect 86467 668 86479 724
rect -1076 248 -1064 304
rect -1008 248 -984 304
rect -928 248 -904 304
rect -848 248 -824 304
rect -768 248 -756 304
rect -1076 224 -756 248
rect -1076 168 -1064 224
rect -1008 168 -984 224
rect -928 168 -904 224
rect -848 168 -824 224
rect -768 168 -756 224
rect -1076 144 -756 168
rect -1076 88 -1064 144
rect -1008 88 -984 144
rect -928 88 -904 144
rect -848 88 -824 144
rect -768 88 -756 144
rect -1076 64 -756 88
rect -1076 8 -1064 64
rect -1008 8 -984 64
rect -928 8 -904 64
rect -848 8 -824 64
rect -768 8 -756 64
rect -1076 -4 -756 8
rect 86159 -4 86479 668
rect 86819 9784 87139 9796
rect 86819 9728 86831 9784
rect 86887 9728 86911 9784
rect 86967 9728 86991 9784
rect 87047 9728 87071 9784
rect 87127 9728 87139 9784
rect 86819 9704 87139 9728
rect 86819 9648 86831 9704
rect 86887 9648 86911 9704
rect 86967 9648 86991 9704
rect 87047 9648 87071 9704
rect 87127 9648 87139 9704
rect 86819 9624 87139 9648
rect 86819 9568 86831 9624
rect 86887 9568 86911 9624
rect 86967 9568 86991 9624
rect 87047 9568 87071 9624
rect 87127 9568 87139 9624
rect 86819 9544 87139 9568
rect 86819 9488 86831 9544
rect 86887 9488 86911 9544
rect 86967 9488 86991 9544
rect 87047 9488 87071 9544
rect 87127 9488 87139 9544
rect 86819 7740 87139 9488
rect 107568 9240 107620 9246
rect 107568 9182 107620 9188
rect 122748 9240 122800 9246
rect 122748 9182 122800 9188
rect 169668 9240 169720 9246
rect 169668 9182 169720 9188
rect 184848 9240 184900 9246
rect 184848 9182 184900 9188
rect 215208 9240 215260 9246
rect 215208 9182 215260 9188
rect 230388 9240 230440 9246
rect 230388 9182 230440 9188
rect 92388 8968 92440 8974
rect 92388 8910 92440 8916
rect 86819 7684 86831 7740
rect 86887 7684 86911 7740
rect 86967 7684 86991 7740
rect 87047 7684 87071 7740
rect 87127 7684 87139 7740
rect 86819 7660 87139 7684
rect 86819 7642 86831 7660
rect 86887 7642 86911 7660
rect 86967 7642 86991 7660
rect 87047 7642 87071 7660
rect 87127 7642 87139 7660
rect 86819 7590 86825 7642
rect 86887 7604 86889 7642
rect 87069 7604 87071 7642
rect 86877 7590 86889 7604
rect 86941 7590 86953 7604
rect 87005 7590 87017 7604
rect 87069 7590 87081 7604
rect 87133 7590 87139 7642
rect 86819 7580 87139 7590
rect 86819 7524 86831 7580
rect 86887 7524 86911 7580
rect 86967 7524 86991 7580
rect 87047 7524 87071 7580
rect 87127 7524 87139 7580
rect 86819 7500 87139 7524
rect 86819 7444 86831 7500
rect 86887 7444 86911 7500
rect 86967 7444 86991 7500
rect 87047 7444 87071 7500
rect 87127 7444 87139 7500
rect 86819 6554 87139 7444
rect 92400 6866 92428 8910
rect 107580 6866 107608 9182
rect 122760 6866 122788 9182
rect 137928 8968 137980 8974
rect 137928 8910 137980 8916
rect 153108 8968 153160 8974
rect 153108 8910 153160 8916
rect 137940 6866 137968 8910
rect 153120 6866 153148 8910
rect 169680 6866 169708 9182
rect 184860 6866 184888 9182
rect 200028 8968 200080 8974
rect 200028 8910 200080 8916
rect 200040 6866 200068 8910
rect 215220 6866 215248 9182
rect 230400 6866 230428 9182
rect 256589 9124 256909 9796
rect 256589 9068 256601 9124
rect 256657 9068 256681 9124
rect 256737 9068 256761 9124
rect 256817 9068 256841 9124
rect 256897 9068 256909 9124
rect 256589 9044 256909 9068
rect 256589 8988 256601 9044
rect 256657 8988 256681 9044
rect 256737 8988 256761 9044
rect 256817 8988 256841 9044
rect 256897 8988 256909 9044
rect 245568 8968 245620 8974
rect 245568 8910 245620 8916
rect 256589 8964 256909 8988
rect 245580 6866 245608 8910
rect 256589 8908 256601 8964
rect 256657 8908 256681 8964
rect 256737 8908 256761 8964
rect 256817 8908 256841 8964
rect 256897 8908 256909 8964
rect 256589 8884 256909 8908
rect 256589 8828 256601 8884
rect 256657 8828 256681 8884
rect 256737 8828 256761 8884
rect 256817 8828 256841 8884
rect 256897 8828 256909 8884
rect 256589 7098 256909 8828
rect 256589 7046 256595 7098
rect 256647 7080 256659 7098
rect 256711 7080 256723 7098
rect 256775 7080 256787 7098
rect 256839 7080 256851 7098
rect 256657 7046 256659 7080
rect 256839 7046 256841 7080
rect 256903 7046 256909 7098
rect 256589 7024 256601 7046
rect 256657 7024 256681 7046
rect 256737 7024 256761 7046
rect 256817 7024 256841 7046
rect 256897 7024 256909 7046
rect 256589 7000 256909 7024
rect 256589 6944 256601 7000
rect 256657 6944 256681 7000
rect 256737 6944 256761 7000
rect 256817 6944 256841 7000
rect 256897 6944 256909 7000
rect 256589 6920 256909 6944
rect 92388 6860 92440 6866
rect 92388 6802 92440 6808
rect 94596 6860 94648 6866
rect 94596 6802 94648 6808
rect 107568 6860 107620 6866
rect 107568 6802 107620 6808
rect 110052 6860 110104 6866
rect 110052 6802 110104 6808
rect 122748 6860 122800 6866
rect 122748 6802 122800 6808
rect 125508 6860 125560 6866
rect 125508 6802 125560 6808
rect 137928 6860 137980 6866
rect 137928 6802 137980 6808
rect 140688 6860 140740 6866
rect 140688 6802 140740 6808
rect 153108 6860 153160 6866
rect 153108 6802 153160 6808
rect 155868 6860 155920 6866
rect 155868 6802 155920 6808
rect 169668 6860 169720 6866
rect 169668 6802 169720 6808
rect 171600 6860 171652 6866
rect 171600 6802 171652 6808
rect 184848 6860 184900 6866
rect 184848 6802 184900 6808
rect 187332 6860 187384 6866
rect 187332 6802 187384 6808
rect 200028 6860 200080 6866
rect 200028 6802 200080 6808
rect 202788 6860 202840 6866
rect 202788 6802 202840 6808
rect 215208 6860 215260 6866
rect 215208 6802 215260 6808
rect 218060 6860 218112 6866
rect 218060 6802 218112 6808
rect 230388 6860 230440 6866
rect 230388 6802 230440 6808
rect 233056 6860 233108 6866
rect 233056 6802 233108 6808
rect 245568 6860 245620 6866
rect 245568 6802 245620 6808
rect 249156 6860 249208 6866
rect 249156 6802 249208 6808
rect 256589 6864 256601 6920
rect 256657 6864 256681 6920
rect 256737 6864 256761 6920
rect 256817 6864 256841 6920
rect 256897 6864 256909 6920
rect 256589 6840 256909 6864
rect 86819 6502 86825 6554
rect 86877 6502 86889 6554
rect 86941 6502 86953 6554
rect 87005 6502 87017 6554
rect 87069 6502 87081 6554
rect 87133 6502 87139 6554
rect 86819 6381 87139 6502
rect 86819 6325 86831 6381
rect 86887 6325 86911 6381
rect 86967 6325 86991 6381
rect 87047 6325 87071 6381
rect 87127 6325 87139 6381
rect 86819 6301 87139 6325
rect 86819 6245 86831 6301
rect 86887 6245 86911 6301
rect 86967 6245 86991 6301
rect 87047 6245 87071 6301
rect 87127 6245 87139 6301
rect 86819 6221 87139 6245
rect 86819 6165 86831 6221
rect 86887 6165 86911 6221
rect 86967 6165 86991 6221
rect 87047 6165 87071 6221
rect 87127 6165 87139 6221
rect 86819 6141 87139 6165
rect 86819 6085 86831 6141
rect 86887 6085 86911 6141
rect 86967 6085 86991 6141
rect 87047 6085 87071 6141
rect 87127 6085 87139 6141
rect 86819 5466 87139 6085
rect 86819 5414 86825 5466
rect 86877 5414 86889 5466
rect 86941 5414 86953 5466
rect 87005 5414 87017 5466
rect 87069 5414 87081 5466
rect 87133 5414 87139 5466
rect 86819 5022 87139 5414
rect 86819 4966 86831 5022
rect 86887 4966 86911 5022
rect 86967 4966 86991 5022
rect 87047 4966 87071 5022
rect 87127 4966 87139 5022
rect 86819 4942 87139 4966
rect 86819 4886 86831 4942
rect 86887 4886 86911 4942
rect 86967 4886 86991 4942
rect 87047 4886 87071 4942
rect 87127 4886 87139 4942
rect 86819 4862 87139 4886
rect 86819 4806 86831 4862
rect 86887 4806 86911 4862
rect 86967 4806 86991 4862
rect 87047 4806 87071 4862
rect 87127 4806 87139 4862
rect 86819 4782 87139 4806
rect 86819 4726 86831 4782
rect 86887 4726 86911 4782
rect 86967 4726 86991 4782
rect 87047 4726 87071 4782
rect 87127 4726 87139 4782
rect 86819 4378 87139 4726
rect 86819 4326 86825 4378
rect 86877 4326 86889 4378
rect 86941 4326 86953 4378
rect 87005 4326 87017 4378
rect 87069 4326 87081 4378
rect 87133 4326 87139 4378
rect 86819 3663 87139 4326
rect 86819 3607 86831 3663
rect 86887 3607 86911 3663
rect 86967 3607 86991 3663
rect 87047 3607 87071 3663
rect 87127 3607 87139 3663
rect 86819 3583 87139 3607
rect 86819 3527 86831 3583
rect 86887 3527 86911 3583
rect 86967 3527 86991 3583
rect 87047 3527 87071 3583
rect 87127 3527 87139 3583
rect 86819 3503 87139 3527
rect 86819 3447 86831 3503
rect 86887 3447 86911 3503
rect 86967 3447 86991 3503
rect 87047 3447 87071 3503
rect 87127 3447 87139 3503
rect 86819 3423 87139 3447
rect 86819 3367 86831 3423
rect 86887 3367 86911 3423
rect 86967 3367 86991 3423
rect 87047 3367 87071 3423
rect 87127 3367 87139 3423
rect 86819 3290 87139 3367
rect 86819 3238 86825 3290
rect 86877 3238 86889 3290
rect 86941 3238 86953 3290
rect 87005 3238 87017 3290
rect 87069 3238 87081 3290
rect 87133 3238 87139 3290
rect 86819 2202 87139 3238
rect 94608 2650 94636 6802
rect 94596 2644 94648 2650
rect 94596 2586 94648 2592
rect 97356 2644 97408 2650
rect 97356 2586 97408 2592
rect 97368 2446 97396 2586
rect 95332 2440 95384 2446
rect 95332 2382 95384 2388
rect 97356 2440 97408 2446
rect 97356 2382 97408 2388
rect 95344 2310 95372 2382
rect 96804 2372 96856 2378
rect 96804 2314 96856 2320
rect 95332 2304 95384 2310
rect 95332 2246 95384 2252
rect 86819 2150 86825 2202
rect 86877 2150 86889 2202
rect 86941 2150 86953 2202
rect 87005 2150 87017 2202
rect 87069 2150 87081 2202
rect 87133 2150 87139 2202
rect 86819 304 87139 2150
rect 95344 1834 95372 2246
rect 96816 2106 96844 2314
rect 110064 2310 110092 6802
rect 125520 2446 125548 6802
rect 136548 2848 136600 2854
rect 136548 2790 136600 2796
rect 136560 2446 136588 2790
rect 140700 2582 140728 6802
rect 155880 2582 155908 6802
rect 171612 3194 171640 6802
rect 171600 3188 171652 3194
rect 171600 3130 171652 3136
rect 140688 2576 140740 2582
rect 140688 2518 140740 2524
rect 155868 2576 155920 2582
rect 155868 2518 155920 2524
rect 138388 2508 138440 2514
rect 138388 2450 138440 2456
rect 110696 2440 110748 2446
rect 110696 2382 110748 2388
rect 113456 2440 113508 2446
rect 113456 2382 113508 2388
rect 125508 2440 125560 2446
rect 125508 2382 125560 2388
rect 136548 2440 136600 2446
rect 136548 2382 136600 2388
rect 138112 2440 138164 2446
rect 138400 2394 138428 2450
rect 171612 2446 171640 3130
rect 187344 2650 187372 6802
rect 187700 2848 187752 2854
rect 187700 2790 187752 2796
rect 187332 2644 187384 2650
rect 187332 2586 187384 2592
rect 138112 2382 138164 2388
rect 110708 2310 110736 2382
rect 112260 2372 112312 2378
rect 112260 2314 112312 2320
rect 110052 2304 110104 2310
rect 110052 2246 110104 2252
rect 110696 2304 110748 2310
rect 110696 2246 110748 2252
rect 110708 2106 110736 2246
rect 96804 2100 96856 2106
rect 96804 2042 96856 2048
rect 110696 2100 110748 2106
rect 110696 2042 110748 2048
rect 112272 1970 112300 2314
rect 113468 2310 113496 2382
rect 135996 2372 136048 2378
rect 135996 2314 136048 2320
rect 113456 2304 113508 2310
rect 113456 2246 113508 2252
rect 125692 2304 125744 2310
rect 125692 2246 125744 2252
rect 112260 1964 112312 1970
rect 112260 1906 112312 1912
rect 95332 1828 95384 1834
rect 95332 1770 95384 1776
rect 113468 1766 113496 2246
rect 125704 1970 125732 2246
rect 125692 1964 125744 1970
rect 125692 1906 125744 1912
rect 113456 1760 113508 1766
rect 113456 1702 113508 1708
rect 136008 950 136036 2314
rect 136560 2038 136588 2382
rect 136824 2372 136876 2378
rect 136824 2314 136876 2320
rect 136548 2032 136600 2038
rect 136548 1974 136600 1980
rect 135996 944 136048 950
rect 135996 886 136048 892
rect 86819 248 86831 304
rect 86887 248 86911 304
rect 86967 248 86991 304
rect 87047 248 87071 304
rect 87127 248 87139 304
rect 136836 270 136864 2314
rect 138124 1970 138152 2382
rect 138216 2366 138428 2394
rect 141700 2440 141752 2446
rect 141700 2382 141752 2388
rect 157156 2440 157208 2446
rect 157156 2382 157208 2388
rect 171600 2440 171652 2446
rect 171600 2382 171652 2388
rect 138216 2310 138244 2366
rect 141712 2310 141740 2382
rect 157168 2310 157196 2382
rect 187712 2310 187740 2790
rect 202800 2650 202828 6802
rect 218072 3194 218100 6802
rect 218060 3188 218112 3194
rect 218060 3130 218112 3136
rect 202972 2848 203024 2854
rect 202972 2790 203024 2796
rect 202788 2644 202840 2650
rect 202788 2586 202840 2592
rect 202984 2446 203012 2790
rect 218072 2446 218100 3130
rect 233068 2650 233096 6802
rect 248420 3392 248472 3398
rect 248420 3334 248472 3340
rect 242164 3188 242216 3194
rect 242164 3130 242216 3136
rect 233056 2644 233108 2650
rect 233056 2586 233108 2592
rect 218244 2576 218296 2582
rect 238024 2576 238076 2582
rect 218244 2518 218296 2524
rect 236826 2544 236882 2553
rect 189540 2440 189592 2446
rect 189540 2382 189592 2388
rect 191380 2440 191432 2446
rect 191380 2382 191432 2388
rect 202972 2440 203024 2446
rect 202972 2382 203024 2388
rect 218060 2440 218112 2446
rect 218060 2382 218112 2388
rect 188620 2372 188672 2378
rect 188620 2314 188672 2320
rect 138204 2304 138256 2310
rect 138204 2246 138256 2252
rect 138296 2304 138348 2310
rect 138296 2246 138348 2252
rect 141700 2304 141752 2310
rect 141700 2246 141752 2252
rect 144368 2304 144420 2310
rect 144368 2246 144420 2252
rect 157156 2304 157208 2310
rect 157156 2246 157208 2252
rect 159824 2304 159876 2310
rect 159824 2246 159876 2252
rect 171876 2304 171928 2310
rect 171876 2246 171928 2252
rect 187700 2304 187752 2310
rect 187700 2246 187752 2252
rect 138112 1964 138164 1970
rect 138112 1906 138164 1912
rect 138308 882 138336 2246
rect 141712 1018 141740 2246
rect 144380 1086 144408 2246
rect 157168 1154 157196 2246
rect 159836 1222 159864 2246
rect 171888 1290 171916 2246
rect 188632 1834 188660 2314
rect 188620 1828 188672 1834
rect 188620 1770 188672 1776
rect 189552 1358 189580 2382
rect 191392 2310 191420 2382
rect 191380 2304 191432 2310
rect 191380 2246 191432 2252
rect 189540 1352 189592 1358
rect 189540 1294 189592 1300
rect 171876 1284 171928 1290
rect 171876 1226 171928 1232
rect 159824 1216 159876 1222
rect 159824 1158 159876 1164
rect 157156 1148 157208 1154
rect 157156 1090 157208 1096
rect 144368 1080 144420 1086
rect 144368 1022 144420 1028
rect 141700 1012 141752 1018
rect 141700 954 141752 960
rect 138296 876 138348 882
rect 138296 818 138348 824
rect 86819 224 87139 248
rect 86819 168 86831 224
rect 86887 168 86911 224
rect 86967 168 86991 224
rect 87047 168 87071 224
rect 87127 168 87139 224
rect 136824 264 136876 270
rect 136824 206 136876 212
rect 86819 144 87139 168
rect 86819 88 86831 144
rect 86887 88 86911 144
rect 86967 88 86991 144
rect 87047 88 87071 144
rect 87127 88 87139 144
rect 86819 64 87139 88
rect 191392 66 191420 2246
rect 202984 202 203012 2382
rect 203892 2372 203944 2378
rect 203892 2314 203944 2320
rect 205916 2372 205968 2378
rect 205916 2314 205968 2320
rect 203904 2106 203932 2314
rect 203892 2100 203944 2106
rect 203892 2042 203944 2048
rect 205928 1766 205956 2314
rect 218256 2106 218284 2518
rect 228180 2508 228232 2514
rect 238024 2518 238076 2524
rect 236826 2479 236882 2488
rect 228180 2450 228232 2456
rect 218244 2100 218296 2106
rect 218244 2042 218296 2048
rect 205916 1760 205968 1766
rect 205916 1702 205968 1708
rect 227260 1352 227312 1358
rect 227260 1294 227312 1300
rect 227812 1352 227864 1358
rect 227812 1294 227864 1300
rect 224224 1080 224276 1086
rect 224224 1022 224276 1028
rect 224236 898 224264 1022
rect 224316 1012 224368 1018
rect 224316 954 224368 960
rect 224144 870 224264 898
rect 224144 746 224172 870
rect 224132 740 224184 746
rect 224132 682 224184 688
rect 224328 354 224356 954
rect 227272 882 227300 1294
rect 227628 1216 227680 1222
rect 227442 1184 227498 1193
rect 227628 1158 227680 1164
rect 227442 1119 227444 1128
rect 227496 1119 227498 1128
rect 227444 1090 227496 1096
rect 227260 876 227312 882
rect 227260 818 227312 824
rect 227640 814 227668 1158
rect 227720 1148 227772 1154
rect 227720 1090 227772 1096
rect 227628 808 227680 814
rect 227628 750 227680 756
rect 227732 678 227760 1090
rect 227720 672 227772 678
rect 227720 614 227772 620
rect 224144 326 224356 354
rect 224144 270 224172 326
rect 224132 264 224184 270
rect 227824 218 227852 1294
rect 228192 814 228220 2450
rect 232688 2372 232740 2378
rect 232688 2314 232740 2320
rect 230664 2304 230716 2310
rect 230664 2246 230716 2252
rect 229376 1284 229428 1290
rect 229376 1226 229428 1232
rect 229468 1284 229520 1290
rect 229468 1226 229520 1232
rect 228640 1080 228692 1086
rect 228640 1022 228692 1028
rect 228732 1080 228784 1086
rect 228732 1022 228784 1028
rect 228652 814 228680 1022
rect 228744 882 228772 1022
rect 228732 876 228784 882
rect 228732 818 228784 824
rect 229388 814 229416 1226
rect 229480 1193 229508 1226
rect 229466 1184 229522 1193
rect 229466 1119 229522 1128
rect 230676 814 230704 2246
rect 231768 2100 231820 2106
rect 231768 2042 231820 2048
rect 231780 1426 231808 2042
rect 232228 1488 232280 1494
rect 232228 1430 232280 1436
rect 231768 1420 231820 1426
rect 231768 1362 231820 1368
rect 231952 1284 232004 1290
rect 231952 1226 232004 1232
rect 228180 808 228232 814
rect 228180 750 228232 756
rect 228640 808 228692 814
rect 228640 750 228692 756
rect 229376 808 229428 814
rect 229376 750 229428 756
rect 230664 808 230716 814
rect 230664 750 230716 756
rect 231964 678 231992 1226
rect 232240 1154 232268 1430
rect 232228 1148 232280 1154
rect 232228 1090 232280 1096
rect 232700 814 232728 2314
rect 234344 2304 234396 2310
rect 234344 2246 234396 2252
rect 234356 814 234384 2246
rect 235540 2032 235592 2038
rect 235540 1974 235592 1980
rect 235264 1488 235316 1494
rect 235264 1430 235316 1436
rect 235276 814 235304 1430
rect 235552 814 235580 1974
rect 236000 1964 236052 1970
rect 236000 1906 236052 1912
rect 236012 814 236040 1906
rect 236840 814 236868 2479
rect 237196 1352 237248 1358
rect 237196 1294 237248 1300
rect 237208 814 237236 1294
rect 238036 814 238064 2518
rect 240140 2508 240192 2514
rect 240140 2450 240192 2456
rect 239588 2304 239640 2310
rect 239588 2246 239640 2252
rect 238484 1896 238536 1902
rect 238484 1838 238536 1844
rect 238496 814 238524 1838
rect 239600 814 239628 2246
rect 239954 1456 240010 1465
rect 239954 1391 240010 1400
rect 239968 1222 239996 1391
rect 239956 1216 240008 1222
rect 239956 1158 240008 1164
rect 240048 1216 240100 1222
rect 240048 1158 240100 1164
rect 240060 814 240088 1158
rect 240152 950 240180 2450
rect 242070 1728 242126 1737
rect 241520 1692 241572 1698
rect 242070 1663 242126 1672
rect 241520 1634 241572 1640
rect 240140 944 240192 950
rect 240140 886 240192 892
rect 241244 876 241296 882
rect 241532 864 241560 1634
rect 241794 1592 241850 1601
rect 241794 1527 241850 1536
rect 241296 836 241560 864
rect 241244 818 241296 824
rect 241808 814 241836 1527
rect 241888 1488 241940 1494
rect 241888 1430 241940 1436
rect 241900 1018 241928 1430
rect 242084 1154 242112 1663
rect 242072 1148 242124 1154
rect 242072 1090 242124 1096
rect 241888 1012 241940 1018
rect 241888 954 241940 960
rect 242176 814 242204 3130
rect 247040 3120 247092 3126
rect 247040 3062 247092 3068
rect 244280 2644 244332 2650
rect 244280 2586 244332 2592
rect 243268 2100 243320 2106
rect 243268 2042 243320 2048
rect 242532 1148 242584 1154
rect 242532 1090 242584 1096
rect 242544 814 242572 1090
rect 243280 882 243308 2042
rect 244188 1964 244240 1970
rect 244188 1906 244240 1912
rect 244096 1828 244148 1834
rect 244096 1770 244148 1776
rect 244108 1612 244136 1770
rect 244200 1766 244228 1906
rect 244188 1760 244240 1766
rect 244188 1702 244240 1708
rect 244108 1584 244228 1612
rect 243544 1556 243596 1562
rect 243544 1498 243596 1504
rect 243556 1290 243584 1498
rect 244002 1456 244058 1465
rect 244002 1391 244004 1400
rect 244056 1391 244058 1400
rect 244004 1362 244056 1368
rect 243544 1284 243596 1290
rect 243544 1226 243596 1232
rect 243912 1284 243964 1290
rect 243912 1226 243964 1232
rect 243636 1216 243688 1222
rect 243636 1158 243688 1164
rect 243268 876 243320 882
rect 243268 818 243320 824
rect 232688 808 232740 814
rect 232688 750 232740 756
rect 234344 808 234396 814
rect 234344 750 234396 756
rect 235264 808 235316 814
rect 235264 750 235316 756
rect 235540 808 235592 814
rect 235540 750 235592 756
rect 236000 808 236052 814
rect 236000 750 236052 756
rect 236828 808 236880 814
rect 236828 750 236880 756
rect 237196 808 237248 814
rect 237196 750 237248 756
rect 238024 808 238076 814
rect 238024 750 238076 756
rect 238484 808 238536 814
rect 238484 750 238536 756
rect 239588 808 239640 814
rect 239588 750 239640 756
rect 240048 808 240100 814
rect 240048 750 240100 756
rect 241796 808 241848 814
rect 241796 750 241848 756
rect 242164 808 242216 814
rect 242164 750 242216 756
rect 242532 808 242584 814
rect 242532 750 242584 756
rect 231952 672 232004 678
rect 231952 614 232004 620
rect 243648 513 243676 1158
rect 243820 808 243872 814
rect 243924 796 243952 1226
rect 244002 1184 244058 1193
rect 244200 1170 244228 1584
rect 244292 1562 244320 2586
rect 247052 2582 247080 3062
rect 248432 3058 248460 3334
rect 248420 3052 248472 3058
rect 248420 2994 248472 3000
rect 248052 2644 248104 2650
rect 248052 2586 248104 2592
rect 247040 2576 247092 2582
rect 247040 2518 247092 2524
rect 248064 2446 248092 2586
rect 248052 2440 248104 2446
rect 248052 2382 248104 2388
rect 244372 1964 244424 1970
rect 244372 1906 244424 1912
rect 244280 1556 244332 1562
rect 244280 1498 244332 1504
rect 244278 1456 244334 1465
rect 244278 1391 244334 1400
rect 244292 1222 244320 1391
rect 244384 1306 244412 1906
rect 246488 1692 246540 1698
rect 246488 1634 246540 1640
rect 246304 1624 246356 1630
rect 244830 1592 244886 1601
rect 246304 1566 246356 1572
rect 244830 1527 244886 1536
rect 244844 1426 244872 1527
rect 244832 1420 244884 1426
rect 244832 1362 244884 1368
rect 244556 1352 244608 1358
rect 244554 1320 244556 1329
rect 244608 1320 244610 1329
rect 244384 1278 244504 1306
rect 244002 1119 244004 1128
rect 244056 1119 244058 1128
rect 244108 1142 244228 1170
rect 244280 1216 244332 1222
rect 244280 1158 244332 1164
rect 244004 1090 244056 1096
rect 244108 814 244136 1142
rect 244476 1000 244504 1278
rect 244554 1255 244610 1264
rect 244832 1284 244884 1290
rect 244832 1226 244884 1232
rect 244740 1216 244792 1222
rect 244646 1184 244702 1193
rect 244740 1158 244792 1164
rect 244646 1119 244702 1128
rect 244660 1018 244688 1119
rect 244292 972 244504 1000
rect 244648 1012 244700 1018
rect 244292 898 244320 972
rect 244648 954 244700 960
rect 244200 882 244320 898
rect 244188 876 244320 882
rect 244240 870 244320 876
rect 244464 876 244516 882
rect 244188 818 244240 824
rect 244464 818 244516 824
rect 243872 768 243952 796
rect 244096 808 244148 814
rect 243820 750 243872 756
rect 244096 750 244148 756
rect 244476 513 244504 818
rect 244556 808 244608 814
rect 244752 796 244780 1158
rect 244844 1154 244872 1226
rect 244832 1148 244884 1154
rect 244832 1090 244884 1096
rect 244924 1148 244976 1154
rect 244924 1090 244976 1096
rect 244936 814 244964 1090
rect 244608 768 244780 796
rect 244924 808 244976 814
rect 244556 750 244608 756
rect 244924 750 244976 756
rect 243634 504 243690 513
rect 243634 439 243690 448
rect 244462 504 244518 513
rect 244462 439 244518 448
rect 245384 400 245436 406
rect 245436 348 246160 354
rect 245384 342 246160 348
rect 245396 338 246160 342
rect 245396 332 246172 338
rect 245396 326 246120 332
rect 246120 274 246172 280
rect 246316 270 246344 1566
rect 246500 1494 246528 1634
rect 246488 1488 246540 1494
rect 248432 1465 248460 2994
rect 249168 2650 249196 6802
rect 256589 6784 256601 6840
rect 256657 6784 256681 6840
rect 256737 6784 256761 6840
rect 256817 6784 256841 6840
rect 256897 6784 256909 6840
rect 256589 6010 256909 6784
rect 256589 5958 256595 6010
rect 256647 5958 256659 6010
rect 256711 5958 256723 6010
rect 256775 5958 256787 6010
rect 256839 5958 256851 6010
rect 256903 5958 256909 6010
rect 256589 5721 256909 5958
rect 256589 5665 256601 5721
rect 256657 5665 256681 5721
rect 256737 5665 256761 5721
rect 256817 5665 256841 5721
rect 256897 5665 256909 5721
rect 256589 5641 256909 5665
rect 256589 5585 256601 5641
rect 256657 5585 256681 5641
rect 256737 5585 256761 5641
rect 256817 5585 256841 5641
rect 256897 5585 256909 5641
rect 256589 5561 256909 5585
rect 256589 5505 256601 5561
rect 256657 5505 256681 5561
rect 256737 5505 256761 5561
rect 256817 5505 256841 5561
rect 256897 5505 256909 5561
rect 256589 5481 256909 5505
rect 256589 5425 256601 5481
rect 256657 5425 256681 5481
rect 256737 5425 256761 5481
rect 256817 5425 256841 5481
rect 256897 5425 256909 5481
rect 256589 4922 256909 5425
rect 256589 4870 256595 4922
rect 256647 4870 256659 4922
rect 256711 4870 256723 4922
rect 256775 4870 256787 4922
rect 256839 4870 256851 4922
rect 256903 4870 256909 4922
rect 256589 4362 256909 4870
rect 256589 4306 256601 4362
rect 256657 4306 256681 4362
rect 256737 4306 256761 4362
rect 256817 4306 256841 4362
rect 256897 4306 256909 4362
rect 256589 4282 256909 4306
rect 256589 4226 256601 4282
rect 256657 4226 256681 4282
rect 256737 4226 256761 4282
rect 256817 4226 256841 4282
rect 256897 4226 256909 4282
rect 256589 4202 256909 4226
rect 256589 4146 256601 4202
rect 256657 4146 256681 4202
rect 256737 4146 256761 4202
rect 256817 4146 256841 4202
rect 256897 4146 256909 4202
rect 256589 4122 256909 4146
rect 256589 4066 256601 4122
rect 256657 4066 256681 4122
rect 256737 4066 256761 4122
rect 256817 4066 256841 4122
rect 256897 4066 256909 4122
rect 256589 3834 256909 4066
rect 256589 3782 256595 3834
rect 256647 3782 256659 3834
rect 256711 3782 256723 3834
rect 256775 3782 256787 3834
rect 256839 3782 256851 3834
rect 256903 3782 256909 3834
rect 256589 3003 256909 3782
rect 249708 2984 249760 2990
rect 249708 2926 249760 2932
rect 256589 2947 256601 3003
rect 256657 2947 256681 3003
rect 256737 2947 256761 3003
rect 256817 2947 256841 3003
rect 256897 2947 256909 3003
rect 249248 2848 249300 2854
rect 249248 2790 249300 2796
rect 249156 2644 249208 2650
rect 249156 2586 249208 2592
rect 249260 2582 249288 2790
rect 249248 2576 249300 2582
rect 249248 2518 249300 2524
rect 249720 1902 249748 2926
rect 256589 2923 256909 2947
rect 256589 2867 256601 2923
rect 256657 2867 256681 2923
rect 256737 2867 256761 2923
rect 256817 2867 256841 2923
rect 256897 2867 256909 2923
rect 256589 2843 256909 2867
rect 256589 2787 256601 2843
rect 256657 2787 256681 2843
rect 256737 2787 256761 2843
rect 256817 2787 256841 2843
rect 256897 2787 256909 2843
rect 256589 2763 256909 2787
rect 256589 2746 256601 2763
rect 256657 2746 256681 2763
rect 256737 2746 256761 2763
rect 256817 2746 256841 2763
rect 256897 2746 256909 2763
rect 256589 2694 256595 2746
rect 256657 2707 256659 2746
rect 256839 2707 256841 2746
rect 256647 2694 256659 2707
rect 256711 2694 256723 2707
rect 256775 2694 256787 2707
rect 256839 2694 256851 2707
rect 256903 2694 256909 2746
rect 250444 2372 250496 2378
rect 250444 2314 250496 2320
rect 249708 1896 249760 1902
rect 249708 1838 249760 1844
rect 249430 1728 249486 1737
rect 249430 1663 249486 1672
rect 246488 1430 246540 1436
rect 248418 1456 248474 1465
rect 248418 1391 248474 1400
rect 249444 1358 249472 1663
rect 250456 1494 250484 2314
rect 250444 1488 250496 1494
rect 250444 1430 250496 1436
rect 249432 1352 249484 1358
rect 246394 1320 246450 1329
rect 249432 1294 249484 1300
rect 246394 1255 246450 1264
rect 224132 206 224184 212
rect 227732 202 227852 218
rect 245844 264 245896 270
rect 246304 264 246356 270
rect 245896 224 246068 252
rect 245844 206 245896 212
rect 246040 218 246068 224
rect 202972 196 203024 202
rect 202972 138 203024 144
rect 227720 196 227852 202
rect 227772 190 227852 196
rect 246040 202 246160 218
rect 246304 206 246356 212
rect 246040 196 246172 202
rect 246040 190 246120 196
rect 227720 138 227772 144
rect 246120 138 246172 144
rect 246408 134 246436 1255
rect 249156 1216 249208 1222
rect 249156 1158 249208 1164
rect 249168 610 249196 1158
rect 249340 1148 249392 1154
rect 249340 1090 249392 1096
rect 249156 604 249208 610
rect 249156 546 249208 552
rect 249352 474 249380 1090
rect 256589 964 256909 2694
rect 256589 908 256601 964
rect 256657 908 256681 964
rect 256737 908 256761 964
rect 256817 908 256841 964
rect 256897 908 256909 964
rect 256589 884 256909 908
rect 256589 828 256601 884
rect 256657 828 256681 884
rect 256737 828 256761 884
rect 256817 828 256841 884
rect 256897 828 256909 884
rect 256589 804 256909 828
rect 256589 748 256601 804
rect 256657 748 256681 804
rect 256737 748 256761 804
rect 256817 748 256841 804
rect 256897 748 256909 804
rect 256589 724 256909 748
rect 256589 668 256601 724
rect 256657 668 256681 724
rect 256737 668 256761 724
rect 256817 668 256841 724
rect 256897 668 256909 724
rect 249340 468 249392 474
rect 249340 410 249392 416
rect 246396 128 246448 134
rect 246396 70 246448 76
rect 86819 8 86831 64
rect 86887 8 86911 64
rect 86967 8 86991 64
rect 87047 8 87071 64
rect 87127 8 87139 64
rect 86819 -4 87139 8
rect 191380 60 191432 66
rect 191380 2 191432 8
rect 256589 -4 256909 668
rect 257249 9784 257569 9796
rect 257249 9728 257261 9784
rect 257317 9728 257341 9784
rect 257397 9728 257421 9784
rect 257477 9728 257501 9784
rect 257557 9728 257569 9784
rect 257249 9704 257569 9728
rect 257249 9648 257261 9704
rect 257317 9648 257341 9704
rect 257397 9648 257421 9704
rect 257477 9648 257501 9704
rect 257557 9648 257569 9704
rect 257249 9624 257569 9648
rect 257249 9568 257261 9624
rect 257317 9568 257341 9624
rect 257397 9568 257421 9624
rect 257477 9568 257501 9624
rect 257557 9568 257569 9624
rect 257249 9544 257569 9568
rect 257249 9488 257261 9544
rect 257317 9488 257341 9544
rect 257397 9488 257421 9544
rect 257477 9488 257501 9544
rect 257557 9488 257569 9544
rect 257249 7740 257569 9488
rect 260472 9240 260524 9246
rect 260472 9182 260524 9188
rect 275928 9240 275980 9246
rect 275928 9182 275980 9188
rect 321468 9240 321520 9246
rect 321468 9182 321520 9188
rect 336832 9240 336884 9246
rect 336832 9182 336884 9188
rect 368388 9240 368440 9246
rect 368388 9182 368440 9188
rect 383568 9240 383620 9246
rect 383568 9182 383620 9188
rect 413928 9240 413980 9246
rect 413928 9182 413980 9188
rect 257249 7684 257261 7740
rect 257317 7684 257341 7740
rect 257397 7684 257421 7740
rect 257477 7684 257501 7740
rect 257557 7684 257569 7740
rect 257249 7660 257569 7684
rect 257249 7642 257261 7660
rect 257317 7642 257341 7660
rect 257397 7642 257421 7660
rect 257477 7642 257501 7660
rect 257557 7642 257569 7660
rect 257249 7590 257255 7642
rect 257317 7604 257319 7642
rect 257499 7604 257501 7642
rect 257307 7590 257319 7604
rect 257371 7590 257383 7604
rect 257435 7590 257447 7604
rect 257499 7590 257511 7604
rect 257563 7590 257569 7642
rect 257249 7580 257569 7590
rect 257249 7524 257261 7580
rect 257317 7524 257341 7580
rect 257397 7524 257421 7580
rect 257477 7524 257501 7580
rect 257557 7524 257569 7580
rect 257249 7500 257569 7524
rect 257249 7444 257261 7500
rect 257317 7444 257341 7500
rect 257397 7444 257421 7500
rect 257477 7444 257501 7500
rect 257557 7444 257569 7500
rect 257249 6554 257569 7444
rect 260484 6866 260512 9182
rect 275940 6866 275968 9182
rect 291108 8968 291160 8974
rect 291108 8910 291160 8916
rect 306288 8968 306340 8974
rect 306288 8910 306340 8916
rect 291120 6866 291148 8910
rect 260472 6860 260524 6866
rect 260472 6802 260524 6808
rect 264336 6860 264388 6866
rect 264336 6802 264388 6808
rect 275928 6860 275980 6866
rect 275928 6802 275980 6808
rect 280068 6860 280120 6866
rect 280068 6802 280120 6808
rect 291108 6860 291160 6866
rect 291108 6802 291160 6808
rect 295524 6860 295576 6866
rect 295524 6802 295576 6808
rect 257249 6502 257255 6554
rect 257307 6502 257319 6554
rect 257371 6502 257383 6554
rect 257435 6502 257447 6554
rect 257499 6502 257511 6554
rect 257563 6502 257569 6554
rect 257249 6381 257569 6502
rect 257249 6325 257261 6381
rect 257317 6325 257341 6381
rect 257397 6325 257421 6381
rect 257477 6325 257501 6381
rect 257557 6325 257569 6381
rect 257249 6301 257569 6325
rect 257249 6245 257261 6301
rect 257317 6245 257341 6301
rect 257397 6245 257421 6301
rect 257477 6245 257501 6301
rect 257557 6245 257569 6301
rect 257249 6221 257569 6245
rect 257249 6165 257261 6221
rect 257317 6165 257341 6221
rect 257397 6165 257421 6221
rect 257477 6165 257501 6221
rect 257557 6165 257569 6221
rect 257249 6141 257569 6165
rect 257249 6085 257261 6141
rect 257317 6085 257341 6141
rect 257397 6085 257421 6141
rect 257477 6085 257501 6141
rect 257557 6085 257569 6141
rect 257249 5466 257569 6085
rect 257249 5414 257255 5466
rect 257307 5414 257319 5466
rect 257371 5414 257383 5466
rect 257435 5414 257447 5466
rect 257499 5414 257511 5466
rect 257563 5414 257569 5466
rect 257249 5022 257569 5414
rect 257249 4966 257261 5022
rect 257317 4966 257341 5022
rect 257397 4966 257421 5022
rect 257477 4966 257501 5022
rect 257557 4966 257569 5022
rect 257249 4942 257569 4966
rect 257249 4886 257261 4942
rect 257317 4886 257341 4942
rect 257397 4886 257421 4942
rect 257477 4886 257501 4942
rect 257557 4886 257569 4942
rect 257249 4862 257569 4886
rect 257249 4806 257261 4862
rect 257317 4806 257341 4862
rect 257397 4806 257421 4862
rect 257477 4806 257501 4862
rect 257557 4806 257569 4862
rect 257249 4782 257569 4806
rect 257249 4726 257261 4782
rect 257317 4726 257341 4782
rect 257397 4726 257421 4782
rect 257477 4726 257501 4782
rect 257557 4726 257569 4782
rect 257249 4378 257569 4726
rect 257249 4326 257255 4378
rect 257307 4326 257319 4378
rect 257371 4326 257383 4378
rect 257435 4326 257447 4378
rect 257499 4326 257511 4378
rect 257563 4326 257569 4378
rect 257249 3663 257569 4326
rect 257249 3607 257261 3663
rect 257317 3607 257341 3663
rect 257397 3607 257421 3663
rect 257477 3607 257501 3663
rect 257557 3607 257569 3663
rect 257249 3583 257569 3607
rect 257249 3527 257261 3583
rect 257317 3527 257341 3583
rect 257397 3527 257421 3583
rect 257477 3527 257501 3583
rect 257557 3527 257569 3583
rect 257249 3503 257569 3527
rect 257249 3447 257261 3503
rect 257317 3447 257341 3503
rect 257397 3447 257421 3503
rect 257477 3447 257501 3503
rect 257557 3447 257569 3503
rect 257249 3423 257569 3447
rect 257249 3367 257261 3423
rect 257317 3367 257341 3423
rect 257397 3367 257421 3423
rect 257477 3367 257501 3423
rect 257557 3367 257569 3423
rect 257249 3290 257569 3367
rect 257249 3238 257255 3290
rect 257307 3238 257319 3290
rect 257371 3238 257383 3290
rect 257435 3238 257447 3290
rect 257499 3238 257511 3290
rect 257563 3238 257569 3290
rect 257249 2202 257569 3238
rect 264348 3058 264376 6802
rect 264336 3052 264388 3058
rect 264336 2994 264388 3000
rect 264348 2446 264376 2994
rect 277216 2848 277268 2854
rect 277216 2790 277268 2796
rect 273352 2644 273404 2650
rect 273352 2586 273404 2592
rect 273364 2446 273392 2586
rect 277228 2446 277256 2790
rect 264336 2440 264388 2446
rect 264336 2382 264388 2388
rect 273352 2440 273404 2446
rect 273352 2382 273404 2388
rect 276020 2440 276072 2446
rect 276020 2382 276072 2388
rect 277216 2440 277268 2446
rect 277216 2382 277268 2388
rect 275560 2372 275612 2378
rect 275560 2314 275612 2320
rect 264612 2304 264664 2310
rect 264612 2246 264664 2252
rect 272524 2304 272576 2310
rect 272524 2246 272576 2252
rect 274732 2304 274784 2310
rect 274732 2246 274784 2252
rect 257249 2150 257255 2202
rect 257307 2150 257319 2202
rect 257371 2150 257383 2202
rect 257435 2150 257447 2202
rect 257499 2150 257511 2202
rect 257563 2150 257569 2202
rect 257249 304 257569 2150
rect 257249 248 257261 304
rect 257317 248 257341 304
rect 257397 248 257421 304
rect 257477 248 257501 304
rect 257557 248 257569 304
rect 264624 270 264652 2246
rect 272536 338 272564 2246
rect 274744 2106 274772 2246
rect 274732 2100 274784 2106
rect 274732 2042 274784 2048
rect 275572 1630 275600 2314
rect 276032 1698 276060 2382
rect 277676 2372 277728 2378
rect 277676 2314 277728 2320
rect 277688 1902 277716 2314
rect 280080 2310 280108 6802
rect 292856 2848 292908 2854
rect 292856 2790 292908 2796
rect 292868 2446 292896 2790
rect 295536 2650 295564 6802
rect 306300 6186 306328 8910
rect 321480 6866 321508 9182
rect 336844 6866 336872 9182
rect 353208 8900 353260 8906
rect 353208 8842 353260 8848
rect 353220 6866 353248 8842
rect 368400 6866 368428 9182
rect 321468 6860 321520 6866
rect 321468 6802 321520 6808
rect 326436 6860 326488 6866
rect 326436 6802 326488 6808
rect 336832 6860 336884 6866
rect 336832 6802 336884 6808
rect 341892 6860 341944 6866
rect 341892 6802 341944 6808
rect 353208 6860 353260 6866
rect 353208 6802 353260 6808
rect 357072 6860 357124 6866
rect 357072 6802 357124 6808
rect 368388 6860 368440 6866
rect 368388 6802 368440 6808
rect 372804 6860 372856 6866
rect 372804 6802 372856 6808
rect 306288 6180 306340 6186
rect 306288 6122 306340 6128
rect 310704 6180 310756 6186
rect 310704 6122 310756 6128
rect 310716 3058 310744 6122
rect 310704 3052 310756 3058
rect 310704 2994 310756 3000
rect 295524 2644 295576 2650
rect 295524 2586 295576 2592
rect 295800 2508 295852 2514
rect 295800 2450 295852 2456
rect 292856 2440 292908 2446
rect 292856 2382 292908 2388
rect 294420 2440 294472 2446
rect 295812 2394 295840 2450
rect 310716 2446 310744 2994
rect 323584 2848 323636 2854
rect 323584 2790 323636 2796
rect 324504 2848 324556 2854
rect 324504 2790 324556 2796
rect 326160 2848 326212 2854
rect 326160 2790 326212 2796
rect 323596 2446 323624 2790
rect 324516 2446 324544 2790
rect 326172 2553 326200 2790
rect 326158 2544 326214 2553
rect 326158 2479 326214 2488
rect 326172 2446 326200 2479
rect 294420 2382 294472 2388
rect 290188 2372 290240 2378
rect 290188 2314 290240 2320
rect 290924 2372 290976 2378
rect 290924 2314 290976 2320
rect 278964 2304 279016 2310
rect 278964 2246 279016 2252
rect 280068 2304 280120 2310
rect 280068 2246 280120 2252
rect 287980 2304 288032 2310
rect 287980 2246 288032 2252
rect 278976 2038 279004 2246
rect 278964 2032 279016 2038
rect 278964 1974 279016 1980
rect 277676 1896 277728 1902
rect 277676 1838 277728 1844
rect 276020 1692 276072 1698
rect 276020 1634 276072 1640
rect 275560 1624 275612 1630
rect 275560 1566 275612 1572
rect 272524 332 272576 338
rect 272524 274 272576 280
rect 257249 224 257569 248
rect 257249 168 257261 224
rect 257317 168 257341 224
rect 257397 168 257421 224
rect 257477 168 257501 224
rect 257557 168 257569 224
rect 264612 264 264664 270
rect 264612 206 264664 212
rect 287992 202 288020 2246
rect 290200 1970 290228 2314
rect 290936 2106 290964 2314
rect 290924 2100 290976 2106
rect 290924 2042 290976 2048
rect 290188 1964 290240 1970
rect 290188 1906 290240 1912
rect 292868 1562 292896 2382
rect 293408 2372 293460 2378
rect 293408 2314 293460 2320
rect 293420 1970 293448 2314
rect 293408 1964 293460 1970
rect 293408 1906 293460 1912
rect 294432 1766 294460 2382
rect 295628 2366 295840 2394
rect 310704 2440 310756 2446
rect 310704 2382 310756 2388
rect 320916 2440 320968 2446
rect 320916 2382 320968 2388
rect 323584 2440 323636 2446
rect 323584 2382 323636 2388
rect 324504 2440 324556 2446
rect 324504 2382 324556 2388
rect 326160 2440 326212 2446
rect 326160 2382 326212 2388
rect 295628 2310 295656 2366
rect 320928 2310 320956 2382
rect 322112 2372 322164 2378
rect 322112 2314 322164 2320
rect 295616 2304 295668 2310
rect 295616 2246 295668 2252
rect 310980 2304 311032 2310
rect 310980 2246 311032 2252
rect 320916 2304 320968 2310
rect 320916 2246 320968 2252
rect 294420 1760 294472 1766
rect 294420 1702 294472 1708
rect 292856 1556 292908 1562
rect 292856 1498 292908 1504
rect 257249 144 257569 168
rect 257249 88 257261 144
rect 257317 88 257341 144
rect 257397 88 257421 144
rect 257477 88 257501 144
rect 257557 88 257569 144
rect 287980 196 288032 202
rect 287980 138 288032 144
rect 310992 134 311020 2246
rect 320928 1834 320956 2246
rect 322124 2038 322152 2314
rect 322112 2032 322164 2038
rect 322112 1974 322164 1980
rect 320916 1828 320968 1834
rect 320916 1770 320968 1776
rect 323596 1426 323624 2382
rect 324136 2372 324188 2378
rect 324136 2314 324188 2320
rect 325332 2372 325384 2378
rect 325332 2314 325384 2320
rect 324148 1698 324176 2314
rect 324136 1692 324188 1698
rect 324136 1634 324188 1640
rect 325344 1562 325372 2314
rect 326448 2310 326476 6802
rect 339592 3528 339644 3534
rect 339592 3470 339644 3476
rect 337384 3460 337436 3466
rect 337384 3402 337436 3408
rect 336464 3392 336516 3398
rect 336464 3334 336516 3340
rect 331588 2848 331640 2854
rect 331588 2790 331640 2796
rect 333060 2848 333112 2854
rect 333060 2790 333112 2796
rect 334624 2848 334676 2854
rect 334624 2790 334676 2796
rect 335728 2848 335780 2854
rect 335728 2790 335780 2796
rect 331600 2446 331628 2790
rect 333072 2446 333100 2790
rect 334636 2446 334664 2790
rect 335740 2446 335768 2790
rect 336476 2446 336504 3334
rect 337396 3058 337424 3402
rect 338212 3392 338264 3398
rect 338212 3334 338264 3340
rect 337384 3052 337436 3058
rect 337384 2994 337436 3000
rect 336832 2984 336884 2990
rect 336832 2926 336884 2932
rect 331588 2440 331640 2446
rect 331588 2382 331640 2388
rect 333060 2440 333112 2446
rect 333060 2382 333112 2388
rect 334624 2440 334676 2446
rect 334624 2382 334676 2388
rect 335728 2440 335780 2446
rect 335728 2382 335780 2388
rect 336464 2440 336516 2446
rect 336464 2382 336516 2388
rect 331312 2372 331364 2378
rect 331312 2314 331364 2320
rect 326436 2304 326488 2310
rect 326436 2246 326488 2252
rect 325332 1556 325384 1562
rect 325332 1498 325384 1504
rect 323584 1420 323636 1426
rect 323584 1362 323636 1368
rect 331324 1290 331352 2314
rect 331600 1766 331628 2382
rect 332600 2372 332652 2378
rect 332600 2314 332652 2320
rect 331588 1760 331640 1766
rect 331588 1702 331640 1708
rect 331312 1284 331364 1290
rect 331312 1226 331364 1232
rect 332612 1086 332640 2314
rect 333072 1086 333100 2382
rect 334072 2372 334124 2378
rect 334072 2314 334124 2320
rect 332600 1080 332652 1086
rect 332600 1022 332652 1028
rect 333060 1080 333112 1086
rect 333060 1022 333112 1028
rect 334084 882 334112 2314
rect 334636 1222 334664 2382
rect 335452 2372 335504 2378
rect 335452 2314 335504 2320
rect 334624 1216 334676 1222
rect 334624 1158 334676 1164
rect 335464 950 335492 2314
rect 335740 1290 335768 2382
rect 335728 1284 335780 1290
rect 335728 1226 335780 1232
rect 335452 944 335504 950
rect 335452 886 335504 892
rect 334072 876 334124 882
rect 334072 818 334124 824
rect 336476 610 336504 2382
rect 336844 1018 336872 2926
rect 338224 2446 338252 3334
rect 339604 3058 339632 3470
rect 339868 3392 339920 3398
rect 339868 3334 339920 3340
rect 339592 3052 339644 3058
rect 339592 2994 339644 3000
rect 339880 2446 339908 3334
rect 341524 2984 341576 2990
rect 341524 2926 341576 2932
rect 340236 2848 340288 2854
rect 340236 2790 340288 2796
rect 340248 2446 340276 2790
rect 338212 2440 338264 2446
rect 337014 2408 337070 2417
rect 338212 2382 338264 2388
rect 339868 2440 339920 2446
rect 339868 2382 339920 2388
rect 340236 2440 340288 2446
rect 340236 2382 340288 2388
rect 337014 2343 337016 2352
rect 337068 2343 337070 2352
rect 337660 2372 337712 2378
rect 337016 2314 337068 2320
rect 337660 2314 337712 2320
rect 337672 1154 337700 2314
rect 338224 1358 338252 2382
rect 339040 2372 339092 2378
rect 339040 2314 339092 2320
rect 338212 1352 338264 1358
rect 338212 1294 338264 1300
rect 337660 1148 337712 1154
rect 337660 1090 337712 1096
rect 336832 1012 336884 1018
rect 336832 954 336884 960
rect 336464 604 336516 610
rect 336464 546 336516 552
rect 339052 474 339080 2314
rect 340248 1494 340276 2382
rect 340788 2372 340840 2378
rect 340788 2314 340840 2320
rect 340236 1488 340288 1494
rect 340236 1430 340288 1436
rect 340800 1426 340828 2314
rect 340788 1420 340840 1426
rect 340788 1362 340840 1368
rect 339040 468 339092 474
rect 339040 410 339092 416
rect 257249 64 257569 88
rect 310980 128 311032 134
rect 310980 70 311032 76
rect 341536 66 341564 2926
rect 341904 2310 341932 6802
rect 357084 3194 357112 6802
rect 357072 3188 357124 3194
rect 357072 3130 357124 3136
rect 342720 3052 342772 3058
rect 342720 2994 342772 3000
rect 342732 2854 342760 2994
rect 342720 2848 342772 2854
rect 342720 2790 342772 2796
rect 341892 2304 341944 2310
rect 341892 2246 341944 2252
rect 342732 1834 342760 2790
rect 357084 2446 357112 3130
rect 367468 2848 367520 2854
rect 367468 2790 367520 2796
rect 370872 2848 370924 2854
rect 370872 2790 370924 2796
rect 367480 2650 367508 2790
rect 367468 2644 367520 2650
rect 367468 2586 367520 2592
rect 367480 2446 367508 2586
rect 370884 2446 370912 2790
rect 372816 2582 372844 6802
rect 383580 6186 383608 9182
rect 398748 8900 398800 8906
rect 398748 8842 398800 8848
rect 398760 6866 398788 8842
rect 413940 6866 413968 9182
rect 427019 9124 427339 9796
rect 427019 9068 427031 9124
rect 427087 9068 427111 9124
rect 427167 9068 427191 9124
rect 427247 9068 427271 9124
rect 427327 9068 427339 9124
rect 427019 9044 427339 9068
rect 427019 8988 427031 9044
rect 427087 8988 427111 9044
rect 427167 8988 427191 9044
rect 427247 8988 427271 9044
rect 427327 8988 427339 9044
rect 427019 8964 427339 8988
rect 427019 8908 427031 8964
rect 427087 8908 427111 8964
rect 427167 8908 427191 8964
rect 427247 8908 427271 8964
rect 427327 8908 427339 8964
rect 427019 8884 427339 8908
rect 427019 8828 427031 8884
rect 427087 8828 427111 8884
rect 427167 8828 427191 8884
rect 427247 8828 427271 8884
rect 427327 8828 427339 8884
rect 427019 7098 427339 8828
rect 427019 7046 427025 7098
rect 427077 7080 427089 7098
rect 427141 7080 427153 7098
rect 427205 7080 427217 7098
rect 427269 7080 427281 7098
rect 427087 7046 427089 7080
rect 427269 7046 427271 7080
rect 427333 7046 427339 7098
rect 427019 7024 427031 7046
rect 427087 7024 427111 7046
rect 427167 7024 427191 7046
rect 427247 7024 427271 7046
rect 427327 7024 427339 7046
rect 427019 7000 427339 7024
rect 427019 6944 427031 7000
rect 427087 6944 427111 7000
rect 427167 6944 427191 7000
rect 427247 6944 427271 7000
rect 427327 6944 427339 7000
rect 427019 6920 427339 6944
rect 398748 6860 398800 6866
rect 398748 6802 398800 6808
rect 403440 6860 403492 6866
rect 403440 6802 403492 6808
rect 413928 6860 413980 6866
rect 413928 6802 413980 6808
rect 419172 6860 419224 6866
rect 419172 6802 419224 6808
rect 427019 6864 427031 6920
rect 427087 6864 427111 6920
rect 427167 6864 427191 6920
rect 427247 6864 427271 6920
rect 427327 6864 427339 6920
rect 427019 6840 427339 6864
rect 383568 6180 383620 6186
rect 383568 6122 383620 6128
rect 388260 6180 388312 6186
rect 388260 6122 388312 6128
rect 372988 2916 373040 2922
rect 372988 2858 373040 2864
rect 372804 2576 372856 2582
rect 372804 2518 372856 2524
rect 373000 2446 373028 2858
rect 382832 2848 382884 2854
rect 382832 2790 382884 2796
rect 386604 2848 386656 2854
rect 386604 2790 386656 2796
rect 357072 2440 357124 2446
rect 357072 2382 357124 2388
rect 367468 2440 367520 2446
rect 367468 2382 367520 2388
rect 370320 2440 370372 2446
rect 370320 2382 370372 2388
rect 370872 2440 370924 2446
rect 370872 2382 370924 2388
rect 372988 2440 373040 2446
rect 372988 2382 373040 2388
rect 368296 2372 368348 2378
rect 368296 2314 368348 2320
rect 357348 2304 357400 2310
rect 357348 2246 357400 2252
rect 342720 1828 342772 1834
rect 342720 1770 342772 1776
rect 357360 1766 357388 2246
rect 357348 1760 357400 1766
rect 357348 1702 357400 1708
rect 368308 1154 368336 2314
rect 369124 2304 369176 2310
rect 369124 2246 369176 2252
rect 369136 1630 369164 2246
rect 370332 1902 370360 2382
rect 382844 2378 382872 2790
rect 386616 2446 386644 2790
rect 388272 2582 388300 6122
rect 403452 3194 403480 6802
rect 403440 3188 403492 3194
rect 403440 3130 403492 3136
rect 388444 3120 388496 3126
rect 388444 3062 388496 3068
rect 388260 2576 388312 2582
rect 388260 2518 388312 2524
rect 388456 2446 388484 3062
rect 403452 2446 403480 3130
rect 417516 2848 417568 2854
rect 417516 2790 417568 2796
rect 418896 2848 418948 2854
rect 418896 2790 418948 2796
rect 417528 2446 417556 2790
rect 418908 2446 418936 2790
rect 386604 2440 386656 2446
rect 386604 2382 386656 2388
rect 388444 2440 388496 2446
rect 388444 2382 388496 2388
rect 403440 2440 403492 2446
rect 403440 2382 403492 2388
rect 417516 2440 417568 2446
rect 417516 2382 417568 2388
rect 418896 2440 418948 2446
rect 418896 2382 418948 2388
rect 370412 2372 370464 2378
rect 370412 2314 370464 2320
rect 382832 2372 382884 2378
rect 382832 2314 382884 2320
rect 383660 2372 383712 2378
rect 383660 2314 383712 2320
rect 370424 1902 370452 2314
rect 370320 1896 370372 1902
rect 370320 1838 370372 1844
rect 370412 1896 370464 1902
rect 370412 1838 370464 1844
rect 383672 1630 383700 2314
rect 384580 2304 384632 2310
rect 384580 2246 384632 2252
rect 384592 2106 384620 2246
rect 384580 2100 384632 2106
rect 384580 2042 384632 2048
rect 386616 1970 386644 2382
rect 387156 2372 387208 2378
rect 387156 2314 387208 2320
rect 416780 2372 416832 2378
rect 416780 2314 416832 2320
rect 386604 1964 386656 1970
rect 386604 1906 386656 1912
rect 369124 1624 369176 1630
rect 369124 1566 369176 1572
rect 383660 1624 383712 1630
rect 383660 1566 383712 1572
rect 387168 1494 387196 2314
rect 403716 2304 403768 2310
rect 403716 2246 403768 2252
rect 415492 2304 415544 2310
rect 415492 2246 415544 2252
rect 387156 1488 387208 1494
rect 387156 1430 387208 1436
rect 368296 1148 368348 1154
rect 368296 1090 368348 1096
rect 403728 1086 403756 2246
rect 415504 2038 415532 2246
rect 416792 2106 416820 2314
rect 416780 2100 416832 2106
rect 416780 2042 416832 2048
rect 415492 2032 415544 2038
rect 415492 1974 415544 1980
rect 417528 1698 417556 2382
rect 417516 1692 417568 1698
rect 417516 1634 417568 1640
rect 418908 1562 418936 2382
rect 419184 2310 419212 6802
rect 427019 6784 427031 6840
rect 427087 6784 427111 6840
rect 427167 6784 427191 6840
rect 427247 6784 427271 6840
rect 427327 6784 427339 6840
rect 427019 6010 427339 6784
rect 427019 5958 427025 6010
rect 427077 5958 427089 6010
rect 427141 5958 427153 6010
rect 427205 5958 427217 6010
rect 427269 5958 427281 6010
rect 427333 5958 427339 6010
rect 427019 5721 427339 5958
rect 427019 5665 427031 5721
rect 427087 5665 427111 5721
rect 427167 5665 427191 5721
rect 427247 5665 427271 5721
rect 427327 5665 427339 5721
rect 427019 5641 427339 5665
rect 427019 5585 427031 5641
rect 427087 5585 427111 5641
rect 427167 5585 427191 5641
rect 427247 5585 427271 5641
rect 427327 5585 427339 5641
rect 427019 5561 427339 5585
rect 427019 5505 427031 5561
rect 427087 5505 427111 5561
rect 427167 5505 427191 5561
rect 427247 5505 427271 5561
rect 427327 5505 427339 5561
rect 427019 5481 427339 5505
rect 427019 5425 427031 5481
rect 427087 5425 427111 5481
rect 427167 5425 427191 5481
rect 427247 5425 427271 5481
rect 427327 5425 427339 5481
rect 427019 4922 427339 5425
rect 427019 4870 427025 4922
rect 427077 4870 427089 4922
rect 427141 4870 427153 4922
rect 427205 4870 427217 4922
rect 427269 4870 427281 4922
rect 427333 4870 427339 4922
rect 427019 4362 427339 4870
rect 427019 4306 427031 4362
rect 427087 4306 427111 4362
rect 427167 4306 427191 4362
rect 427247 4306 427271 4362
rect 427327 4306 427339 4362
rect 427019 4282 427339 4306
rect 427019 4226 427031 4282
rect 427087 4226 427111 4282
rect 427167 4226 427191 4282
rect 427247 4226 427271 4282
rect 427327 4226 427339 4282
rect 427019 4202 427339 4226
rect 427019 4146 427031 4202
rect 427087 4146 427111 4202
rect 427167 4146 427191 4202
rect 427247 4146 427271 4202
rect 427327 4146 427339 4202
rect 427019 4122 427339 4146
rect 427019 4066 427031 4122
rect 427087 4066 427111 4122
rect 427167 4066 427191 4122
rect 427247 4066 427271 4122
rect 427327 4066 427339 4122
rect 427019 3834 427339 4066
rect 427019 3782 427025 3834
rect 427077 3782 427089 3834
rect 427141 3782 427153 3834
rect 427205 3782 427217 3834
rect 427269 3782 427281 3834
rect 427333 3782 427339 3834
rect 426900 3392 426952 3398
rect 426900 3334 426952 3340
rect 426912 3194 426940 3334
rect 426900 3188 426952 3194
rect 426900 3130 426952 3136
rect 427019 3003 427339 3782
rect 427019 2947 427031 3003
rect 427087 2947 427111 3003
rect 427167 2947 427191 3003
rect 427247 2947 427271 3003
rect 427327 2947 427339 3003
rect 427019 2923 427339 2947
rect 427019 2867 427031 2923
rect 427087 2867 427111 2923
rect 427167 2867 427191 2923
rect 427247 2867 427271 2923
rect 427327 2867 427339 2923
rect 427019 2843 427339 2867
rect 427019 2787 427031 2843
rect 427087 2787 427111 2843
rect 427167 2787 427191 2843
rect 427247 2787 427271 2843
rect 427327 2787 427339 2843
rect 427019 2763 427339 2787
rect 427019 2746 427031 2763
rect 427087 2746 427111 2763
rect 427167 2746 427191 2763
rect 427247 2746 427271 2763
rect 427327 2746 427339 2763
rect 427019 2694 427025 2746
rect 427087 2707 427089 2746
rect 427269 2707 427271 2746
rect 427077 2694 427089 2707
rect 427141 2694 427153 2707
rect 427205 2694 427217 2707
rect 427269 2694 427281 2707
rect 427333 2694 427339 2746
rect 419172 2304 419224 2310
rect 419172 2246 419224 2252
rect 418896 1556 418948 1562
rect 418896 1498 418948 1504
rect 403716 1080 403768 1086
rect 403716 1022 403768 1028
rect 427019 964 427339 2694
rect 427019 908 427031 964
rect 427087 908 427111 964
rect 427167 908 427191 964
rect 427247 908 427271 964
rect 427327 908 427339 964
rect 427019 884 427339 908
rect 427019 828 427031 884
rect 427087 828 427111 884
rect 427167 828 427191 884
rect 427247 828 427271 884
rect 427327 828 427339 884
rect 427019 804 427339 828
rect 427019 748 427031 804
rect 427087 748 427111 804
rect 427167 748 427191 804
rect 427247 748 427271 804
rect 427327 748 427339 804
rect 427019 724 427339 748
rect 427019 668 427031 724
rect 427087 668 427111 724
rect 427167 668 427191 724
rect 427247 668 427271 724
rect 427327 668 427339 724
rect 257249 8 257261 64
rect 257317 8 257341 64
rect 257397 8 257421 64
rect 257477 8 257501 64
rect 257557 8 257569 64
rect 257249 -4 257569 8
rect 341524 60 341576 66
rect 341524 2 341576 8
rect 427019 -4 427339 668
rect 427679 9784 427999 9796
rect 427679 9728 427691 9784
rect 427747 9728 427771 9784
rect 427827 9728 427851 9784
rect 427907 9728 427931 9784
rect 427987 9728 427999 9784
rect 427679 9704 427999 9728
rect 427679 9648 427691 9704
rect 427747 9648 427771 9704
rect 427827 9648 427851 9704
rect 427907 9648 427931 9704
rect 427987 9648 427999 9704
rect 427679 9624 427999 9648
rect 427679 9568 427691 9624
rect 427747 9568 427771 9624
rect 427827 9568 427851 9624
rect 427907 9568 427931 9624
rect 427987 9568 427999 9624
rect 427679 9544 427999 9568
rect 427679 9488 427691 9544
rect 427747 9488 427771 9544
rect 427827 9488 427851 9544
rect 427907 9488 427931 9544
rect 427987 9488 427999 9544
rect 427679 7740 427999 9488
rect 429108 9240 429160 9246
rect 429108 9182 429160 9188
rect 459468 9240 459520 9246
rect 459468 9182 459520 9188
rect 474648 9240 474700 9246
rect 474648 9182 474700 9188
rect 520924 9240 520976 9246
rect 520924 9182 520976 9188
rect 536748 9240 536800 9246
rect 536748 9182 536800 9188
rect 567108 9240 567160 9246
rect 567108 9182 567160 9188
rect 582288 9240 582340 9246
rect 582288 9182 582340 9188
rect 427679 7684 427691 7740
rect 427747 7684 427771 7740
rect 427827 7684 427851 7740
rect 427907 7684 427931 7740
rect 427987 7684 427999 7740
rect 427679 7660 427999 7684
rect 427679 7642 427691 7660
rect 427747 7642 427771 7660
rect 427827 7642 427851 7660
rect 427907 7642 427931 7660
rect 427987 7642 427999 7660
rect 427679 7590 427685 7642
rect 427747 7604 427749 7642
rect 427929 7604 427931 7642
rect 427737 7590 427749 7604
rect 427801 7590 427813 7604
rect 427865 7590 427877 7604
rect 427929 7590 427941 7604
rect 427993 7590 427999 7642
rect 427679 7580 427999 7590
rect 427679 7524 427691 7580
rect 427747 7524 427771 7580
rect 427827 7524 427851 7580
rect 427907 7524 427931 7580
rect 427987 7524 427999 7580
rect 427679 7500 427999 7524
rect 427679 7444 427691 7500
rect 427747 7444 427771 7500
rect 427827 7444 427851 7500
rect 427907 7444 427931 7500
rect 427987 7444 427999 7500
rect 427679 6554 427999 7444
rect 429120 6866 429148 9182
rect 444104 8968 444156 8974
rect 444104 8910 444156 8916
rect 444116 6866 444144 8910
rect 429108 6860 429160 6866
rect 429108 6802 429160 6808
rect 434628 6860 434680 6866
rect 434628 6802 434680 6808
rect 444104 6860 444156 6866
rect 444104 6802 444156 6808
rect 449900 6860 449952 6866
rect 449900 6802 449952 6808
rect 427679 6502 427685 6554
rect 427737 6502 427749 6554
rect 427801 6502 427813 6554
rect 427865 6502 427877 6554
rect 427929 6502 427941 6554
rect 427993 6502 427999 6554
rect 427679 6381 427999 6502
rect 427679 6325 427691 6381
rect 427747 6325 427771 6381
rect 427827 6325 427851 6381
rect 427907 6325 427931 6381
rect 427987 6325 427999 6381
rect 427679 6301 427999 6325
rect 427679 6245 427691 6301
rect 427747 6245 427771 6301
rect 427827 6245 427851 6301
rect 427907 6245 427931 6301
rect 427987 6245 427999 6301
rect 427679 6221 427999 6245
rect 427679 6165 427691 6221
rect 427747 6165 427771 6221
rect 427827 6165 427851 6221
rect 427907 6165 427931 6221
rect 427987 6165 427999 6221
rect 427679 6141 427999 6165
rect 427679 6085 427691 6141
rect 427747 6085 427771 6141
rect 427827 6085 427851 6141
rect 427907 6085 427931 6141
rect 427987 6085 427999 6141
rect 427679 5466 427999 6085
rect 427679 5414 427685 5466
rect 427737 5414 427749 5466
rect 427801 5414 427813 5466
rect 427865 5414 427877 5466
rect 427929 5414 427941 5466
rect 427993 5414 427999 5466
rect 427679 5022 427999 5414
rect 427679 4966 427691 5022
rect 427747 4966 427771 5022
rect 427827 4966 427851 5022
rect 427907 4966 427931 5022
rect 427987 4966 427999 5022
rect 427679 4942 427999 4966
rect 427679 4886 427691 4942
rect 427747 4886 427771 4942
rect 427827 4886 427851 4942
rect 427907 4886 427931 4942
rect 427987 4886 427999 4942
rect 427679 4862 427999 4886
rect 427679 4806 427691 4862
rect 427747 4806 427771 4862
rect 427827 4806 427851 4862
rect 427907 4806 427931 4862
rect 427987 4806 427999 4862
rect 427679 4782 427999 4806
rect 427679 4726 427691 4782
rect 427747 4726 427771 4782
rect 427827 4726 427851 4782
rect 427907 4726 427931 4782
rect 427987 4726 427999 4782
rect 427679 4378 427999 4726
rect 427679 4326 427685 4378
rect 427737 4326 427749 4378
rect 427801 4326 427813 4378
rect 427865 4326 427877 4378
rect 427929 4326 427941 4378
rect 427993 4326 427999 4378
rect 427679 3663 427999 4326
rect 427679 3607 427691 3663
rect 427747 3607 427771 3663
rect 427827 3607 427851 3663
rect 427907 3607 427931 3663
rect 427987 3607 427999 3663
rect 427679 3583 427999 3607
rect 427679 3527 427691 3583
rect 427747 3527 427771 3583
rect 427827 3527 427851 3583
rect 427907 3527 427931 3583
rect 427987 3527 427999 3583
rect 427679 3503 427999 3527
rect 427679 3447 427691 3503
rect 427747 3447 427771 3503
rect 427827 3447 427851 3503
rect 427907 3447 427931 3503
rect 427987 3447 427999 3503
rect 432972 3528 433024 3534
rect 432972 3470 433024 3476
rect 433432 3528 433484 3534
rect 433432 3470 433484 3476
rect 427679 3423 427999 3447
rect 427679 3367 427691 3423
rect 427747 3367 427771 3423
rect 427827 3367 427851 3423
rect 427907 3367 427931 3423
rect 427987 3367 427999 3423
rect 431684 3460 431736 3466
rect 431684 3402 431736 3408
rect 427679 3290 427999 3367
rect 427679 3238 427685 3290
rect 427737 3238 427749 3290
rect 427801 3238 427813 3290
rect 427865 3238 427877 3290
rect 427929 3238 427941 3290
rect 427993 3238 427999 3290
rect 427679 2202 427999 3238
rect 430764 3052 430816 3058
rect 430764 2994 430816 3000
rect 430776 2854 430804 2994
rect 430764 2848 430816 2854
rect 430764 2790 430816 2796
rect 430776 2417 430804 2790
rect 431696 2446 431724 3402
rect 432984 3058 433012 3470
rect 433340 3392 433392 3398
rect 433340 3334 433392 3340
rect 433352 3194 433380 3334
rect 433340 3188 433392 3194
rect 433340 3130 433392 3136
rect 432972 3052 433024 3058
rect 432972 2994 433024 3000
rect 431868 2984 431920 2990
rect 431868 2926 431920 2932
rect 431880 2553 431908 2926
rect 431866 2544 431922 2553
rect 431866 2479 431922 2488
rect 433352 2446 433380 3130
rect 433444 2446 433472 3470
rect 433524 3460 433576 3466
rect 433524 3402 433576 3408
rect 433536 3058 433564 3402
rect 434536 3392 434588 3398
rect 434536 3334 434588 3340
rect 433524 3052 433576 3058
rect 433524 2994 433576 3000
rect 434548 2446 434576 3334
rect 431684 2440 431736 2446
rect 430762 2408 430818 2417
rect 428188 2372 428240 2378
rect 428188 2314 428240 2320
rect 429752 2372 429804 2378
rect 431684 2382 431736 2388
rect 433340 2440 433392 2446
rect 433340 2382 433392 2388
rect 433432 2440 433484 2446
rect 433432 2382 433484 2388
rect 434536 2440 434588 2446
rect 434536 2382 434588 2388
rect 430762 2343 430818 2352
rect 432880 2372 432932 2378
rect 429752 2314 429804 2320
rect 432880 2314 432932 2320
rect 427679 2150 427685 2202
rect 427737 2150 427749 2202
rect 427801 2150 427813 2202
rect 427865 2150 427877 2202
rect 427929 2150 427941 2202
rect 427993 2150 427999 2202
rect 427679 304 427999 2150
rect 428200 1222 428228 2314
rect 429108 2304 429160 2310
rect 429108 2246 429160 2252
rect 429120 2038 429148 2246
rect 429108 2032 429160 2038
rect 429108 1974 429160 1980
rect 429764 1290 429792 2314
rect 430948 2304 431000 2310
rect 430948 2246 431000 2252
rect 430960 1766 430988 2246
rect 430948 1760 431000 1766
rect 430948 1702 431000 1708
rect 432892 1358 432920 2314
rect 434548 1426 434576 2382
rect 434640 2310 434668 6802
rect 449912 3126 449940 6802
rect 459480 6186 459508 9182
rect 474660 6866 474688 9182
rect 489828 8968 489880 8974
rect 489828 8910 489880 8916
rect 505008 8968 505060 8974
rect 505008 8910 505060 8916
rect 474648 6860 474700 6866
rect 474648 6802 474700 6808
rect 478880 6860 478932 6866
rect 478880 6802 478932 6808
rect 459468 6180 459520 6186
rect 459468 6122 459520 6128
rect 464988 6180 465040 6186
rect 464988 6122 465040 6128
rect 449900 3120 449952 3126
rect 449900 3062 449952 3068
rect 435456 3052 435508 3058
rect 435456 2994 435508 3000
rect 435468 2854 435496 2994
rect 435456 2848 435508 2854
rect 435456 2790 435508 2796
rect 435364 2372 435416 2378
rect 435364 2314 435416 2320
rect 434628 2304 434680 2310
rect 434628 2246 434680 2252
rect 435376 1834 435404 2314
rect 435364 1828 435416 1834
rect 435364 1770 435416 1776
rect 435468 1698 435496 2790
rect 449912 2378 449940 3062
rect 463240 3052 463292 3058
rect 463240 2994 463292 3000
rect 463252 2854 463280 2994
rect 463240 2848 463292 2854
rect 463240 2790 463292 2796
rect 461860 2440 461912 2446
rect 461860 2382 461912 2388
rect 449900 2372 449952 2378
rect 449900 2314 449952 2320
rect 461872 2310 461900 2382
rect 436836 2304 436888 2310
rect 436836 2246 436888 2252
rect 450084 2304 450136 2310
rect 450084 2246 450136 2252
rect 461860 2304 461912 2310
rect 461860 2246 461912 2252
rect 436848 1834 436876 2246
rect 450096 2038 450124 2246
rect 450084 2032 450136 2038
rect 450084 1974 450136 1980
rect 436836 1828 436888 1834
rect 436836 1770 436888 1776
rect 435456 1692 435508 1698
rect 435456 1634 435508 1640
rect 434536 1420 434588 1426
rect 434536 1362 434588 1368
rect 432880 1352 432932 1358
rect 432880 1294 432932 1300
rect 429752 1284 429804 1290
rect 429752 1226 429804 1232
rect 428188 1216 428240 1222
rect 428188 1158 428240 1164
rect 461872 1154 461900 2246
rect 463252 1902 463280 2790
rect 463332 2372 463384 2378
rect 463332 2314 463384 2320
rect 463344 2038 463372 2314
rect 465000 2310 465028 6122
rect 478696 3052 478748 3058
rect 478696 2994 478748 3000
rect 478708 2854 478736 2994
rect 465264 2848 465316 2854
rect 465264 2790 465316 2796
rect 478696 2848 478748 2854
rect 478696 2790 478748 2796
rect 465276 2650 465304 2790
rect 465264 2644 465316 2650
rect 465264 2586 465316 2592
rect 465276 2446 465304 2586
rect 478708 2582 478736 2790
rect 478892 2650 478920 6802
rect 489840 6186 489868 8910
rect 505020 6866 505048 8910
rect 520936 6866 520964 9182
rect 505008 6860 505060 6866
rect 505008 6802 505060 6808
rect 510528 6860 510580 6866
rect 510528 6802 510580 6808
rect 520924 6860 520976 6866
rect 520924 6802 520976 6808
rect 527088 6860 527140 6866
rect 527088 6802 527140 6808
rect 489828 6180 489880 6186
rect 489828 6122 489880 6128
rect 496176 6180 496228 6186
rect 496176 6122 496228 6128
rect 496188 3126 496216 6122
rect 496176 3120 496228 3126
rect 496176 3062 496228 3068
rect 480720 2848 480772 2854
rect 480720 2790 480772 2796
rect 478880 2644 478932 2650
rect 478880 2586 478932 2592
rect 478696 2576 478748 2582
rect 478696 2518 478748 2524
rect 480732 2446 480760 2790
rect 496188 2446 496216 3062
rect 510540 2650 510568 6802
rect 526996 3528 527048 3534
rect 526996 3470 527048 3476
rect 527008 2990 527036 3470
rect 526996 2984 527048 2990
rect 526996 2926 527048 2932
rect 511632 2848 511684 2854
rect 511632 2790 511684 2796
rect 510528 2644 510580 2650
rect 510528 2586 510580 2592
rect 511644 2446 511672 2790
rect 525064 2576 525116 2582
rect 525062 2544 525064 2553
rect 525116 2544 525118 2553
rect 525062 2479 525118 2488
rect 525076 2446 525104 2479
rect 465264 2440 465316 2446
rect 465264 2382 465316 2388
rect 477316 2440 477368 2446
rect 477316 2382 477368 2388
rect 480720 2440 480772 2446
rect 480720 2382 480772 2388
rect 496176 2440 496228 2446
rect 496176 2382 496228 2388
rect 509700 2440 509752 2446
rect 509700 2382 509752 2388
rect 511632 2440 511684 2446
rect 511632 2382 511684 2388
rect 525064 2440 525116 2446
rect 525064 2382 525116 2388
rect 477328 2310 477356 2382
rect 464988 2304 465040 2310
rect 464988 2246 465040 2252
rect 477316 2304 477368 2310
rect 477316 2246 477368 2252
rect 463332 2032 463384 2038
rect 463332 1974 463384 1980
rect 463240 1896 463292 1902
rect 463240 1838 463292 1844
rect 477328 1630 477356 2246
rect 477316 1624 477368 1630
rect 477316 1566 477368 1572
rect 480732 1494 480760 2382
rect 496452 2304 496504 2310
rect 496452 2246 496504 2252
rect 496464 1766 496492 2246
rect 509712 2106 509740 2382
rect 511644 2310 511672 2382
rect 527100 2310 527128 6802
rect 536760 6186 536788 9182
rect 551928 8900 551980 8906
rect 551928 8842 551980 8848
rect 551940 6866 551968 8842
rect 551928 6860 551980 6866
rect 551928 6802 551980 6808
rect 556160 6860 556212 6866
rect 556160 6802 556212 6808
rect 536748 6180 536800 6186
rect 536748 6122 536800 6128
rect 542268 6180 542320 6186
rect 542268 6122 542320 6128
rect 527548 3460 527600 3466
rect 527548 3402 527600 3408
rect 527560 2446 527588 3402
rect 528192 3052 528244 3058
rect 528192 2994 528244 3000
rect 539508 3052 539560 3058
rect 539508 2994 539560 3000
rect 528204 2854 528232 2994
rect 528192 2848 528244 2854
rect 528192 2790 528244 2796
rect 528836 2848 528888 2854
rect 528836 2790 528888 2796
rect 527548 2440 527600 2446
rect 527548 2382 527600 2388
rect 511632 2304 511684 2310
rect 511632 2246 511684 2252
rect 527088 2304 527140 2310
rect 527088 2246 527140 2252
rect 528204 2106 528232 2790
rect 528848 2446 528876 2790
rect 528836 2440 528888 2446
rect 528836 2382 528888 2388
rect 528284 2372 528336 2378
rect 528284 2314 528336 2320
rect 509700 2100 509752 2106
rect 509700 2042 509752 2048
rect 528192 2100 528244 2106
rect 528192 2042 528244 2048
rect 496452 1760 496504 1766
rect 496452 1702 496504 1708
rect 528296 1698 528324 2314
rect 528848 1902 528876 2382
rect 529756 2372 529808 2378
rect 529756 2314 529808 2320
rect 528836 1896 528888 1902
rect 528836 1838 528888 1844
rect 529768 1834 529796 2314
rect 539520 2310 539548 2994
rect 542280 2446 542308 6122
rect 542268 2440 542320 2446
rect 542268 2382 542320 2388
rect 556172 2310 556200 6802
rect 567120 6186 567148 9182
rect 582300 6866 582328 9182
rect 597449 9124 597769 9796
rect 597449 9068 597461 9124
rect 597517 9068 597541 9124
rect 597597 9068 597621 9124
rect 597677 9068 597701 9124
rect 597757 9068 597769 9124
rect 597449 9044 597769 9068
rect 597449 8988 597461 9044
rect 597517 8988 597541 9044
rect 597597 8988 597621 9044
rect 597677 8988 597701 9044
rect 597757 8988 597769 9044
rect 597284 8968 597336 8974
rect 597284 8910 597336 8916
rect 597449 8964 597769 8988
rect 597296 6866 597324 8910
rect 597449 8908 597461 8964
rect 597517 8908 597541 8964
rect 597597 8908 597621 8964
rect 597677 8908 597701 8964
rect 597757 8908 597769 8964
rect 597449 8884 597769 8908
rect 597449 8828 597461 8884
rect 597517 8828 597541 8884
rect 597597 8828 597621 8884
rect 597677 8828 597701 8884
rect 597757 8828 597769 8884
rect 597449 7098 597769 8828
rect 597449 7046 597455 7098
rect 597507 7080 597519 7098
rect 597571 7080 597583 7098
rect 597635 7080 597647 7098
rect 597699 7080 597711 7098
rect 597517 7046 597519 7080
rect 597699 7046 597701 7080
rect 597763 7046 597769 7098
rect 597449 7024 597461 7046
rect 597517 7024 597541 7046
rect 597597 7024 597621 7046
rect 597677 7024 597701 7046
rect 597757 7024 597769 7046
rect 597449 7000 597769 7024
rect 597449 6944 597461 7000
rect 597517 6944 597541 7000
rect 597597 6944 597621 7000
rect 597677 6944 597701 7000
rect 597757 6944 597769 7000
rect 597449 6920 597769 6944
rect 582288 6860 582340 6866
rect 582288 6802 582340 6808
rect 588912 6860 588964 6866
rect 588912 6802 588964 6808
rect 597284 6860 597336 6866
rect 597284 6802 597336 6808
rect 597449 6864 597461 6920
rect 597517 6864 597541 6920
rect 597597 6864 597621 6920
rect 597677 6864 597701 6920
rect 597757 6864 597769 6920
rect 597449 6840 597769 6864
rect 567108 6180 567160 6186
rect 567108 6122 567160 6128
rect 572628 6180 572680 6186
rect 572628 6122 572680 6128
rect 558092 2848 558144 2854
rect 558092 2790 558144 2796
rect 558104 2446 558132 2790
rect 558092 2440 558144 2446
rect 558092 2382 558144 2388
rect 572640 2310 572668 6122
rect 588924 3194 588952 6802
rect 597449 6784 597461 6840
rect 597517 6784 597541 6840
rect 597597 6784 597621 6840
rect 597677 6784 597701 6840
rect 597757 6784 597769 6840
rect 597449 6010 597769 6784
rect 597449 5958 597455 6010
rect 597507 5958 597519 6010
rect 597571 5958 597583 6010
rect 597635 5958 597647 6010
rect 597699 5958 597711 6010
rect 597763 5958 597769 6010
rect 597449 5721 597769 5958
rect 597449 5665 597461 5721
rect 597517 5665 597541 5721
rect 597597 5665 597621 5721
rect 597677 5665 597701 5721
rect 597757 5665 597769 5721
rect 597449 5641 597769 5665
rect 597449 5585 597461 5641
rect 597517 5585 597541 5641
rect 597597 5585 597621 5641
rect 597677 5585 597701 5641
rect 597757 5585 597769 5641
rect 597449 5561 597769 5585
rect 597449 5505 597461 5561
rect 597517 5505 597541 5561
rect 597597 5505 597621 5561
rect 597677 5505 597701 5561
rect 597757 5505 597769 5561
rect 597449 5481 597769 5505
rect 597449 5425 597461 5481
rect 597517 5425 597541 5481
rect 597597 5425 597621 5481
rect 597677 5425 597701 5481
rect 597757 5425 597769 5481
rect 597449 4922 597769 5425
rect 597449 4870 597455 4922
rect 597507 4870 597519 4922
rect 597571 4870 597583 4922
rect 597635 4870 597647 4922
rect 597699 4870 597711 4922
rect 597763 4870 597769 4922
rect 597449 4362 597769 4870
rect 597449 4306 597461 4362
rect 597517 4306 597541 4362
rect 597597 4306 597621 4362
rect 597677 4306 597701 4362
rect 597757 4306 597769 4362
rect 597449 4282 597769 4306
rect 597449 4226 597461 4282
rect 597517 4226 597541 4282
rect 597597 4226 597621 4282
rect 597677 4226 597701 4282
rect 597757 4226 597769 4282
rect 597449 4202 597769 4226
rect 597449 4146 597461 4202
rect 597517 4146 597541 4202
rect 597597 4146 597621 4202
rect 597677 4146 597701 4202
rect 597757 4146 597769 4202
rect 597449 4122 597769 4146
rect 597449 4066 597461 4122
rect 597517 4066 597541 4122
rect 597597 4066 597621 4122
rect 597677 4066 597701 4122
rect 597757 4066 597769 4122
rect 597449 3834 597769 4066
rect 597449 3782 597455 3834
rect 597507 3782 597519 3834
rect 597571 3782 597583 3834
rect 597635 3782 597647 3834
rect 597699 3782 597711 3834
rect 597763 3782 597769 3834
rect 588912 3188 588964 3194
rect 588912 3130 588964 3136
rect 573916 2984 573968 2990
rect 573916 2926 573968 2932
rect 573928 2446 573956 2926
rect 588924 2446 588952 3130
rect 597449 3003 597769 3782
rect 597449 2947 597461 3003
rect 597517 2947 597541 3003
rect 597597 2947 597621 3003
rect 597677 2947 597701 3003
rect 597757 2947 597769 3003
rect 597449 2923 597769 2947
rect 597449 2867 597461 2923
rect 597517 2867 597541 2923
rect 597597 2867 597621 2923
rect 597677 2867 597701 2923
rect 597757 2867 597769 2923
rect 597449 2843 597769 2867
rect 597449 2787 597461 2843
rect 597517 2787 597541 2843
rect 597597 2787 597621 2843
rect 597677 2787 597701 2843
rect 597757 2787 597769 2843
rect 597449 2763 597769 2787
rect 597449 2746 597461 2763
rect 597517 2746 597541 2763
rect 597597 2746 597621 2763
rect 597677 2746 597701 2763
rect 597757 2746 597769 2763
rect 597449 2694 597455 2746
rect 597517 2707 597519 2746
rect 597699 2707 597701 2746
rect 597507 2694 597519 2707
rect 597571 2694 597583 2707
rect 597635 2694 597647 2707
rect 597699 2694 597711 2707
rect 597763 2694 597769 2746
rect 573916 2440 573968 2446
rect 573916 2382 573968 2388
rect 588912 2440 588964 2446
rect 588912 2382 588964 2388
rect 530952 2304 531004 2310
rect 530952 2246 531004 2252
rect 539508 2304 539560 2310
rect 539508 2246 539560 2252
rect 555332 2304 555384 2310
rect 555332 2246 555384 2252
rect 556160 2304 556212 2310
rect 556160 2246 556212 2252
rect 572628 2304 572680 2310
rect 572628 2246 572680 2252
rect 589188 2304 589240 2310
rect 589188 2246 589240 2252
rect 530964 1970 530992 2246
rect 555344 2038 555372 2246
rect 589200 2106 589228 2246
rect 589188 2100 589240 2106
rect 589188 2042 589240 2048
rect 555332 2032 555384 2038
rect 555332 1974 555384 1980
rect 530952 1964 531004 1970
rect 530952 1906 531004 1912
rect 529756 1828 529808 1834
rect 529756 1770 529808 1776
rect 528284 1692 528336 1698
rect 528284 1634 528336 1640
rect 480720 1488 480772 1494
rect 480720 1430 480772 1436
rect 461860 1148 461912 1154
rect 461860 1090 461912 1096
rect 427679 248 427691 304
rect 427747 248 427771 304
rect 427827 248 427851 304
rect 427907 248 427931 304
rect 427987 248 427999 304
rect 427679 224 427999 248
rect 427679 168 427691 224
rect 427747 168 427771 224
rect 427827 168 427851 224
rect 427907 168 427931 224
rect 427987 168 427999 224
rect 427679 144 427999 168
rect 427679 88 427691 144
rect 427747 88 427771 144
rect 427827 88 427851 144
rect 427907 88 427931 144
rect 427987 88 427999 144
rect 427679 64 427999 88
rect 427679 8 427691 64
rect 427747 8 427771 64
rect 427827 8 427851 64
rect 427907 8 427931 64
rect 427987 8 427999 64
rect 427679 -4 427999 8
rect 597449 964 597769 2694
rect 597449 908 597461 964
rect 597517 908 597541 964
rect 597597 908 597621 964
rect 597677 908 597701 964
rect 597757 908 597769 964
rect 597449 884 597769 908
rect 597449 828 597461 884
rect 597517 828 597541 884
rect 597597 828 597621 884
rect 597677 828 597701 884
rect 597757 828 597769 884
rect 597449 804 597769 828
rect 597449 748 597461 804
rect 597517 748 597541 804
rect 597597 748 597621 804
rect 597677 748 597701 804
rect 597757 748 597769 804
rect 597449 724 597769 748
rect 597449 668 597461 724
rect 597517 668 597541 724
rect 597597 668 597621 724
rect 597677 668 597701 724
rect 597757 668 597769 724
rect 597449 -4 597769 668
rect 598109 9784 598429 9796
rect 598109 9728 598121 9784
rect 598177 9728 598201 9784
rect 598257 9728 598281 9784
rect 598337 9728 598361 9784
rect 598417 9728 598429 9784
rect 598109 9704 598429 9728
rect 598109 9648 598121 9704
rect 598177 9648 598201 9704
rect 598257 9648 598281 9704
rect 598337 9648 598361 9704
rect 598417 9648 598429 9704
rect 598109 9624 598429 9648
rect 598109 9568 598121 9624
rect 598177 9568 598201 9624
rect 598257 9568 598281 9624
rect 598337 9568 598361 9624
rect 598417 9568 598429 9624
rect 598109 9544 598429 9568
rect 598109 9488 598121 9544
rect 598177 9488 598201 9544
rect 598257 9488 598281 9544
rect 598337 9488 598361 9544
rect 598417 9488 598429 9544
rect 598109 7740 598429 9488
rect 684684 9784 685004 9796
rect 684684 9728 684696 9784
rect 684752 9728 684776 9784
rect 684832 9728 684856 9784
rect 684912 9728 684936 9784
rect 684992 9728 685004 9784
rect 684684 9704 685004 9728
rect 684684 9648 684696 9704
rect 684752 9648 684776 9704
rect 684832 9648 684856 9704
rect 684912 9648 684936 9704
rect 684992 9648 685004 9704
rect 684684 9624 685004 9648
rect 684684 9568 684696 9624
rect 684752 9568 684776 9624
rect 684832 9568 684856 9624
rect 684912 9568 684936 9624
rect 684992 9568 685004 9624
rect 684684 9544 685004 9568
rect 684684 9488 684696 9544
rect 684752 9488 684776 9544
rect 684832 9488 684856 9544
rect 684912 9488 684936 9544
rect 684992 9488 685004 9544
rect 612648 9240 612700 9246
rect 612648 9182 612700 9188
rect 627644 9240 627696 9246
rect 627644 9182 627696 9188
rect 673368 9240 673420 9246
rect 673368 9182 673420 9188
rect 598109 7684 598121 7740
rect 598177 7684 598201 7740
rect 598257 7684 598281 7740
rect 598337 7684 598361 7740
rect 598417 7684 598429 7740
rect 598109 7660 598429 7684
rect 598109 7642 598121 7660
rect 598177 7642 598201 7660
rect 598257 7642 598281 7660
rect 598337 7642 598361 7660
rect 598417 7642 598429 7660
rect 598109 7590 598115 7642
rect 598177 7604 598179 7642
rect 598359 7604 598361 7642
rect 598167 7590 598179 7604
rect 598231 7590 598243 7604
rect 598295 7590 598307 7604
rect 598359 7590 598371 7604
rect 598423 7590 598429 7642
rect 598109 7580 598429 7590
rect 598109 7524 598121 7580
rect 598177 7524 598201 7580
rect 598257 7524 598281 7580
rect 598337 7524 598361 7580
rect 598417 7524 598429 7580
rect 598109 7500 598429 7524
rect 598109 7444 598121 7500
rect 598177 7444 598201 7500
rect 598257 7444 598281 7500
rect 598337 7444 598361 7500
rect 598417 7444 598429 7500
rect 598109 6554 598429 7444
rect 604644 6860 604696 6866
rect 604644 6802 604696 6808
rect 598109 6502 598115 6554
rect 598167 6502 598179 6554
rect 598231 6502 598243 6554
rect 598295 6502 598307 6554
rect 598359 6502 598371 6554
rect 598423 6502 598429 6554
rect 598109 6381 598429 6502
rect 598109 6325 598121 6381
rect 598177 6325 598201 6381
rect 598257 6325 598281 6381
rect 598337 6325 598361 6381
rect 598417 6325 598429 6381
rect 598109 6301 598429 6325
rect 598109 6245 598121 6301
rect 598177 6245 598201 6301
rect 598257 6245 598281 6301
rect 598337 6245 598361 6301
rect 598417 6245 598429 6301
rect 598109 6221 598429 6245
rect 598109 6165 598121 6221
rect 598177 6165 598201 6221
rect 598257 6165 598281 6221
rect 598337 6165 598361 6221
rect 598417 6165 598429 6221
rect 598109 6141 598429 6165
rect 598109 6085 598121 6141
rect 598177 6085 598201 6141
rect 598257 6085 598281 6141
rect 598337 6085 598361 6141
rect 598417 6085 598429 6141
rect 598109 5466 598429 6085
rect 598109 5414 598115 5466
rect 598167 5414 598179 5466
rect 598231 5414 598243 5466
rect 598295 5414 598307 5466
rect 598359 5414 598371 5466
rect 598423 5414 598429 5466
rect 598109 5022 598429 5414
rect 598109 4966 598121 5022
rect 598177 4966 598201 5022
rect 598257 4966 598281 5022
rect 598337 4966 598361 5022
rect 598417 4966 598429 5022
rect 598109 4942 598429 4966
rect 598109 4886 598121 4942
rect 598177 4886 598201 4942
rect 598257 4886 598281 4942
rect 598337 4886 598361 4942
rect 598417 4886 598429 4942
rect 598109 4862 598429 4886
rect 598109 4806 598121 4862
rect 598177 4806 598201 4862
rect 598257 4806 598281 4862
rect 598337 4806 598361 4862
rect 598417 4806 598429 4862
rect 598109 4782 598429 4806
rect 598109 4726 598121 4782
rect 598177 4726 598201 4782
rect 598257 4726 598281 4782
rect 598337 4726 598361 4782
rect 598417 4726 598429 4782
rect 598109 4378 598429 4726
rect 598109 4326 598115 4378
rect 598167 4326 598179 4378
rect 598231 4326 598243 4378
rect 598295 4326 598307 4378
rect 598359 4326 598371 4378
rect 598423 4326 598429 4378
rect 598109 3663 598429 4326
rect 598109 3607 598121 3663
rect 598177 3607 598201 3663
rect 598257 3607 598281 3663
rect 598337 3607 598361 3663
rect 598417 3607 598429 3663
rect 598109 3583 598429 3607
rect 598109 3527 598121 3583
rect 598177 3527 598201 3583
rect 598257 3527 598281 3583
rect 598337 3527 598361 3583
rect 598417 3527 598429 3583
rect 598109 3503 598429 3527
rect 598109 3447 598121 3503
rect 598177 3447 598201 3503
rect 598257 3447 598281 3503
rect 598337 3447 598361 3503
rect 598417 3447 598429 3503
rect 598109 3423 598429 3447
rect 598109 3367 598121 3423
rect 598177 3367 598201 3423
rect 598257 3367 598281 3423
rect 598337 3367 598361 3423
rect 598417 3367 598429 3423
rect 598109 3290 598429 3367
rect 598109 3238 598115 3290
rect 598167 3238 598179 3290
rect 598231 3238 598243 3290
rect 598295 3238 598307 3290
rect 598359 3238 598371 3290
rect 598423 3238 598429 3290
rect 598109 2202 598429 3238
rect 604460 2848 604512 2854
rect 604460 2790 604512 2796
rect 604472 2650 604500 2790
rect 604656 2650 604684 6802
rect 612660 6186 612688 9182
rect 627656 6186 627684 9182
rect 643008 8968 643060 8974
rect 643008 8910 643060 8916
rect 658188 8968 658240 8974
rect 658188 8910 658240 8916
rect 643020 6186 643048 8910
rect 658200 6866 658228 8910
rect 658188 6860 658240 6866
rect 658188 6802 658240 6808
rect 666468 6860 666520 6866
rect 666468 6802 666520 6808
rect 612648 6180 612700 6186
rect 612648 6122 612700 6128
rect 620100 6180 620152 6186
rect 620100 6122 620152 6128
rect 627644 6180 627696 6186
rect 627644 6122 627696 6128
rect 635556 6180 635608 6186
rect 635556 6122 635608 6128
rect 643008 6180 643060 6186
rect 643008 6122 643060 6128
rect 651012 6180 651064 6186
rect 651012 6122 651064 6128
rect 619824 2848 619876 2854
rect 619824 2790 619876 2796
rect 604460 2644 604512 2650
rect 604460 2586 604512 2592
rect 604644 2644 604696 2650
rect 604644 2586 604696 2592
rect 604472 2446 604500 2586
rect 619836 2582 619864 2790
rect 620112 2650 620140 6122
rect 620100 2644 620152 2650
rect 620100 2586 620152 2592
rect 625436 2644 625488 2650
rect 625436 2586 625488 2592
rect 619824 2576 619876 2582
rect 619824 2518 619876 2524
rect 619836 2446 619864 2518
rect 625448 2446 625476 2586
rect 635568 2446 635596 6122
rect 650736 2848 650788 2854
rect 650736 2790 650788 2796
rect 604460 2440 604512 2446
rect 604460 2382 604512 2388
rect 619824 2440 619876 2446
rect 619824 2382 619876 2388
rect 625436 2440 625488 2446
rect 625436 2382 625488 2388
rect 635556 2440 635608 2446
rect 635556 2382 635608 2388
rect 650748 2378 650776 2790
rect 651024 2582 651052 6122
rect 666192 2848 666244 2854
rect 666192 2790 666244 2796
rect 651012 2576 651064 2582
rect 651012 2518 651064 2524
rect 666204 2514 666232 2790
rect 666480 2582 666508 6802
rect 673380 6186 673408 9182
rect 684024 9124 684344 9136
rect 684024 9068 684036 9124
rect 684092 9068 684116 9124
rect 684172 9068 684196 9124
rect 684252 9068 684276 9124
rect 684332 9068 684344 9124
rect 684024 9044 684344 9068
rect 684024 8988 684036 9044
rect 684092 8988 684116 9044
rect 684172 8988 684196 9044
rect 684252 8988 684276 9044
rect 684332 8988 684344 9044
rect 684024 8964 684344 8988
rect 684024 8908 684036 8964
rect 684092 8908 684116 8964
rect 684172 8908 684196 8964
rect 684252 8908 684276 8964
rect 684332 8908 684344 8964
rect 684024 8884 684344 8908
rect 684024 8828 684036 8884
rect 684092 8828 684116 8884
rect 684172 8828 684196 8884
rect 684252 8828 684276 8884
rect 684332 8828 684344 8884
rect 684024 7080 684344 8828
rect 684024 7024 684036 7080
rect 684092 7024 684116 7080
rect 684172 7024 684196 7080
rect 684252 7024 684276 7080
rect 684332 7024 684344 7080
rect 684024 7000 684344 7024
rect 684024 6944 684036 7000
rect 684092 6944 684116 7000
rect 684172 6944 684196 7000
rect 684252 6944 684276 7000
rect 684332 6944 684344 7000
rect 684024 6920 684344 6944
rect 684024 6864 684036 6920
rect 684092 6864 684116 6920
rect 684172 6864 684196 6920
rect 684252 6864 684276 6920
rect 684332 6864 684344 6920
rect 684024 6840 684344 6864
rect 684024 6784 684036 6840
rect 684092 6784 684116 6840
rect 684172 6784 684196 6840
rect 684252 6784 684276 6840
rect 684332 6784 684344 6840
rect 673368 6180 673420 6186
rect 673368 6122 673420 6128
rect 681740 6180 681792 6186
rect 681740 6122 681792 6128
rect 681752 3194 681780 6122
rect 684024 5721 684344 6784
rect 684024 5665 684036 5721
rect 684092 5665 684116 5721
rect 684172 5665 684196 5721
rect 684252 5665 684276 5721
rect 684332 5665 684344 5721
rect 684024 5641 684344 5665
rect 684024 5585 684036 5641
rect 684092 5585 684116 5641
rect 684172 5585 684196 5641
rect 684252 5585 684276 5641
rect 684332 5585 684344 5641
rect 684024 5561 684344 5585
rect 684024 5505 684036 5561
rect 684092 5505 684116 5561
rect 684172 5505 684196 5561
rect 684252 5505 684276 5561
rect 684332 5505 684344 5561
rect 684024 5481 684344 5505
rect 684024 5425 684036 5481
rect 684092 5425 684116 5481
rect 684172 5425 684196 5481
rect 684252 5425 684276 5481
rect 684332 5425 684344 5481
rect 684024 4362 684344 5425
rect 684024 4306 684036 4362
rect 684092 4306 684116 4362
rect 684172 4306 684196 4362
rect 684252 4306 684276 4362
rect 684332 4306 684344 4362
rect 684024 4282 684344 4306
rect 684024 4226 684036 4282
rect 684092 4226 684116 4282
rect 684172 4226 684196 4282
rect 684252 4226 684276 4282
rect 684332 4226 684344 4282
rect 684024 4202 684344 4226
rect 684024 4146 684036 4202
rect 684092 4146 684116 4202
rect 684172 4146 684196 4202
rect 684252 4146 684276 4202
rect 684332 4146 684344 4202
rect 684024 4122 684344 4146
rect 684024 4066 684036 4122
rect 684092 4066 684116 4122
rect 684172 4066 684196 4122
rect 684252 4066 684276 4122
rect 684332 4066 684344 4122
rect 681740 3188 681792 3194
rect 681740 3130 681792 3136
rect 666468 2576 666520 2582
rect 666468 2518 666520 2524
rect 666192 2508 666244 2514
rect 666192 2450 666244 2456
rect 681752 2446 681780 3130
rect 684024 3003 684344 4066
rect 684024 2947 684036 3003
rect 684092 2947 684116 3003
rect 684172 2947 684196 3003
rect 684252 2947 684276 3003
rect 684332 2947 684344 3003
rect 684024 2923 684344 2947
rect 684024 2867 684036 2923
rect 684092 2867 684116 2923
rect 684172 2867 684196 2923
rect 684252 2867 684276 2923
rect 684332 2867 684344 2923
rect 684024 2843 684344 2867
rect 684024 2787 684036 2843
rect 684092 2787 684116 2843
rect 684172 2787 684196 2843
rect 684252 2787 684276 2843
rect 684332 2787 684344 2843
rect 684024 2763 684344 2787
rect 684024 2707 684036 2763
rect 684092 2707 684116 2763
rect 684172 2707 684196 2763
rect 684252 2707 684276 2763
rect 684332 2707 684344 2763
rect 681740 2440 681792 2446
rect 681740 2382 681792 2388
rect 623044 2372 623096 2378
rect 623044 2314 623096 2320
rect 624884 2372 624936 2378
rect 624884 2314 624936 2320
rect 650736 2372 650788 2378
rect 650736 2314 650788 2320
rect 598109 2150 598115 2202
rect 598167 2150 598179 2202
rect 598231 2150 598243 2202
rect 598295 2150 598307 2202
rect 598359 2150 598371 2202
rect 598423 2150 598429 2202
rect 598109 304 598429 2150
rect 623056 1902 623084 2314
rect 624896 1970 624924 2314
rect 624884 1964 624936 1970
rect 624884 1906 624936 1912
rect 623044 1896 623096 1902
rect 623044 1838 623096 1844
rect 684024 964 684344 2707
rect 684024 908 684036 964
rect 684092 908 684116 964
rect 684172 908 684196 964
rect 684252 908 684276 964
rect 684332 908 684344 964
rect 684024 884 684344 908
rect 684024 828 684036 884
rect 684092 828 684116 884
rect 684172 828 684196 884
rect 684252 828 684276 884
rect 684332 828 684344 884
rect 684024 804 684344 828
rect 684024 748 684036 804
rect 684092 748 684116 804
rect 684172 748 684196 804
rect 684252 748 684276 804
rect 684332 748 684344 804
rect 684024 724 684344 748
rect 684024 668 684036 724
rect 684092 668 684116 724
rect 684172 668 684196 724
rect 684252 668 684276 724
rect 684332 668 684344 724
rect 684024 656 684344 668
rect 684684 7740 685004 9488
rect 684684 7684 684696 7740
rect 684752 7684 684776 7740
rect 684832 7684 684856 7740
rect 684912 7684 684936 7740
rect 684992 7684 685004 7740
rect 684684 7660 685004 7684
rect 684684 7604 684696 7660
rect 684752 7604 684776 7660
rect 684832 7604 684856 7660
rect 684912 7604 684936 7660
rect 684992 7604 685004 7660
rect 684684 7580 685004 7604
rect 684684 7524 684696 7580
rect 684752 7524 684776 7580
rect 684832 7524 684856 7580
rect 684912 7524 684936 7580
rect 684992 7524 685004 7580
rect 684684 7500 685004 7524
rect 684684 7444 684696 7500
rect 684752 7444 684776 7500
rect 684832 7444 684856 7500
rect 684912 7444 684936 7500
rect 684992 7444 685004 7500
rect 684684 6381 685004 7444
rect 684684 6325 684696 6381
rect 684752 6325 684776 6381
rect 684832 6325 684856 6381
rect 684912 6325 684936 6381
rect 684992 6325 685004 6381
rect 684684 6301 685004 6325
rect 684684 6245 684696 6301
rect 684752 6245 684776 6301
rect 684832 6245 684856 6301
rect 684912 6245 684936 6301
rect 684992 6245 685004 6301
rect 684684 6221 685004 6245
rect 684684 6165 684696 6221
rect 684752 6165 684776 6221
rect 684832 6165 684856 6221
rect 684912 6165 684936 6221
rect 684992 6165 685004 6221
rect 684684 6141 685004 6165
rect 684684 6085 684696 6141
rect 684752 6085 684776 6141
rect 684832 6085 684856 6141
rect 684912 6085 684936 6141
rect 684992 6085 685004 6141
rect 684684 5022 685004 6085
rect 684684 4966 684696 5022
rect 684752 4966 684776 5022
rect 684832 4966 684856 5022
rect 684912 4966 684936 5022
rect 684992 4966 685004 5022
rect 684684 4942 685004 4966
rect 684684 4886 684696 4942
rect 684752 4886 684776 4942
rect 684832 4886 684856 4942
rect 684912 4886 684936 4942
rect 684992 4886 685004 4942
rect 684684 4862 685004 4886
rect 684684 4806 684696 4862
rect 684752 4806 684776 4862
rect 684832 4806 684856 4862
rect 684912 4806 684936 4862
rect 684992 4806 685004 4862
rect 684684 4782 685004 4806
rect 684684 4726 684696 4782
rect 684752 4726 684776 4782
rect 684832 4726 684856 4782
rect 684912 4726 684936 4782
rect 684992 4726 685004 4782
rect 684684 3663 685004 4726
rect 684684 3607 684696 3663
rect 684752 3607 684776 3663
rect 684832 3607 684856 3663
rect 684912 3607 684936 3663
rect 684992 3607 685004 3663
rect 684684 3583 685004 3607
rect 684684 3527 684696 3583
rect 684752 3527 684776 3583
rect 684832 3527 684856 3583
rect 684912 3527 684936 3583
rect 684992 3527 685004 3583
rect 684684 3503 685004 3527
rect 684684 3447 684696 3503
rect 684752 3447 684776 3503
rect 684832 3447 684856 3503
rect 684912 3447 684936 3503
rect 684992 3447 685004 3503
rect 684684 3423 685004 3447
rect 684684 3367 684696 3423
rect 684752 3367 684776 3423
rect 684832 3367 684856 3423
rect 684912 3367 684936 3423
rect 684992 3367 685004 3423
rect 598109 248 598121 304
rect 598177 248 598201 304
rect 598257 248 598281 304
rect 598337 248 598361 304
rect 598417 248 598429 304
rect 598109 224 598429 248
rect 598109 168 598121 224
rect 598177 168 598201 224
rect 598257 168 598281 224
rect 598337 168 598361 224
rect 598417 168 598429 224
rect 598109 144 598429 168
rect 598109 88 598121 144
rect 598177 88 598201 144
rect 598257 88 598281 144
rect 598337 88 598361 144
rect 598417 88 598429 144
rect 598109 64 598429 88
rect 598109 8 598121 64
rect 598177 8 598201 64
rect 598257 8 598281 64
rect 598337 8 598361 64
rect 598417 8 598429 64
rect 598109 -4 598429 8
rect 684684 304 685004 3367
rect 684684 248 684696 304
rect 684752 248 684776 304
rect 684832 248 684856 304
rect 684912 248 684936 304
rect 684992 248 685004 304
rect 684684 224 685004 248
rect 684684 168 684696 224
rect 684752 168 684776 224
rect 684832 168 684856 224
rect 684912 168 684936 224
rect 684992 168 685004 224
rect 684684 144 685004 168
rect 684684 88 684696 144
rect 684752 88 684776 144
rect 684832 88 684856 144
rect 684912 88 684936 144
rect 684992 88 685004 144
rect 684684 64 685004 88
rect 684684 8 684696 64
rect 684752 8 684776 64
rect 684832 8 684856 64
rect 684912 8 684936 64
rect 684992 8 685004 64
rect 684684 -4 685004 8
<< via2 >>
rect -1064 9728 -1008 9784
rect -984 9728 -928 9784
rect -904 9728 -848 9784
rect -824 9728 -768 9784
rect -1064 9648 -1008 9704
rect -984 9648 -928 9704
rect -904 9648 -848 9704
rect -824 9648 -768 9704
rect -1064 9568 -1008 9624
rect -984 9568 -928 9624
rect -904 9568 -848 9624
rect -824 9568 -768 9624
rect -1064 9488 -1008 9544
rect -984 9488 -928 9544
rect -904 9488 -848 9544
rect -824 9488 -768 9544
rect -1064 7684 -1008 7740
rect -984 7684 -928 7740
rect -904 7684 -848 7740
rect -824 7684 -768 7740
rect -1064 7604 -1008 7660
rect -984 7604 -928 7660
rect -904 7604 -848 7660
rect -824 7604 -768 7660
rect -1064 7524 -1008 7580
rect -984 7524 -928 7580
rect -904 7524 -848 7580
rect -824 7524 -768 7580
rect -1064 7444 -1008 7500
rect -984 7444 -928 7500
rect -904 7444 -848 7500
rect -824 7444 -768 7500
rect -1064 6325 -1008 6381
rect -984 6325 -928 6381
rect -904 6325 -848 6381
rect -824 6325 -768 6381
rect -1064 6245 -1008 6301
rect -984 6245 -928 6301
rect -904 6245 -848 6301
rect -824 6245 -768 6301
rect -1064 6165 -1008 6221
rect -984 6165 -928 6221
rect -904 6165 -848 6221
rect -824 6165 -768 6221
rect -1064 6085 -1008 6141
rect -984 6085 -928 6141
rect -904 6085 -848 6141
rect -824 6085 -768 6141
rect -1064 4966 -1008 5022
rect -984 4966 -928 5022
rect -904 4966 -848 5022
rect -824 4966 -768 5022
rect -1064 4886 -1008 4942
rect -984 4886 -928 4942
rect -904 4886 -848 4942
rect -824 4886 -768 4942
rect -1064 4806 -1008 4862
rect -984 4806 -928 4862
rect -904 4806 -848 4862
rect -824 4806 -768 4862
rect -1064 4726 -1008 4782
rect -984 4726 -928 4782
rect -904 4726 -848 4782
rect -824 4726 -768 4782
rect -1064 3607 -1008 3663
rect -984 3607 -928 3663
rect -904 3607 -848 3663
rect -824 3607 -768 3663
rect -1064 3527 -1008 3583
rect -984 3527 -928 3583
rect -904 3527 -848 3583
rect -824 3527 -768 3583
rect -1064 3447 -1008 3503
rect -984 3447 -928 3503
rect -904 3447 -848 3503
rect -824 3447 -768 3503
rect -1064 3367 -1008 3423
rect -984 3367 -928 3423
rect -904 3367 -848 3423
rect -824 3367 -768 3423
rect -404 9068 -348 9124
rect -324 9068 -268 9124
rect -244 9068 -188 9124
rect -164 9068 -108 9124
rect -404 8988 -348 9044
rect -324 8988 -268 9044
rect -244 8988 -188 9044
rect -164 8988 -108 9044
rect -404 8908 -348 8964
rect -324 8908 -268 8964
rect -244 8908 -188 8964
rect -164 8908 -108 8964
rect -404 8828 -348 8884
rect -324 8828 -268 8884
rect -244 8828 -188 8884
rect -164 8828 -108 8884
rect -404 7024 -348 7080
rect -324 7024 -268 7080
rect -244 7024 -188 7080
rect -164 7024 -108 7080
rect -404 6944 -348 7000
rect -324 6944 -268 7000
rect -244 6944 -188 7000
rect -164 6944 -108 7000
rect -404 6864 -348 6920
rect -324 6864 -268 6920
rect -244 6864 -188 6920
rect -164 6864 -108 6920
rect -404 6784 -348 6840
rect -324 6784 -268 6840
rect -244 6784 -188 6840
rect -164 6784 -108 6840
rect -404 5665 -348 5721
rect -324 5665 -268 5721
rect -244 5665 -188 5721
rect -164 5665 -108 5721
rect -404 5585 -348 5641
rect -324 5585 -268 5641
rect -244 5585 -188 5641
rect -164 5585 -108 5641
rect -404 5505 -348 5561
rect -324 5505 -268 5561
rect -244 5505 -188 5561
rect -164 5505 -108 5561
rect -404 5425 -348 5481
rect -324 5425 -268 5481
rect -244 5425 -188 5481
rect -164 5425 -108 5481
rect -404 4306 -348 4362
rect -324 4306 -268 4362
rect -244 4306 -188 4362
rect -164 4306 -108 4362
rect -404 4226 -348 4282
rect -324 4226 -268 4282
rect -244 4226 -188 4282
rect -164 4226 -108 4282
rect -404 4146 -348 4202
rect -324 4146 -268 4202
rect -244 4146 -188 4202
rect -164 4146 -108 4202
rect -404 4066 -348 4122
rect -324 4066 -268 4122
rect -244 4066 -188 4122
rect -164 4066 -108 4122
rect -404 2947 -348 3003
rect -324 2947 -268 3003
rect -244 2947 -188 3003
rect -164 2947 -108 3003
rect -404 2867 -348 2923
rect -324 2867 -268 2923
rect -244 2867 -188 2923
rect -164 2867 -108 2923
rect -404 2787 -348 2843
rect -324 2787 -268 2843
rect -244 2787 -188 2843
rect -164 2787 -108 2843
rect -404 2707 -348 2763
rect -324 2707 -268 2763
rect -244 2707 -188 2763
rect -164 2707 -108 2763
rect 86171 9068 86227 9124
rect 86251 9068 86307 9124
rect 86331 9068 86387 9124
rect 86411 9068 86467 9124
rect 86171 8988 86227 9044
rect 86251 8988 86307 9044
rect 86331 8988 86387 9044
rect 86411 8988 86467 9044
rect 86171 8908 86227 8964
rect 86251 8908 86307 8964
rect 86331 8908 86387 8964
rect 86411 8908 86467 8964
rect 86171 8828 86227 8884
rect 86251 8828 86307 8884
rect 86331 8828 86387 8884
rect 86411 8828 86467 8884
rect 86171 7046 86217 7080
rect 86217 7046 86227 7080
rect 86251 7046 86281 7080
rect 86281 7046 86293 7080
rect 86293 7046 86307 7080
rect 86331 7046 86345 7080
rect 86345 7046 86357 7080
rect 86357 7046 86387 7080
rect 86411 7046 86421 7080
rect 86421 7046 86467 7080
rect 86171 7024 86227 7046
rect 86251 7024 86307 7046
rect 86331 7024 86387 7046
rect 86411 7024 86467 7046
rect 86171 6944 86227 7000
rect 86251 6944 86307 7000
rect 86331 6944 86387 7000
rect 86411 6944 86467 7000
rect 86171 6864 86227 6920
rect 86251 6864 86307 6920
rect 86331 6864 86387 6920
rect 86411 6864 86467 6920
rect 86171 6784 86227 6840
rect 86251 6784 86307 6840
rect 86331 6784 86387 6840
rect 86411 6784 86467 6840
rect 86171 5665 86227 5721
rect 86251 5665 86307 5721
rect 86331 5665 86387 5721
rect 86411 5665 86467 5721
rect 86171 5585 86227 5641
rect 86251 5585 86307 5641
rect 86331 5585 86387 5641
rect 86411 5585 86467 5641
rect 86171 5505 86227 5561
rect 86251 5505 86307 5561
rect 86331 5505 86387 5561
rect 86411 5505 86467 5561
rect 86171 5425 86227 5481
rect 86251 5425 86307 5481
rect 86331 5425 86387 5481
rect 86411 5425 86467 5481
rect 86171 4306 86227 4362
rect 86251 4306 86307 4362
rect 86331 4306 86387 4362
rect 86411 4306 86467 4362
rect 86171 4226 86227 4282
rect 86251 4226 86307 4282
rect 86331 4226 86387 4282
rect 86411 4226 86467 4282
rect 86171 4146 86227 4202
rect 86251 4146 86307 4202
rect 86331 4146 86387 4202
rect 86411 4146 86467 4202
rect 86171 4066 86227 4122
rect 86251 4066 86307 4122
rect 86331 4066 86387 4122
rect 86411 4066 86467 4122
rect 86171 2947 86227 3003
rect 86251 2947 86307 3003
rect 86331 2947 86387 3003
rect 86411 2947 86467 3003
rect 86171 2867 86227 2923
rect 86251 2867 86307 2923
rect 86331 2867 86387 2923
rect 86411 2867 86467 2923
rect 86171 2787 86227 2843
rect 86251 2787 86307 2843
rect 86331 2787 86387 2843
rect 86411 2787 86467 2843
rect 86171 2746 86227 2763
rect 86251 2746 86307 2763
rect 86331 2746 86387 2763
rect 86411 2746 86467 2763
rect 86171 2707 86217 2746
rect 86217 2707 86227 2746
rect 86251 2707 86281 2746
rect 86281 2707 86293 2746
rect 86293 2707 86307 2746
rect 86331 2707 86345 2746
rect 86345 2707 86357 2746
rect 86357 2707 86387 2746
rect 86411 2707 86421 2746
rect 86421 2707 86467 2746
rect -404 908 -348 964
rect -324 908 -268 964
rect -244 908 -188 964
rect -164 908 -108 964
rect -404 828 -348 884
rect -324 828 -268 884
rect -244 828 -188 884
rect -164 828 -108 884
rect -404 748 -348 804
rect -324 748 -268 804
rect -244 748 -188 804
rect -164 748 -108 804
rect -404 668 -348 724
rect -324 668 -268 724
rect -244 668 -188 724
rect -164 668 -108 724
rect 86171 908 86227 964
rect 86251 908 86307 964
rect 86331 908 86387 964
rect 86411 908 86467 964
rect 86171 828 86227 884
rect 86251 828 86307 884
rect 86331 828 86387 884
rect 86411 828 86467 884
rect 86171 748 86227 804
rect 86251 748 86307 804
rect 86331 748 86387 804
rect 86411 748 86467 804
rect 86171 668 86227 724
rect 86251 668 86307 724
rect 86331 668 86387 724
rect 86411 668 86467 724
rect -1064 248 -1008 304
rect -984 248 -928 304
rect -904 248 -848 304
rect -824 248 -768 304
rect -1064 168 -1008 224
rect -984 168 -928 224
rect -904 168 -848 224
rect -824 168 -768 224
rect -1064 88 -1008 144
rect -984 88 -928 144
rect -904 88 -848 144
rect -824 88 -768 144
rect -1064 8 -1008 64
rect -984 8 -928 64
rect -904 8 -848 64
rect -824 8 -768 64
rect 86831 9728 86887 9784
rect 86911 9728 86967 9784
rect 86991 9728 87047 9784
rect 87071 9728 87127 9784
rect 86831 9648 86887 9704
rect 86911 9648 86967 9704
rect 86991 9648 87047 9704
rect 87071 9648 87127 9704
rect 86831 9568 86887 9624
rect 86911 9568 86967 9624
rect 86991 9568 87047 9624
rect 87071 9568 87127 9624
rect 86831 9488 86887 9544
rect 86911 9488 86967 9544
rect 86991 9488 87047 9544
rect 87071 9488 87127 9544
rect 86831 7684 86887 7740
rect 86911 7684 86967 7740
rect 86991 7684 87047 7740
rect 87071 7684 87127 7740
rect 86831 7642 86887 7660
rect 86911 7642 86967 7660
rect 86991 7642 87047 7660
rect 87071 7642 87127 7660
rect 86831 7604 86877 7642
rect 86877 7604 86887 7642
rect 86911 7604 86941 7642
rect 86941 7604 86953 7642
rect 86953 7604 86967 7642
rect 86991 7604 87005 7642
rect 87005 7604 87017 7642
rect 87017 7604 87047 7642
rect 87071 7604 87081 7642
rect 87081 7604 87127 7642
rect 86831 7524 86887 7580
rect 86911 7524 86967 7580
rect 86991 7524 87047 7580
rect 87071 7524 87127 7580
rect 86831 7444 86887 7500
rect 86911 7444 86967 7500
rect 86991 7444 87047 7500
rect 87071 7444 87127 7500
rect 256601 9068 256657 9124
rect 256681 9068 256737 9124
rect 256761 9068 256817 9124
rect 256841 9068 256897 9124
rect 256601 8988 256657 9044
rect 256681 8988 256737 9044
rect 256761 8988 256817 9044
rect 256841 8988 256897 9044
rect 256601 8908 256657 8964
rect 256681 8908 256737 8964
rect 256761 8908 256817 8964
rect 256841 8908 256897 8964
rect 256601 8828 256657 8884
rect 256681 8828 256737 8884
rect 256761 8828 256817 8884
rect 256841 8828 256897 8884
rect 256601 7046 256647 7080
rect 256647 7046 256657 7080
rect 256681 7046 256711 7080
rect 256711 7046 256723 7080
rect 256723 7046 256737 7080
rect 256761 7046 256775 7080
rect 256775 7046 256787 7080
rect 256787 7046 256817 7080
rect 256841 7046 256851 7080
rect 256851 7046 256897 7080
rect 256601 7024 256657 7046
rect 256681 7024 256737 7046
rect 256761 7024 256817 7046
rect 256841 7024 256897 7046
rect 256601 6944 256657 7000
rect 256681 6944 256737 7000
rect 256761 6944 256817 7000
rect 256841 6944 256897 7000
rect 256601 6864 256657 6920
rect 256681 6864 256737 6920
rect 256761 6864 256817 6920
rect 256841 6864 256897 6920
rect 86831 6325 86887 6381
rect 86911 6325 86967 6381
rect 86991 6325 87047 6381
rect 87071 6325 87127 6381
rect 86831 6245 86887 6301
rect 86911 6245 86967 6301
rect 86991 6245 87047 6301
rect 87071 6245 87127 6301
rect 86831 6165 86887 6221
rect 86911 6165 86967 6221
rect 86991 6165 87047 6221
rect 87071 6165 87127 6221
rect 86831 6085 86887 6141
rect 86911 6085 86967 6141
rect 86991 6085 87047 6141
rect 87071 6085 87127 6141
rect 86831 4966 86887 5022
rect 86911 4966 86967 5022
rect 86991 4966 87047 5022
rect 87071 4966 87127 5022
rect 86831 4886 86887 4942
rect 86911 4886 86967 4942
rect 86991 4886 87047 4942
rect 87071 4886 87127 4942
rect 86831 4806 86887 4862
rect 86911 4806 86967 4862
rect 86991 4806 87047 4862
rect 87071 4806 87127 4862
rect 86831 4726 86887 4782
rect 86911 4726 86967 4782
rect 86991 4726 87047 4782
rect 87071 4726 87127 4782
rect 86831 3607 86887 3663
rect 86911 3607 86967 3663
rect 86991 3607 87047 3663
rect 87071 3607 87127 3663
rect 86831 3527 86887 3583
rect 86911 3527 86967 3583
rect 86991 3527 87047 3583
rect 87071 3527 87127 3583
rect 86831 3447 86887 3503
rect 86911 3447 86967 3503
rect 86991 3447 87047 3503
rect 87071 3447 87127 3503
rect 86831 3367 86887 3423
rect 86911 3367 86967 3423
rect 86991 3367 87047 3423
rect 87071 3367 87127 3423
rect 86831 248 86887 304
rect 86911 248 86967 304
rect 86991 248 87047 304
rect 87071 248 87127 304
rect 86831 168 86887 224
rect 86911 168 86967 224
rect 86991 168 87047 224
rect 87071 168 87127 224
rect 86831 88 86887 144
rect 86911 88 86967 144
rect 86991 88 87047 144
rect 87071 88 87127 144
rect 236826 2488 236882 2544
rect 227442 1148 227498 1184
rect 227442 1128 227444 1148
rect 227444 1128 227496 1148
rect 227496 1128 227498 1148
rect 229466 1128 229522 1184
rect 239954 1400 240010 1456
rect 242070 1672 242126 1728
rect 241794 1536 241850 1592
rect 244002 1420 244058 1456
rect 244002 1400 244004 1420
rect 244004 1400 244056 1420
rect 244056 1400 244058 1420
rect 244002 1148 244058 1184
rect 244278 1400 244334 1456
rect 244830 1536 244886 1592
rect 244002 1128 244004 1148
rect 244004 1128 244056 1148
rect 244056 1128 244058 1148
rect 244554 1300 244556 1320
rect 244556 1300 244608 1320
rect 244608 1300 244610 1320
rect 244554 1264 244610 1300
rect 244646 1128 244702 1184
rect 243634 448 243690 504
rect 244462 448 244518 504
rect 256601 6784 256657 6840
rect 256681 6784 256737 6840
rect 256761 6784 256817 6840
rect 256841 6784 256897 6840
rect 256601 5665 256657 5721
rect 256681 5665 256737 5721
rect 256761 5665 256817 5721
rect 256841 5665 256897 5721
rect 256601 5585 256657 5641
rect 256681 5585 256737 5641
rect 256761 5585 256817 5641
rect 256841 5585 256897 5641
rect 256601 5505 256657 5561
rect 256681 5505 256737 5561
rect 256761 5505 256817 5561
rect 256841 5505 256897 5561
rect 256601 5425 256657 5481
rect 256681 5425 256737 5481
rect 256761 5425 256817 5481
rect 256841 5425 256897 5481
rect 256601 4306 256657 4362
rect 256681 4306 256737 4362
rect 256761 4306 256817 4362
rect 256841 4306 256897 4362
rect 256601 4226 256657 4282
rect 256681 4226 256737 4282
rect 256761 4226 256817 4282
rect 256841 4226 256897 4282
rect 256601 4146 256657 4202
rect 256681 4146 256737 4202
rect 256761 4146 256817 4202
rect 256841 4146 256897 4202
rect 256601 4066 256657 4122
rect 256681 4066 256737 4122
rect 256761 4066 256817 4122
rect 256841 4066 256897 4122
rect 256601 2947 256657 3003
rect 256681 2947 256737 3003
rect 256761 2947 256817 3003
rect 256841 2947 256897 3003
rect 256601 2867 256657 2923
rect 256681 2867 256737 2923
rect 256761 2867 256817 2923
rect 256841 2867 256897 2923
rect 256601 2787 256657 2843
rect 256681 2787 256737 2843
rect 256761 2787 256817 2843
rect 256841 2787 256897 2843
rect 256601 2746 256657 2763
rect 256681 2746 256737 2763
rect 256761 2746 256817 2763
rect 256841 2746 256897 2763
rect 256601 2707 256647 2746
rect 256647 2707 256657 2746
rect 256681 2707 256711 2746
rect 256711 2707 256723 2746
rect 256723 2707 256737 2746
rect 256761 2707 256775 2746
rect 256775 2707 256787 2746
rect 256787 2707 256817 2746
rect 256841 2707 256851 2746
rect 256851 2707 256897 2746
rect 249430 1672 249486 1728
rect 248418 1400 248474 1456
rect 246394 1264 246450 1320
rect 256601 908 256657 964
rect 256681 908 256737 964
rect 256761 908 256817 964
rect 256841 908 256897 964
rect 256601 828 256657 884
rect 256681 828 256737 884
rect 256761 828 256817 884
rect 256841 828 256897 884
rect 256601 748 256657 804
rect 256681 748 256737 804
rect 256761 748 256817 804
rect 256841 748 256897 804
rect 256601 668 256657 724
rect 256681 668 256737 724
rect 256761 668 256817 724
rect 256841 668 256897 724
rect 86831 8 86887 64
rect 86911 8 86967 64
rect 86991 8 87047 64
rect 87071 8 87127 64
rect 257261 9728 257317 9784
rect 257341 9728 257397 9784
rect 257421 9728 257477 9784
rect 257501 9728 257557 9784
rect 257261 9648 257317 9704
rect 257341 9648 257397 9704
rect 257421 9648 257477 9704
rect 257501 9648 257557 9704
rect 257261 9568 257317 9624
rect 257341 9568 257397 9624
rect 257421 9568 257477 9624
rect 257501 9568 257557 9624
rect 257261 9488 257317 9544
rect 257341 9488 257397 9544
rect 257421 9488 257477 9544
rect 257501 9488 257557 9544
rect 257261 7684 257317 7740
rect 257341 7684 257397 7740
rect 257421 7684 257477 7740
rect 257501 7684 257557 7740
rect 257261 7642 257317 7660
rect 257341 7642 257397 7660
rect 257421 7642 257477 7660
rect 257501 7642 257557 7660
rect 257261 7604 257307 7642
rect 257307 7604 257317 7642
rect 257341 7604 257371 7642
rect 257371 7604 257383 7642
rect 257383 7604 257397 7642
rect 257421 7604 257435 7642
rect 257435 7604 257447 7642
rect 257447 7604 257477 7642
rect 257501 7604 257511 7642
rect 257511 7604 257557 7642
rect 257261 7524 257317 7580
rect 257341 7524 257397 7580
rect 257421 7524 257477 7580
rect 257501 7524 257557 7580
rect 257261 7444 257317 7500
rect 257341 7444 257397 7500
rect 257421 7444 257477 7500
rect 257501 7444 257557 7500
rect 257261 6325 257317 6381
rect 257341 6325 257397 6381
rect 257421 6325 257477 6381
rect 257501 6325 257557 6381
rect 257261 6245 257317 6301
rect 257341 6245 257397 6301
rect 257421 6245 257477 6301
rect 257501 6245 257557 6301
rect 257261 6165 257317 6221
rect 257341 6165 257397 6221
rect 257421 6165 257477 6221
rect 257501 6165 257557 6221
rect 257261 6085 257317 6141
rect 257341 6085 257397 6141
rect 257421 6085 257477 6141
rect 257501 6085 257557 6141
rect 257261 4966 257317 5022
rect 257341 4966 257397 5022
rect 257421 4966 257477 5022
rect 257501 4966 257557 5022
rect 257261 4886 257317 4942
rect 257341 4886 257397 4942
rect 257421 4886 257477 4942
rect 257501 4886 257557 4942
rect 257261 4806 257317 4862
rect 257341 4806 257397 4862
rect 257421 4806 257477 4862
rect 257501 4806 257557 4862
rect 257261 4726 257317 4782
rect 257341 4726 257397 4782
rect 257421 4726 257477 4782
rect 257501 4726 257557 4782
rect 257261 3607 257317 3663
rect 257341 3607 257397 3663
rect 257421 3607 257477 3663
rect 257501 3607 257557 3663
rect 257261 3527 257317 3583
rect 257341 3527 257397 3583
rect 257421 3527 257477 3583
rect 257501 3527 257557 3583
rect 257261 3447 257317 3503
rect 257341 3447 257397 3503
rect 257421 3447 257477 3503
rect 257501 3447 257557 3503
rect 257261 3367 257317 3423
rect 257341 3367 257397 3423
rect 257421 3367 257477 3423
rect 257501 3367 257557 3423
rect 257261 248 257317 304
rect 257341 248 257397 304
rect 257421 248 257477 304
rect 257501 248 257557 304
rect 326158 2488 326214 2544
rect 257261 168 257317 224
rect 257341 168 257397 224
rect 257421 168 257477 224
rect 257501 168 257557 224
rect 257261 88 257317 144
rect 257341 88 257397 144
rect 257421 88 257477 144
rect 257501 88 257557 144
rect 337014 2372 337070 2408
rect 337014 2352 337016 2372
rect 337016 2352 337068 2372
rect 337068 2352 337070 2372
rect 427031 9068 427087 9124
rect 427111 9068 427167 9124
rect 427191 9068 427247 9124
rect 427271 9068 427327 9124
rect 427031 8988 427087 9044
rect 427111 8988 427167 9044
rect 427191 8988 427247 9044
rect 427271 8988 427327 9044
rect 427031 8908 427087 8964
rect 427111 8908 427167 8964
rect 427191 8908 427247 8964
rect 427271 8908 427327 8964
rect 427031 8828 427087 8884
rect 427111 8828 427167 8884
rect 427191 8828 427247 8884
rect 427271 8828 427327 8884
rect 427031 7046 427077 7080
rect 427077 7046 427087 7080
rect 427111 7046 427141 7080
rect 427141 7046 427153 7080
rect 427153 7046 427167 7080
rect 427191 7046 427205 7080
rect 427205 7046 427217 7080
rect 427217 7046 427247 7080
rect 427271 7046 427281 7080
rect 427281 7046 427327 7080
rect 427031 7024 427087 7046
rect 427111 7024 427167 7046
rect 427191 7024 427247 7046
rect 427271 7024 427327 7046
rect 427031 6944 427087 7000
rect 427111 6944 427167 7000
rect 427191 6944 427247 7000
rect 427271 6944 427327 7000
rect 427031 6864 427087 6920
rect 427111 6864 427167 6920
rect 427191 6864 427247 6920
rect 427271 6864 427327 6920
rect 427031 6784 427087 6840
rect 427111 6784 427167 6840
rect 427191 6784 427247 6840
rect 427271 6784 427327 6840
rect 427031 5665 427087 5721
rect 427111 5665 427167 5721
rect 427191 5665 427247 5721
rect 427271 5665 427327 5721
rect 427031 5585 427087 5641
rect 427111 5585 427167 5641
rect 427191 5585 427247 5641
rect 427271 5585 427327 5641
rect 427031 5505 427087 5561
rect 427111 5505 427167 5561
rect 427191 5505 427247 5561
rect 427271 5505 427327 5561
rect 427031 5425 427087 5481
rect 427111 5425 427167 5481
rect 427191 5425 427247 5481
rect 427271 5425 427327 5481
rect 427031 4306 427087 4362
rect 427111 4306 427167 4362
rect 427191 4306 427247 4362
rect 427271 4306 427327 4362
rect 427031 4226 427087 4282
rect 427111 4226 427167 4282
rect 427191 4226 427247 4282
rect 427271 4226 427327 4282
rect 427031 4146 427087 4202
rect 427111 4146 427167 4202
rect 427191 4146 427247 4202
rect 427271 4146 427327 4202
rect 427031 4066 427087 4122
rect 427111 4066 427167 4122
rect 427191 4066 427247 4122
rect 427271 4066 427327 4122
rect 427031 2947 427087 3003
rect 427111 2947 427167 3003
rect 427191 2947 427247 3003
rect 427271 2947 427327 3003
rect 427031 2867 427087 2923
rect 427111 2867 427167 2923
rect 427191 2867 427247 2923
rect 427271 2867 427327 2923
rect 427031 2787 427087 2843
rect 427111 2787 427167 2843
rect 427191 2787 427247 2843
rect 427271 2787 427327 2843
rect 427031 2746 427087 2763
rect 427111 2746 427167 2763
rect 427191 2746 427247 2763
rect 427271 2746 427327 2763
rect 427031 2707 427077 2746
rect 427077 2707 427087 2746
rect 427111 2707 427141 2746
rect 427141 2707 427153 2746
rect 427153 2707 427167 2746
rect 427191 2707 427205 2746
rect 427205 2707 427217 2746
rect 427217 2707 427247 2746
rect 427271 2707 427281 2746
rect 427281 2707 427327 2746
rect 427031 908 427087 964
rect 427111 908 427167 964
rect 427191 908 427247 964
rect 427271 908 427327 964
rect 427031 828 427087 884
rect 427111 828 427167 884
rect 427191 828 427247 884
rect 427271 828 427327 884
rect 427031 748 427087 804
rect 427111 748 427167 804
rect 427191 748 427247 804
rect 427271 748 427327 804
rect 427031 668 427087 724
rect 427111 668 427167 724
rect 427191 668 427247 724
rect 427271 668 427327 724
rect 257261 8 257317 64
rect 257341 8 257397 64
rect 257421 8 257477 64
rect 257501 8 257557 64
rect 427691 9728 427747 9784
rect 427771 9728 427827 9784
rect 427851 9728 427907 9784
rect 427931 9728 427987 9784
rect 427691 9648 427747 9704
rect 427771 9648 427827 9704
rect 427851 9648 427907 9704
rect 427931 9648 427987 9704
rect 427691 9568 427747 9624
rect 427771 9568 427827 9624
rect 427851 9568 427907 9624
rect 427931 9568 427987 9624
rect 427691 9488 427747 9544
rect 427771 9488 427827 9544
rect 427851 9488 427907 9544
rect 427931 9488 427987 9544
rect 427691 7684 427747 7740
rect 427771 7684 427827 7740
rect 427851 7684 427907 7740
rect 427931 7684 427987 7740
rect 427691 7642 427747 7660
rect 427771 7642 427827 7660
rect 427851 7642 427907 7660
rect 427931 7642 427987 7660
rect 427691 7604 427737 7642
rect 427737 7604 427747 7642
rect 427771 7604 427801 7642
rect 427801 7604 427813 7642
rect 427813 7604 427827 7642
rect 427851 7604 427865 7642
rect 427865 7604 427877 7642
rect 427877 7604 427907 7642
rect 427931 7604 427941 7642
rect 427941 7604 427987 7642
rect 427691 7524 427747 7580
rect 427771 7524 427827 7580
rect 427851 7524 427907 7580
rect 427931 7524 427987 7580
rect 427691 7444 427747 7500
rect 427771 7444 427827 7500
rect 427851 7444 427907 7500
rect 427931 7444 427987 7500
rect 427691 6325 427747 6381
rect 427771 6325 427827 6381
rect 427851 6325 427907 6381
rect 427931 6325 427987 6381
rect 427691 6245 427747 6301
rect 427771 6245 427827 6301
rect 427851 6245 427907 6301
rect 427931 6245 427987 6301
rect 427691 6165 427747 6221
rect 427771 6165 427827 6221
rect 427851 6165 427907 6221
rect 427931 6165 427987 6221
rect 427691 6085 427747 6141
rect 427771 6085 427827 6141
rect 427851 6085 427907 6141
rect 427931 6085 427987 6141
rect 427691 4966 427747 5022
rect 427771 4966 427827 5022
rect 427851 4966 427907 5022
rect 427931 4966 427987 5022
rect 427691 4886 427747 4942
rect 427771 4886 427827 4942
rect 427851 4886 427907 4942
rect 427931 4886 427987 4942
rect 427691 4806 427747 4862
rect 427771 4806 427827 4862
rect 427851 4806 427907 4862
rect 427931 4806 427987 4862
rect 427691 4726 427747 4782
rect 427771 4726 427827 4782
rect 427851 4726 427907 4782
rect 427931 4726 427987 4782
rect 427691 3607 427747 3663
rect 427771 3607 427827 3663
rect 427851 3607 427907 3663
rect 427931 3607 427987 3663
rect 427691 3527 427747 3583
rect 427771 3527 427827 3583
rect 427851 3527 427907 3583
rect 427931 3527 427987 3583
rect 427691 3447 427747 3503
rect 427771 3447 427827 3503
rect 427851 3447 427907 3503
rect 427931 3447 427987 3503
rect 427691 3367 427747 3423
rect 427771 3367 427827 3423
rect 427851 3367 427907 3423
rect 427931 3367 427987 3423
rect 431866 2488 431922 2544
rect 430762 2352 430818 2408
rect 525062 2524 525064 2544
rect 525064 2524 525116 2544
rect 525116 2524 525118 2544
rect 525062 2488 525118 2524
rect 597461 9068 597517 9124
rect 597541 9068 597597 9124
rect 597621 9068 597677 9124
rect 597701 9068 597757 9124
rect 597461 8988 597517 9044
rect 597541 8988 597597 9044
rect 597621 8988 597677 9044
rect 597701 8988 597757 9044
rect 597461 8908 597517 8964
rect 597541 8908 597597 8964
rect 597621 8908 597677 8964
rect 597701 8908 597757 8964
rect 597461 8828 597517 8884
rect 597541 8828 597597 8884
rect 597621 8828 597677 8884
rect 597701 8828 597757 8884
rect 597461 7046 597507 7080
rect 597507 7046 597517 7080
rect 597541 7046 597571 7080
rect 597571 7046 597583 7080
rect 597583 7046 597597 7080
rect 597621 7046 597635 7080
rect 597635 7046 597647 7080
rect 597647 7046 597677 7080
rect 597701 7046 597711 7080
rect 597711 7046 597757 7080
rect 597461 7024 597517 7046
rect 597541 7024 597597 7046
rect 597621 7024 597677 7046
rect 597701 7024 597757 7046
rect 597461 6944 597517 7000
rect 597541 6944 597597 7000
rect 597621 6944 597677 7000
rect 597701 6944 597757 7000
rect 597461 6864 597517 6920
rect 597541 6864 597597 6920
rect 597621 6864 597677 6920
rect 597701 6864 597757 6920
rect 597461 6784 597517 6840
rect 597541 6784 597597 6840
rect 597621 6784 597677 6840
rect 597701 6784 597757 6840
rect 597461 5665 597517 5721
rect 597541 5665 597597 5721
rect 597621 5665 597677 5721
rect 597701 5665 597757 5721
rect 597461 5585 597517 5641
rect 597541 5585 597597 5641
rect 597621 5585 597677 5641
rect 597701 5585 597757 5641
rect 597461 5505 597517 5561
rect 597541 5505 597597 5561
rect 597621 5505 597677 5561
rect 597701 5505 597757 5561
rect 597461 5425 597517 5481
rect 597541 5425 597597 5481
rect 597621 5425 597677 5481
rect 597701 5425 597757 5481
rect 597461 4306 597517 4362
rect 597541 4306 597597 4362
rect 597621 4306 597677 4362
rect 597701 4306 597757 4362
rect 597461 4226 597517 4282
rect 597541 4226 597597 4282
rect 597621 4226 597677 4282
rect 597701 4226 597757 4282
rect 597461 4146 597517 4202
rect 597541 4146 597597 4202
rect 597621 4146 597677 4202
rect 597701 4146 597757 4202
rect 597461 4066 597517 4122
rect 597541 4066 597597 4122
rect 597621 4066 597677 4122
rect 597701 4066 597757 4122
rect 597461 2947 597517 3003
rect 597541 2947 597597 3003
rect 597621 2947 597677 3003
rect 597701 2947 597757 3003
rect 597461 2867 597517 2923
rect 597541 2867 597597 2923
rect 597621 2867 597677 2923
rect 597701 2867 597757 2923
rect 597461 2787 597517 2843
rect 597541 2787 597597 2843
rect 597621 2787 597677 2843
rect 597701 2787 597757 2843
rect 597461 2746 597517 2763
rect 597541 2746 597597 2763
rect 597621 2746 597677 2763
rect 597701 2746 597757 2763
rect 597461 2707 597507 2746
rect 597507 2707 597517 2746
rect 597541 2707 597571 2746
rect 597571 2707 597583 2746
rect 597583 2707 597597 2746
rect 597621 2707 597635 2746
rect 597635 2707 597647 2746
rect 597647 2707 597677 2746
rect 597701 2707 597711 2746
rect 597711 2707 597757 2746
rect 427691 248 427747 304
rect 427771 248 427827 304
rect 427851 248 427907 304
rect 427931 248 427987 304
rect 427691 168 427747 224
rect 427771 168 427827 224
rect 427851 168 427907 224
rect 427931 168 427987 224
rect 427691 88 427747 144
rect 427771 88 427827 144
rect 427851 88 427907 144
rect 427931 88 427987 144
rect 427691 8 427747 64
rect 427771 8 427827 64
rect 427851 8 427907 64
rect 427931 8 427987 64
rect 597461 908 597517 964
rect 597541 908 597597 964
rect 597621 908 597677 964
rect 597701 908 597757 964
rect 597461 828 597517 884
rect 597541 828 597597 884
rect 597621 828 597677 884
rect 597701 828 597757 884
rect 597461 748 597517 804
rect 597541 748 597597 804
rect 597621 748 597677 804
rect 597701 748 597757 804
rect 597461 668 597517 724
rect 597541 668 597597 724
rect 597621 668 597677 724
rect 597701 668 597757 724
rect 598121 9728 598177 9784
rect 598201 9728 598257 9784
rect 598281 9728 598337 9784
rect 598361 9728 598417 9784
rect 598121 9648 598177 9704
rect 598201 9648 598257 9704
rect 598281 9648 598337 9704
rect 598361 9648 598417 9704
rect 598121 9568 598177 9624
rect 598201 9568 598257 9624
rect 598281 9568 598337 9624
rect 598361 9568 598417 9624
rect 598121 9488 598177 9544
rect 598201 9488 598257 9544
rect 598281 9488 598337 9544
rect 598361 9488 598417 9544
rect 684696 9728 684752 9784
rect 684776 9728 684832 9784
rect 684856 9728 684912 9784
rect 684936 9728 684992 9784
rect 684696 9648 684752 9704
rect 684776 9648 684832 9704
rect 684856 9648 684912 9704
rect 684936 9648 684992 9704
rect 684696 9568 684752 9624
rect 684776 9568 684832 9624
rect 684856 9568 684912 9624
rect 684936 9568 684992 9624
rect 684696 9488 684752 9544
rect 684776 9488 684832 9544
rect 684856 9488 684912 9544
rect 684936 9488 684992 9544
rect 598121 7684 598177 7740
rect 598201 7684 598257 7740
rect 598281 7684 598337 7740
rect 598361 7684 598417 7740
rect 598121 7642 598177 7660
rect 598201 7642 598257 7660
rect 598281 7642 598337 7660
rect 598361 7642 598417 7660
rect 598121 7604 598167 7642
rect 598167 7604 598177 7642
rect 598201 7604 598231 7642
rect 598231 7604 598243 7642
rect 598243 7604 598257 7642
rect 598281 7604 598295 7642
rect 598295 7604 598307 7642
rect 598307 7604 598337 7642
rect 598361 7604 598371 7642
rect 598371 7604 598417 7642
rect 598121 7524 598177 7580
rect 598201 7524 598257 7580
rect 598281 7524 598337 7580
rect 598361 7524 598417 7580
rect 598121 7444 598177 7500
rect 598201 7444 598257 7500
rect 598281 7444 598337 7500
rect 598361 7444 598417 7500
rect 598121 6325 598177 6381
rect 598201 6325 598257 6381
rect 598281 6325 598337 6381
rect 598361 6325 598417 6381
rect 598121 6245 598177 6301
rect 598201 6245 598257 6301
rect 598281 6245 598337 6301
rect 598361 6245 598417 6301
rect 598121 6165 598177 6221
rect 598201 6165 598257 6221
rect 598281 6165 598337 6221
rect 598361 6165 598417 6221
rect 598121 6085 598177 6141
rect 598201 6085 598257 6141
rect 598281 6085 598337 6141
rect 598361 6085 598417 6141
rect 598121 4966 598177 5022
rect 598201 4966 598257 5022
rect 598281 4966 598337 5022
rect 598361 4966 598417 5022
rect 598121 4886 598177 4942
rect 598201 4886 598257 4942
rect 598281 4886 598337 4942
rect 598361 4886 598417 4942
rect 598121 4806 598177 4862
rect 598201 4806 598257 4862
rect 598281 4806 598337 4862
rect 598361 4806 598417 4862
rect 598121 4726 598177 4782
rect 598201 4726 598257 4782
rect 598281 4726 598337 4782
rect 598361 4726 598417 4782
rect 598121 3607 598177 3663
rect 598201 3607 598257 3663
rect 598281 3607 598337 3663
rect 598361 3607 598417 3663
rect 598121 3527 598177 3583
rect 598201 3527 598257 3583
rect 598281 3527 598337 3583
rect 598361 3527 598417 3583
rect 598121 3447 598177 3503
rect 598201 3447 598257 3503
rect 598281 3447 598337 3503
rect 598361 3447 598417 3503
rect 598121 3367 598177 3423
rect 598201 3367 598257 3423
rect 598281 3367 598337 3423
rect 598361 3367 598417 3423
rect 684036 9068 684092 9124
rect 684116 9068 684172 9124
rect 684196 9068 684252 9124
rect 684276 9068 684332 9124
rect 684036 8988 684092 9044
rect 684116 8988 684172 9044
rect 684196 8988 684252 9044
rect 684276 8988 684332 9044
rect 684036 8908 684092 8964
rect 684116 8908 684172 8964
rect 684196 8908 684252 8964
rect 684276 8908 684332 8964
rect 684036 8828 684092 8884
rect 684116 8828 684172 8884
rect 684196 8828 684252 8884
rect 684276 8828 684332 8884
rect 684036 7024 684092 7080
rect 684116 7024 684172 7080
rect 684196 7024 684252 7080
rect 684276 7024 684332 7080
rect 684036 6944 684092 7000
rect 684116 6944 684172 7000
rect 684196 6944 684252 7000
rect 684276 6944 684332 7000
rect 684036 6864 684092 6920
rect 684116 6864 684172 6920
rect 684196 6864 684252 6920
rect 684276 6864 684332 6920
rect 684036 6784 684092 6840
rect 684116 6784 684172 6840
rect 684196 6784 684252 6840
rect 684276 6784 684332 6840
rect 684036 5665 684092 5721
rect 684116 5665 684172 5721
rect 684196 5665 684252 5721
rect 684276 5665 684332 5721
rect 684036 5585 684092 5641
rect 684116 5585 684172 5641
rect 684196 5585 684252 5641
rect 684276 5585 684332 5641
rect 684036 5505 684092 5561
rect 684116 5505 684172 5561
rect 684196 5505 684252 5561
rect 684276 5505 684332 5561
rect 684036 5425 684092 5481
rect 684116 5425 684172 5481
rect 684196 5425 684252 5481
rect 684276 5425 684332 5481
rect 684036 4306 684092 4362
rect 684116 4306 684172 4362
rect 684196 4306 684252 4362
rect 684276 4306 684332 4362
rect 684036 4226 684092 4282
rect 684116 4226 684172 4282
rect 684196 4226 684252 4282
rect 684276 4226 684332 4282
rect 684036 4146 684092 4202
rect 684116 4146 684172 4202
rect 684196 4146 684252 4202
rect 684276 4146 684332 4202
rect 684036 4066 684092 4122
rect 684116 4066 684172 4122
rect 684196 4066 684252 4122
rect 684276 4066 684332 4122
rect 684036 2947 684092 3003
rect 684116 2947 684172 3003
rect 684196 2947 684252 3003
rect 684276 2947 684332 3003
rect 684036 2867 684092 2923
rect 684116 2867 684172 2923
rect 684196 2867 684252 2923
rect 684276 2867 684332 2923
rect 684036 2787 684092 2843
rect 684116 2787 684172 2843
rect 684196 2787 684252 2843
rect 684276 2787 684332 2843
rect 684036 2707 684092 2763
rect 684116 2707 684172 2763
rect 684196 2707 684252 2763
rect 684276 2707 684332 2763
rect 684036 908 684092 964
rect 684116 908 684172 964
rect 684196 908 684252 964
rect 684276 908 684332 964
rect 684036 828 684092 884
rect 684116 828 684172 884
rect 684196 828 684252 884
rect 684276 828 684332 884
rect 684036 748 684092 804
rect 684116 748 684172 804
rect 684196 748 684252 804
rect 684276 748 684332 804
rect 684036 668 684092 724
rect 684116 668 684172 724
rect 684196 668 684252 724
rect 684276 668 684332 724
rect 684696 7684 684752 7740
rect 684776 7684 684832 7740
rect 684856 7684 684912 7740
rect 684936 7684 684992 7740
rect 684696 7604 684752 7660
rect 684776 7604 684832 7660
rect 684856 7604 684912 7660
rect 684936 7604 684992 7660
rect 684696 7524 684752 7580
rect 684776 7524 684832 7580
rect 684856 7524 684912 7580
rect 684936 7524 684992 7580
rect 684696 7444 684752 7500
rect 684776 7444 684832 7500
rect 684856 7444 684912 7500
rect 684936 7444 684992 7500
rect 684696 6325 684752 6381
rect 684776 6325 684832 6381
rect 684856 6325 684912 6381
rect 684936 6325 684992 6381
rect 684696 6245 684752 6301
rect 684776 6245 684832 6301
rect 684856 6245 684912 6301
rect 684936 6245 684992 6301
rect 684696 6165 684752 6221
rect 684776 6165 684832 6221
rect 684856 6165 684912 6221
rect 684936 6165 684992 6221
rect 684696 6085 684752 6141
rect 684776 6085 684832 6141
rect 684856 6085 684912 6141
rect 684936 6085 684992 6141
rect 684696 4966 684752 5022
rect 684776 4966 684832 5022
rect 684856 4966 684912 5022
rect 684936 4966 684992 5022
rect 684696 4886 684752 4942
rect 684776 4886 684832 4942
rect 684856 4886 684912 4942
rect 684936 4886 684992 4942
rect 684696 4806 684752 4862
rect 684776 4806 684832 4862
rect 684856 4806 684912 4862
rect 684936 4806 684992 4862
rect 684696 4726 684752 4782
rect 684776 4726 684832 4782
rect 684856 4726 684912 4782
rect 684936 4726 684992 4782
rect 684696 3607 684752 3663
rect 684776 3607 684832 3663
rect 684856 3607 684912 3663
rect 684936 3607 684992 3663
rect 684696 3527 684752 3583
rect 684776 3527 684832 3583
rect 684856 3527 684912 3583
rect 684936 3527 684992 3583
rect 684696 3447 684752 3503
rect 684776 3447 684832 3503
rect 684856 3447 684912 3503
rect 684936 3447 684992 3503
rect 684696 3367 684752 3423
rect 684776 3367 684832 3423
rect 684856 3367 684912 3423
rect 684936 3367 684992 3423
rect 598121 248 598177 304
rect 598201 248 598257 304
rect 598281 248 598337 304
rect 598361 248 598417 304
rect 598121 168 598177 224
rect 598201 168 598257 224
rect 598281 168 598337 224
rect 598361 168 598417 224
rect 598121 88 598177 144
rect 598201 88 598257 144
rect 598281 88 598337 144
rect 598361 88 598417 144
rect 598121 8 598177 64
rect 598201 8 598257 64
rect 598281 8 598337 64
rect 598361 8 598417 64
rect 684696 248 684752 304
rect 684776 248 684832 304
rect 684856 248 684912 304
rect 684936 248 684992 304
rect 684696 168 684752 224
rect 684776 168 684832 224
rect 684856 168 684912 224
rect 684936 168 684992 224
rect 684696 88 684752 144
rect 684776 88 684832 144
rect 684856 88 684912 144
rect 684936 88 684992 144
rect 684696 8 684752 64
rect 684776 8 684832 64
rect 684856 8 684912 64
rect 684936 8 684992 64
<< metal3 >>
rect -1076 9784 685004 9796
rect -1076 9728 -1064 9784
rect -1008 9728 -984 9784
rect -928 9728 -904 9784
rect -848 9728 -824 9784
rect -768 9728 86831 9784
rect 86887 9728 86911 9784
rect 86967 9728 86991 9784
rect 87047 9728 87071 9784
rect 87127 9728 257261 9784
rect 257317 9728 257341 9784
rect 257397 9728 257421 9784
rect 257477 9728 257501 9784
rect 257557 9728 427691 9784
rect 427747 9728 427771 9784
rect 427827 9728 427851 9784
rect 427907 9728 427931 9784
rect 427987 9728 598121 9784
rect 598177 9728 598201 9784
rect 598257 9728 598281 9784
rect 598337 9728 598361 9784
rect 598417 9728 684696 9784
rect 684752 9728 684776 9784
rect 684832 9728 684856 9784
rect 684912 9728 684936 9784
rect 684992 9728 685004 9784
rect -1076 9704 685004 9728
rect -1076 9648 -1064 9704
rect -1008 9648 -984 9704
rect -928 9648 -904 9704
rect -848 9648 -824 9704
rect -768 9648 86831 9704
rect 86887 9648 86911 9704
rect 86967 9648 86991 9704
rect 87047 9648 87071 9704
rect 87127 9648 257261 9704
rect 257317 9648 257341 9704
rect 257397 9648 257421 9704
rect 257477 9648 257501 9704
rect 257557 9648 427691 9704
rect 427747 9648 427771 9704
rect 427827 9648 427851 9704
rect 427907 9648 427931 9704
rect 427987 9648 598121 9704
rect 598177 9648 598201 9704
rect 598257 9648 598281 9704
rect 598337 9648 598361 9704
rect 598417 9648 684696 9704
rect 684752 9648 684776 9704
rect 684832 9648 684856 9704
rect 684912 9648 684936 9704
rect 684992 9648 685004 9704
rect -1076 9624 685004 9648
rect -1076 9568 -1064 9624
rect -1008 9568 -984 9624
rect -928 9568 -904 9624
rect -848 9568 -824 9624
rect -768 9568 86831 9624
rect 86887 9568 86911 9624
rect 86967 9568 86991 9624
rect 87047 9568 87071 9624
rect 87127 9568 257261 9624
rect 257317 9568 257341 9624
rect 257397 9568 257421 9624
rect 257477 9568 257501 9624
rect 257557 9568 427691 9624
rect 427747 9568 427771 9624
rect 427827 9568 427851 9624
rect 427907 9568 427931 9624
rect 427987 9568 598121 9624
rect 598177 9568 598201 9624
rect 598257 9568 598281 9624
rect 598337 9568 598361 9624
rect 598417 9568 684696 9624
rect 684752 9568 684776 9624
rect 684832 9568 684856 9624
rect 684912 9568 684936 9624
rect 684992 9568 685004 9624
rect -1076 9544 685004 9568
rect -1076 9488 -1064 9544
rect -1008 9488 -984 9544
rect -928 9488 -904 9544
rect -848 9488 -824 9544
rect -768 9488 86831 9544
rect 86887 9488 86911 9544
rect 86967 9488 86991 9544
rect 87047 9488 87071 9544
rect 87127 9488 257261 9544
rect 257317 9488 257341 9544
rect 257397 9488 257421 9544
rect 257477 9488 257501 9544
rect 257557 9488 427691 9544
rect 427747 9488 427771 9544
rect 427827 9488 427851 9544
rect 427907 9488 427931 9544
rect 427987 9488 598121 9544
rect 598177 9488 598201 9544
rect 598257 9488 598281 9544
rect 598337 9488 598361 9544
rect 598417 9488 684696 9544
rect 684752 9488 684776 9544
rect 684832 9488 684856 9544
rect 684912 9488 684936 9544
rect 684992 9488 685004 9544
rect -1076 9476 685004 9488
rect -416 9124 684344 9136
rect -416 9068 -404 9124
rect -348 9068 -324 9124
rect -268 9068 -244 9124
rect -188 9068 -164 9124
rect -108 9068 86171 9124
rect 86227 9068 86251 9124
rect 86307 9068 86331 9124
rect 86387 9068 86411 9124
rect 86467 9068 256601 9124
rect 256657 9068 256681 9124
rect 256737 9068 256761 9124
rect 256817 9068 256841 9124
rect 256897 9068 427031 9124
rect 427087 9068 427111 9124
rect 427167 9068 427191 9124
rect 427247 9068 427271 9124
rect 427327 9068 597461 9124
rect 597517 9068 597541 9124
rect 597597 9068 597621 9124
rect 597677 9068 597701 9124
rect 597757 9068 684036 9124
rect 684092 9068 684116 9124
rect 684172 9068 684196 9124
rect 684252 9068 684276 9124
rect 684332 9068 684344 9124
rect -416 9044 684344 9068
rect -416 8988 -404 9044
rect -348 8988 -324 9044
rect -268 8988 -244 9044
rect -188 8988 -164 9044
rect -108 8988 86171 9044
rect 86227 8988 86251 9044
rect 86307 8988 86331 9044
rect 86387 8988 86411 9044
rect 86467 8988 256601 9044
rect 256657 8988 256681 9044
rect 256737 8988 256761 9044
rect 256817 8988 256841 9044
rect 256897 8988 427031 9044
rect 427087 8988 427111 9044
rect 427167 8988 427191 9044
rect 427247 8988 427271 9044
rect 427327 8988 597461 9044
rect 597517 8988 597541 9044
rect 597597 8988 597621 9044
rect 597677 8988 597701 9044
rect 597757 8988 684036 9044
rect 684092 8988 684116 9044
rect 684172 8988 684196 9044
rect 684252 8988 684276 9044
rect 684332 8988 684344 9044
rect -416 8964 684344 8988
rect -416 8908 -404 8964
rect -348 8908 -324 8964
rect -268 8908 -244 8964
rect -188 8908 -164 8964
rect -108 8908 86171 8964
rect 86227 8908 86251 8964
rect 86307 8908 86331 8964
rect 86387 8908 86411 8964
rect 86467 8908 256601 8964
rect 256657 8908 256681 8964
rect 256737 8908 256761 8964
rect 256817 8908 256841 8964
rect 256897 8908 427031 8964
rect 427087 8908 427111 8964
rect 427167 8908 427191 8964
rect 427247 8908 427271 8964
rect 427327 8908 597461 8964
rect 597517 8908 597541 8964
rect 597597 8908 597621 8964
rect 597677 8908 597701 8964
rect 597757 8908 684036 8964
rect 684092 8908 684116 8964
rect 684172 8908 684196 8964
rect 684252 8908 684276 8964
rect 684332 8908 684344 8964
rect -416 8884 684344 8908
rect -416 8828 -404 8884
rect -348 8828 -324 8884
rect -268 8828 -244 8884
rect -188 8828 -164 8884
rect -108 8828 86171 8884
rect 86227 8828 86251 8884
rect 86307 8828 86331 8884
rect 86387 8828 86411 8884
rect 86467 8828 256601 8884
rect 256657 8828 256681 8884
rect 256737 8828 256761 8884
rect 256817 8828 256841 8884
rect 256897 8828 427031 8884
rect 427087 8828 427111 8884
rect 427167 8828 427191 8884
rect 427247 8828 427271 8884
rect 427327 8828 597461 8884
rect 597517 8828 597541 8884
rect 597597 8828 597621 8884
rect 597677 8828 597701 8884
rect 597757 8828 684036 8884
rect 684092 8828 684116 8884
rect 684172 8828 684196 8884
rect 684252 8828 684276 8884
rect 684332 8828 684344 8884
rect -416 8816 684344 8828
rect -1076 7740 685004 7752
rect -1076 7684 -1064 7740
rect -1008 7684 -984 7740
rect -928 7684 -904 7740
rect -848 7684 -824 7740
rect -768 7684 86831 7740
rect 86887 7684 86911 7740
rect 86967 7684 86991 7740
rect 87047 7684 87071 7740
rect 87127 7684 257261 7740
rect 257317 7684 257341 7740
rect 257397 7684 257421 7740
rect 257477 7684 257501 7740
rect 257557 7684 427691 7740
rect 427747 7684 427771 7740
rect 427827 7684 427851 7740
rect 427907 7684 427931 7740
rect 427987 7684 598121 7740
rect 598177 7684 598201 7740
rect 598257 7684 598281 7740
rect 598337 7684 598361 7740
rect 598417 7684 684696 7740
rect 684752 7684 684776 7740
rect 684832 7684 684856 7740
rect 684912 7684 684936 7740
rect 684992 7684 685004 7740
rect -1076 7660 685004 7684
rect -1076 7604 -1064 7660
rect -1008 7604 -984 7660
rect -928 7604 -904 7660
rect -848 7604 -824 7660
rect -768 7604 86831 7660
rect 86887 7604 86911 7660
rect 86967 7604 86991 7660
rect 87047 7604 87071 7660
rect 87127 7604 257261 7660
rect 257317 7604 257341 7660
rect 257397 7604 257421 7660
rect 257477 7604 257501 7660
rect 257557 7604 427691 7660
rect 427747 7604 427771 7660
rect 427827 7604 427851 7660
rect 427907 7604 427931 7660
rect 427987 7604 598121 7660
rect 598177 7604 598201 7660
rect 598257 7604 598281 7660
rect 598337 7604 598361 7660
rect 598417 7604 684696 7660
rect 684752 7604 684776 7660
rect 684832 7604 684856 7660
rect 684912 7604 684936 7660
rect 684992 7604 685004 7660
rect -1076 7580 685004 7604
rect -1076 7524 -1064 7580
rect -1008 7524 -984 7580
rect -928 7524 -904 7580
rect -848 7524 -824 7580
rect -768 7524 86831 7580
rect 86887 7524 86911 7580
rect 86967 7524 86991 7580
rect 87047 7524 87071 7580
rect 87127 7524 257261 7580
rect 257317 7524 257341 7580
rect 257397 7524 257421 7580
rect 257477 7524 257501 7580
rect 257557 7524 427691 7580
rect 427747 7524 427771 7580
rect 427827 7524 427851 7580
rect 427907 7524 427931 7580
rect 427987 7524 598121 7580
rect 598177 7524 598201 7580
rect 598257 7524 598281 7580
rect 598337 7524 598361 7580
rect 598417 7524 684696 7580
rect 684752 7524 684776 7580
rect 684832 7524 684856 7580
rect 684912 7524 684936 7580
rect 684992 7524 685004 7580
rect -1076 7500 685004 7524
rect -1076 7444 -1064 7500
rect -1008 7444 -984 7500
rect -928 7444 -904 7500
rect -848 7444 -824 7500
rect -768 7444 86831 7500
rect 86887 7444 86911 7500
rect 86967 7444 86991 7500
rect 87047 7444 87071 7500
rect 87127 7444 257261 7500
rect 257317 7444 257341 7500
rect 257397 7444 257421 7500
rect 257477 7444 257501 7500
rect 257557 7444 427691 7500
rect 427747 7444 427771 7500
rect 427827 7444 427851 7500
rect 427907 7444 427931 7500
rect 427987 7444 598121 7500
rect 598177 7444 598201 7500
rect 598257 7444 598281 7500
rect 598337 7444 598361 7500
rect 598417 7444 684696 7500
rect 684752 7444 684776 7500
rect 684832 7444 684856 7500
rect 684912 7444 684936 7500
rect 684992 7444 685004 7500
rect -1076 7432 685004 7444
rect -1076 7080 685004 7092
rect -1076 7024 -404 7080
rect -348 7024 -324 7080
rect -268 7024 -244 7080
rect -188 7024 -164 7080
rect -108 7024 86171 7080
rect 86227 7024 86251 7080
rect 86307 7024 86331 7080
rect 86387 7024 86411 7080
rect 86467 7024 256601 7080
rect 256657 7024 256681 7080
rect 256737 7024 256761 7080
rect 256817 7024 256841 7080
rect 256897 7024 427031 7080
rect 427087 7024 427111 7080
rect 427167 7024 427191 7080
rect 427247 7024 427271 7080
rect 427327 7024 597461 7080
rect 597517 7024 597541 7080
rect 597597 7024 597621 7080
rect 597677 7024 597701 7080
rect 597757 7024 684036 7080
rect 684092 7024 684116 7080
rect 684172 7024 684196 7080
rect 684252 7024 684276 7080
rect 684332 7024 685004 7080
rect -1076 7000 685004 7024
rect -1076 6944 -404 7000
rect -348 6944 -324 7000
rect -268 6944 -244 7000
rect -188 6944 -164 7000
rect -108 6944 86171 7000
rect 86227 6944 86251 7000
rect 86307 6944 86331 7000
rect 86387 6944 86411 7000
rect 86467 6944 256601 7000
rect 256657 6944 256681 7000
rect 256737 6944 256761 7000
rect 256817 6944 256841 7000
rect 256897 6944 427031 7000
rect 427087 6944 427111 7000
rect 427167 6944 427191 7000
rect 427247 6944 427271 7000
rect 427327 6944 597461 7000
rect 597517 6944 597541 7000
rect 597597 6944 597621 7000
rect 597677 6944 597701 7000
rect 597757 6944 684036 7000
rect 684092 6944 684116 7000
rect 684172 6944 684196 7000
rect 684252 6944 684276 7000
rect 684332 6944 685004 7000
rect -1076 6920 685004 6944
rect -1076 6864 -404 6920
rect -348 6864 -324 6920
rect -268 6864 -244 6920
rect -188 6864 -164 6920
rect -108 6864 86171 6920
rect 86227 6864 86251 6920
rect 86307 6864 86331 6920
rect 86387 6864 86411 6920
rect 86467 6864 256601 6920
rect 256657 6864 256681 6920
rect 256737 6864 256761 6920
rect 256817 6864 256841 6920
rect 256897 6864 427031 6920
rect 427087 6864 427111 6920
rect 427167 6864 427191 6920
rect 427247 6864 427271 6920
rect 427327 6864 597461 6920
rect 597517 6864 597541 6920
rect 597597 6864 597621 6920
rect 597677 6864 597701 6920
rect 597757 6864 684036 6920
rect 684092 6864 684116 6920
rect 684172 6864 684196 6920
rect 684252 6864 684276 6920
rect 684332 6864 685004 6920
rect -1076 6840 685004 6864
rect -1076 6784 -404 6840
rect -348 6784 -324 6840
rect -268 6784 -244 6840
rect -188 6784 -164 6840
rect -108 6784 86171 6840
rect 86227 6784 86251 6840
rect 86307 6784 86331 6840
rect 86387 6784 86411 6840
rect 86467 6784 256601 6840
rect 256657 6784 256681 6840
rect 256737 6784 256761 6840
rect 256817 6784 256841 6840
rect 256897 6784 427031 6840
rect 427087 6784 427111 6840
rect 427167 6784 427191 6840
rect 427247 6784 427271 6840
rect 427327 6784 597461 6840
rect 597517 6784 597541 6840
rect 597597 6784 597621 6840
rect 597677 6784 597701 6840
rect 597757 6784 684036 6840
rect 684092 6784 684116 6840
rect 684172 6784 684196 6840
rect 684252 6784 684276 6840
rect 684332 6784 685004 6840
rect -1076 6772 685004 6784
rect -1076 6381 685004 6393
rect -1076 6325 -1064 6381
rect -1008 6325 -984 6381
rect -928 6325 -904 6381
rect -848 6325 -824 6381
rect -768 6325 86831 6381
rect 86887 6325 86911 6381
rect 86967 6325 86991 6381
rect 87047 6325 87071 6381
rect 87127 6325 257261 6381
rect 257317 6325 257341 6381
rect 257397 6325 257421 6381
rect 257477 6325 257501 6381
rect 257557 6325 427691 6381
rect 427747 6325 427771 6381
rect 427827 6325 427851 6381
rect 427907 6325 427931 6381
rect 427987 6325 598121 6381
rect 598177 6325 598201 6381
rect 598257 6325 598281 6381
rect 598337 6325 598361 6381
rect 598417 6325 684696 6381
rect 684752 6325 684776 6381
rect 684832 6325 684856 6381
rect 684912 6325 684936 6381
rect 684992 6325 685004 6381
rect -1076 6301 685004 6325
rect -1076 6245 -1064 6301
rect -1008 6245 -984 6301
rect -928 6245 -904 6301
rect -848 6245 -824 6301
rect -768 6245 86831 6301
rect 86887 6245 86911 6301
rect 86967 6245 86991 6301
rect 87047 6245 87071 6301
rect 87127 6245 257261 6301
rect 257317 6245 257341 6301
rect 257397 6245 257421 6301
rect 257477 6245 257501 6301
rect 257557 6245 427691 6301
rect 427747 6245 427771 6301
rect 427827 6245 427851 6301
rect 427907 6245 427931 6301
rect 427987 6245 598121 6301
rect 598177 6245 598201 6301
rect 598257 6245 598281 6301
rect 598337 6245 598361 6301
rect 598417 6245 684696 6301
rect 684752 6245 684776 6301
rect 684832 6245 684856 6301
rect 684912 6245 684936 6301
rect 684992 6245 685004 6301
rect -1076 6221 685004 6245
rect -1076 6165 -1064 6221
rect -1008 6165 -984 6221
rect -928 6165 -904 6221
rect -848 6165 -824 6221
rect -768 6165 86831 6221
rect 86887 6165 86911 6221
rect 86967 6165 86991 6221
rect 87047 6165 87071 6221
rect 87127 6165 257261 6221
rect 257317 6165 257341 6221
rect 257397 6165 257421 6221
rect 257477 6165 257501 6221
rect 257557 6165 427691 6221
rect 427747 6165 427771 6221
rect 427827 6165 427851 6221
rect 427907 6165 427931 6221
rect 427987 6165 598121 6221
rect 598177 6165 598201 6221
rect 598257 6165 598281 6221
rect 598337 6165 598361 6221
rect 598417 6165 684696 6221
rect 684752 6165 684776 6221
rect 684832 6165 684856 6221
rect 684912 6165 684936 6221
rect 684992 6165 685004 6221
rect -1076 6141 685004 6165
rect -1076 6085 -1064 6141
rect -1008 6085 -984 6141
rect -928 6085 -904 6141
rect -848 6085 -824 6141
rect -768 6085 86831 6141
rect 86887 6085 86911 6141
rect 86967 6085 86991 6141
rect 87047 6085 87071 6141
rect 87127 6085 257261 6141
rect 257317 6085 257341 6141
rect 257397 6085 257421 6141
rect 257477 6085 257501 6141
rect 257557 6085 427691 6141
rect 427747 6085 427771 6141
rect 427827 6085 427851 6141
rect 427907 6085 427931 6141
rect 427987 6085 598121 6141
rect 598177 6085 598201 6141
rect 598257 6085 598281 6141
rect 598337 6085 598361 6141
rect 598417 6085 684696 6141
rect 684752 6085 684776 6141
rect 684832 6085 684856 6141
rect 684912 6085 684936 6141
rect 684992 6085 685004 6141
rect -1076 6073 685004 6085
rect -1076 5721 685004 5733
rect -1076 5665 -404 5721
rect -348 5665 -324 5721
rect -268 5665 -244 5721
rect -188 5665 -164 5721
rect -108 5665 86171 5721
rect 86227 5665 86251 5721
rect 86307 5665 86331 5721
rect 86387 5665 86411 5721
rect 86467 5665 256601 5721
rect 256657 5665 256681 5721
rect 256737 5665 256761 5721
rect 256817 5665 256841 5721
rect 256897 5665 427031 5721
rect 427087 5665 427111 5721
rect 427167 5665 427191 5721
rect 427247 5665 427271 5721
rect 427327 5665 597461 5721
rect 597517 5665 597541 5721
rect 597597 5665 597621 5721
rect 597677 5665 597701 5721
rect 597757 5665 684036 5721
rect 684092 5665 684116 5721
rect 684172 5665 684196 5721
rect 684252 5665 684276 5721
rect 684332 5665 685004 5721
rect -1076 5641 685004 5665
rect -1076 5585 -404 5641
rect -348 5585 -324 5641
rect -268 5585 -244 5641
rect -188 5585 -164 5641
rect -108 5585 86171 5641
rect 86227 5585 86251 5641
rect 86307 5585 86331 5641
rect 86387 5585 86411 5641
rect 86467 5585 256601 5641
rect 256657 5585 256681 5641
rect 256737 5585 256761 5641
rect 256817 5585 256841 5641
rect 256897 5585 427031 5641
rect 427087 5585 427111 5641
rect 427167 5585 427191 5641
rect 427247 5585 427271 5641
rect 427327 5585 597461 5641
rect 597517 5585 597541 5641
rect 597597 5585 597621 5641
rect 597677 5585 597701 5641
rect 597757 5585 684036 5641
rect 684092 5585 684116 5641
rect 684172 5585 684196 5641
rect 684252 5585 684276 5641
rect 684332 5585 685004 5641
rect -1076 5561 685004 5585
rect -1076 5505 -404 5561
rect -348 5505 -324 5561
rect -268 5505 -244 5561
rect -188 5505 -164 5561
rect -108 5505 86171 5561
rect 86227 5505 86251 5561
rect 86307 5505 86331 5561
rect 86387 5505 86411 5561
rect 86467 5505 256601 5561
rect 256657 5505 256681 5561
rect 256737 5505 256761 5561
rect 256817 5505 256841 5561
rect 256897 5505 427031 5561
rect 427087 5505 427111 5561
rect 427167 5505 427191 5561
rect 427247 5505 427271 5561
rect 427327 5505 597461 5561
rect 597517 5505 597541 5561
rect 597597 5505 597621 5561
rect 597677 5505 597701 5561
rect 597757 5505 684036 5561
rect 684092 5505 684116 5561
rect 684172 5505 684196 5561
rect 684252 5505 684276 5561
rect 684332 5505 685004 5561
rect -1076 5481 685004 5505
rect -1076 5425 -404 5481
rect -348 5425 -324 5481
rect -268 5425 -244 5481
rect -188 5425 -164 5481
rect -108 5425 86171 5481
rect 86227 5425 86251 5481
rect 86307 5425 86331 5481
rect 86387 5425 86411 5481
rect 86467 5425 256601 5481
rect 256657 5425 256681 5481
rect 256737 5425 256761 5481
rect 256817 5425 256841 5481
rect 256897 5425 427031 5481
rect 427087 5425 427111 5481
rect 427167 5425 427191 5481
rect 427247 5425 427271 5481
rect 427327 5425 597461 5481
rect 597517 5425 597541 5481
rect 597597 5425 597621 5481
rect 597677 5425 597701 5481
rect 597757 5425 684036 5481
rect 684092 5425 684116 5481
rect 684172 5425 684196 5481
rect 684252 5425 684276 5481
rect 684332 5425 685004 5481
rect -1076 5413 685004 5425
rect -1076 5022 685004 5034
rect -1076 4966 -1064 5022
rect -1008 4966 -984 5022
rect -928 4966 -904 5022
rect -848 4966 -824 5022
rect -768 4966 86831 5022
rect 86887 4966 86911 5022
rect 86967 4966 86991 5022
rect 87047 4966 87071 5022
rect 87127 4966 257261 5022
rect 257317 4966 257341 5022
rect 257397 4966 257421 5022
rect 257477 4966 257501 5022
rect 257557 4966 427691 5022
rect 427747 4966 427771 5022
rect 427827 4966 427851 5022
rect 427907 4966 427931 5022
rect 427987 4966 598121 5022
rect 598177 4966 598201 5022
rect 598257 4966 598281 5022
rect 598337 4966 598361 5022
rect 598417 4966 684696 5022
rect 684752 4966 684776 5022
rect 684832 4966 684856 5022
rect 684912 4966 684936 5022
rect 684992 4966 685004 5022
rect -1076 4942 685004 4966
rect -1076 4886 -1064 4942
rect -1008 4886 -984 4942
rect -928 4886 -904 4942
rect -848 4886 -824 4942
rect -768 4886 86831 4942
rect 86887 4886 86911 4942
rect 86967 4886 86991 4942
rect 87047 4886 87071 4942
rect 87127 4886 257261 4942
rect 257317 4886 257341 4942
rect 257397 4886 257421 4942
rect 257477 4886 257501 4942
rect 257557 4886 427691 4942
rect 427747 4886 427771 4942
rect 427827 4886 427851 4942
rect 427907 4886 427931 4942
rect 427987 4886 598121 4942
rect 598177 4886 598201 4942
rect 598257 4886 598281 4942
rect 598337 4886 598361 4942
rect 598417 4886 684696 4942
rect 684752 4886 684776 4942
rect 684832 4886 684856 4942
rect 684912 4886 684936 4942
rect 684992 4886 685004 4942
rect -1076 4862 685004 4886
rect -1076 4806 -1064 4862
rect -1008 4806 -984 4862
rect -928 4806 -904 4862
rect -848 4806 -824 4862
rect -768 4806 86831 4862
rect 86887 4806 86911 4862
rect 86967 4806 86991 4862
rect 87047 4806 87071 4862
rect 87127 4806 257261 4862
rect 257317 4806 257341 4862
rect 257397 4806 257421 4862
rect 257477 4806 257501 4862
rect 257557 4806 427691 4862
rect 427747 4806 427771 4862
rect 427827 4806 427851 4862
rect 427907 4806 427931 4862
rect 427987 4806 598121 4862
rect 598177 4806 598201 4862
rect 598257 4806 598281 4862
rect 598337 4806 598361 4862
rect 598417 4806 684696 4862
rect 684752 4806 684776 4862
rect 684832 4806 684856 4862
rect 684912 4806 684936 4862
rect 684992 4806 685004 4862
rect -1076 4782 685004 4806
rect -1076 4726 -1064 4782
rect -1008 4726 -984 4782
rect -928 4726 -904 4782
rect -848 4726 -824 4782
rect -768 4726 86831 4782
rect 86887 4726 86911 4782
rect 86967 4726 86991 4782
rect 87047 4726 87071 4782
rect 87127 4726 257261 4782
rect 257317 4726 257341 4782
rect 257397 4726 257421 4782
rect 257477 4726 257501 4782
rect 257557 4726 427691 4782
rect 427747 4726 427771 4782
rect 427827 4726 427851 4782
rect 427907 4726 427931 4782
rect 427987 4726 598121 4782
rect 598177 4726 598201 4782
rect 598257 4726 598281 4782
rect 598337 4726 598361 4782
rect 598417 4726 684696 4782
rect 684752 4726 684776 4782
rect 684832 4726 684856 4782
rect 684912 4726 684936 4782
rect 684992 4726 685004 4782
rect -1076 4714 685004 4726
rect -1076 4362 685004 4374
rect -1076 4306 -404 4362
rect -348 4306 -324 4362
rect -268 4306 -244 4362
rect -188 4306 -164 4362
rect -108 4306 86171 4362
rect 86227 4306 86251 4362
rect 86307 4306 86331 4362
rect 86387 4306 86411 4362
rect 86467 4306 256601 4362
rect 256657 4306 256681 4362
rect 256737 4306 256761 4362
rect 256817 4306 256841 4362
rect 256897 4306 427031 4362
rect 427087 4306 427111 4362
rect 427167 4306 427191 4362
rect 427247 4306 427271 4362
rect 427327 4306 597461 4362
rect 597517 4306 597541 4362
rect 597597 4306 597621 4362
rect 597677 4306 597701 4362
rect 597757 4306 684036 4362
rect 684092 4306 684116 4362
rect 684172 4306 684196 4362
rect 684252 4306 684276 4362
rect 684332 4306 685004 4362
rect -1076 4282 685004 4306
rect -1076 4226 -404 4282
rect -348 4226 -324 4282
rect -268 4226 -244 4282
rect -188 4226 -164 4282
rect -108 4226 86171 4282
rect 86227 4226 86251 4282
rect 86307 4226 86331 4282
rect 86387 4226 86411 4282
rect 86467 4226 256601 4282
rect 256657 4226 256681 4282
rect 256737 4226 256761 4282
rect 256817 4226 256841 4282
rect 256897 4226 427031 4282
rect 427087 4226 427111 4282
rect 427167 4226 427191 4282
rect 427247 4226 427271 4282
rect 427327 4226 597461 4282
rect 597517 4226 597541 4282
rect 597597 4226 597621 4282
rect 597677 4226 597701 4282
rect 597757 4226 684036 4282
rect 684092 4226 684116 4282
rect 684172 4226 684196 4282
rect 684252 4226 684276 4282
rect 684332 4226 685004 4282
rect -1076 4202 685004 4226
rect -1076 4146 -404 4202
rect -348 4146 -324 4202
rect -268 4146 -244 4202
rect -188 4146 -164 4202
rect -108 4146 86171 4202
rect 86227 4146 86251 4202
rect 86307 4146 86331 4202
rect 86387 4146 86411 4202
rect 86467 4146 256601 4202
rect 256657 4146 256681 4202
rect 256737 4146 256761 4202
rect 256817 4146 256841 4202
rect 256897 4146 427031 4202
rect 427087 4146 427111 4202
rect 427167 4146 427191 4202
rect 427247 4146 427271 4202
rect 427327 4146 597461 4202
rect 597517 4146 597541 4202
rect 597597 4146 597621 4202
rect 597677 4146 597701 4202
rect 597757 4146 684036 4202
rect 684092 4146 684116 4202
rect 684172 4146 684196 4202
rect 684252 4146 684276 4202
rect 684332 4146 685004 4202
rect -1076 4122 685004 4146
rect -1076 4066 -404 4122
rect -348 4066 -324 4122
rect -268 4066 -244 4122
rect -188 4066 -164 4122
rect -108 4066 86171 4122
rect 86227 4066 86251 4122
rect 86307 4066 86331 4122
rect 86387 4066 86411 4122
rect 86467 4066 256601 4122
rect 256657 4066 256681 4122
rect 256737 4066 256761 4122
rect 256817 4066 256841 4122
rect 256897 4066 427031 4122
rect 427087 4066 427111 4122
rect 427167 4066 427191 4122
rect 427247 4066 427271 4122
rect 427327 4066 597461 4122
rect 597517 4066 597541 4122
rect 597597 4066 597621 4122
rect 597677 4066 597701 4122
rect 597757 4066 684036 4122
rect 684092 4066 684116 4122
rect 684172 4066 684196 4122
rect 684252 4066 684276 4122
rect 684332 4066 685004 4122
rect -1076 4054 685004 4066
rect -1076 3663 685004 3675
rect -1076 3607 -1064 3663
rect -1008 3607 -984 3663
rect -928 3607 -904 3663
rect -848 3607 -824 3663
rect -768 3607 86831 3663
rect 86887 3607 86911 3663
rect 86967 3607 86991 3663
rect 87047 3607 87071 3663
rect 87127 3607 257261 3663
rect 257317 3607 257341 3663
rect 257397 3607 257421 3663
rect 257477 3607 257501 3663
rect 257557 3607 427691 3663
rect 427747 3607 427771 3663
rect 427827 3607 427851 3663
rect 427907 3607 427931 3663
rect 427987 3607 598121 3663
rect 598177 3607 598201 3663
rect 598257 3607 598281 3663
rect 598337 3607 598361 3663
rect 598417 3607 684696 3663
rect 684752 3607 684776 3663
rect 684832 3607 684856 3663
rect 684912 3607 684936 3663
rect 684992 3607 685004 3663
rect -1076 3583 685004 3607
rect -1076 3527 -1064 3583
rect -1008 3527 -984 3583
rect -928 3527 -904 3583
rect -848 3527 -824 3583
rect -768 3527 86831 3583
rect 86887 3527 86911 3583
rect 86967 3527 86991 3583
rect 87047 3527 87071 3583
rect 87127 3527 257261 3583
rect 257317 3527 257341 3583
rect 257397 3527 257421 3583
rect 257477 3527 257501 3583
rect 257557 3527 427691 3583
rect 427747 3527 427771 3583
rect 427827 3527 427851 3583
rect 427907 3527 427931 3583
rect 427987 3527 598121 3583
rect 598177 3527 598201 3583
rect 598257 3527 598281 3583
rect 598337 3527 598361 3583
rect 598417 3527 684696 3583
rect 684752 3527 684776 3583
rect 684832 3527 684856 3583
rect 684912 3527 684936 3583
rect 684992 3527 685004 3583
rect -1076 3503 685004 3527
rect -1076 3447 -1064 3503
rect -1008 3447 -984 3503
rect -928 3447 -904 3503
rect -848 3447 -824 3503
rect -768 3447 86831 3503
rect 86887 3447 86911 3503
rect 86967 3447 86991 3503
rect 87047 3447 87071 3503
rect 87127 3447 257261 3503
rect 257317 3447 257341 3503
rect 257397 3447 257421 3503
rect 257477 3447 257501 3503
rect 257557 3447 427691 3503
rect 427747 3447 427771 3503
rect 427827 3447 427851 3503
rect 427907 3447 427931 3503
rect 427987 3447 598121 3503
rect 598177 3447 598201 3503
rect 598257 3447 598281 3503
rect 598337 3447 598361 3503
rect 598417 3447 684696 3503
rect 684752 3447 684776 3503
rect 684832 3447 684856 3503
rect 684912 3447 684936 3503
rect 684992 3447 685004 3503
rect -1076 3423 685004 3447
rect -1076 3367 -1064 3423
rect -1008 3367 -984 3423
rect -928 3367 -904 3423
rect -848 3367 -824 3423
rect -768 3367 86831 3423
rect 86887 3367 86911 3423
rect 86967 3367 86991 3423
rect 87047 3367 87071 3423
rect 87127 3367 257261 3423
rect 257317 3367 257341 3423
rect 257397 3367 257421 3423
rect 257477 3367 257501 3423
rect 257557 3367 427691 3423
rect 427747 3367 427771 3423
rect 427827 3367 427851 3423
rect 427907 3367 427931 3423
rect 427987 3367 598121 3423
rect 598177 3367 598201 3423
rect 598257 3367 598281 3423
rect 598337 3367 598361 3423
rect 598417 3367 684696 3423
rect 684752 3367 684776 3423
rect 684832 3367 684856 3423
rect 684912 3367 684936 3423
rect 684992 3367 685004 3423
rect -1076 3355 685004 3367
rect -1076 3003 685004 3015
rect -1076 2947 -404 3003
rect -348 2947 -324 3003
rect -268 2947 -244 3003
rect -188 2947 -164 3003
rect -108 2947 86171 3003
rect 86227 2947 86251 3003
rect 86307 2947 86331 3003
rect 86387 2947 86411 3003
rect 86467 2947 256601 3003
rect 256657 2947 256681 3003
rect 256737 2947 256761 3003
rect 256817 2947 256841 3003
rect 256897 2947 427031 3003
rect 427087 2947 427111 3003
rect 427167 2947 427191 3003
rect 427247 2947 427271 3003
rect 427327 2947 597461 3003
rect 597517 2947 597541 3003
rect 597597 2947 597621 3003
rect 597677 2947 597701 3003
rect 597757 2947 684036 3003
rect 684092 2947 684116 3003
rect 684172 2947 684196 3003
rect 684252 2947 684276 3003
rect 684332 2947 685004 3003
rect -1076 2923 685004 2947
rect -1076 2867 -404 2923
rect -348 2867 -324 2923
rect -268 2867 -244 2923
rect -188 2867 -164 2923
rect -108 2867 86171 2923
rect 86227 2867 86251 2923
rect 86307 2867 86331 2923
rect 86387 2867 86411 2923
rect 86467 2867 256601 2923
rect 256657 2867 256681 2923
rect 256737 2867 256761 2923
rect 256817 2867 256841 2923
rect 256897 2867 427031 2923
rect 427087 2867 427111 2923
rect 427167 2867 427191 2923
rect 427247 2867 427271 2923
rect 427327 2867 597461 2923
rect 597517 2867 597541 2923
rect 597597 2867 597621 2923
rect 597677 2867 597701 2923
rect 597757 2867 684036 2923
rect 684092 2867 684116 2923
rect 684172 2867 684196 2923
rect 684252 2867 684276 2923
rect 684332 2867 685004 2923
rect -1076 2843 685004 2867
rect -1076 2787 -404 2843
rect -348 2787 -324 2843
rect -268 2787 -244 2843
rect -188 2787 -164 2843
rect -108 2787 86171 2843
rect 86227 2787 86251 2843
rect 86307 2787 86331 2843
rect 86387 2787 86411 2843
rect 86467 2787 256601 2843
rect 256657 2787 256681 2843
rect 256737 2787 256761 2843
rect 256817 2787 256841 2843
rect 256897 2787 427031 2843
rect 427087 2787 427111 2843
rect 427167 2787 427191 2843
rect 427247 2787 427271 2843
rect 427327 2787 597461 2843
rect 597517 2787 597541 2843
rect 597597 2787 597621 2843
rect 597677 2787 597701 2843
rect 597757 2787 684036 2843
rect 684092 2787 684116 2843
rect 684172 2787 684196 2843
rect 684252 2787 684276 2843
rect 684332 2787 685004 2843
rect -1076 2763 685004 2787
rect -1076 2707 -404 2763
rect -348 2707 -324 2763
rect -268 2707 -244 2763
rect -188 2707 -164 2763
rect -108 2707 86171 2763
rect 86227 2707 86251 2763
rect 86307 2707 86331 2763
rect 86387 2707 86411 2763
rect 86467 2707 256601 2763
rect 256657 2707 256681 2763
rect 256737 2707 256761 2763
rect 256817 2707 256841 2763
rect 256897 2707 427031 2763
rect 427087 2707 427111 2763
rect 427167 2707 427191 2763
rect 427247 2707 427271 2763
rect 427327 2707 597461 2763
rect 597517 2707 597541 2763
rect 597597 2707 597621 2763
rect 597677 2707 597701 2763
rect 597757 2707 684036 2763
rect 684092 2707 684116 2763
rect 684172 2707 684196 2763
rect 684252 2707 684276 2763
rect 684332 2707 685004 2763
rect -1076 2695 685004 2707
rect 236821 2546 236887 2549
rect 326153 2546 326219 2549
rect 236821 2544 326219 2546
rect 236821 2488 236826 2544
rect 236882 2488 326158 2544
rect 326214 2488 326219 2544
rect 236821 2486 326219 2488
rect 236821 2483 236887 2486
rect 326153 2483 326219 2486
rect 431861 2546 431927 2549
rect 525057 2546 525123 2549
rect 431861 2544 525123 2546
rect 431861 2488 431866 2544
rect 431922 2488 525062 2544
rect 525118 2488 525123 2544
rect 431861 2486 525123 2488
rect 431861 2483 431927 2486
rect 525057 2483 525123 2486
rect 337009 2410 337075 2413
rect 430757 2410 430823 2413
rect 337009 2408 430823 2410
rect 337009 2352 337014 2408
rect 337070 2352 430762 2408
rect 430818 2352 430823 2408
rect 337009 2350 430823 2352
rect 337009 2347 337075 2350
rect 430757 2347 430823 2350
rect 242065 1730 242131 1733
rect 249425 1730 249491 1733
rect 242065 1728 249491 1730
rect 242065 1672 242070 1728
rect 242126 1672 249430 1728
rect 249486 1672 249491 1728
rect 242065 1670 249491 1672
rect 242065 1667 242131 1670
rect 249425 1667 249491 1670
rect 241789 1594 241855 1597
rect 244825 1594 244891 1597
rect 241789 1592 244891 1594
rect 241789 1536 241794 1592
rect 241850 1536 244830 1592
rect 244886 1536 244891 1592
rect 241789 1534 244891 1536
rect 241789 1531 241855 1534
rect 244825 1531 244891 1534
rect 239949 1458 240015 1461
rect 243997 1458 244063 1461
rect 239949 1456 244063 1458
rect 239949 1400 239954 1456
rect 240010 1400 244002 1456
rect 244058 1400 244063 1456
rect 239949 1398 244063 1400
rect 239949 1395 240015 1398
rect 243997 1395 244063 1398
rect 244273 1458 244339 1461
rect 248413 1458 248479 1461
rect 244273 1456 248479 1458
rect 244273 1400 244278 1456
rect 244334 1400 248418 1456
rect 248474 1400 248479 1456
rect 244273 1398 248479 1400
rect 244273 1395 244339 1398
rect 248413 1395 248479 1398
rect 244549 1322 244615 1325
rect 246389 1322 246455 1325
rect 244549 1320 246455 1322
rect 244549 1264 244554 1320
rect 244610 1264 246394 1320
rect 246450 1264 246455 1320
rect 244549 1262 246455 1264
rect 244549 1259 244615 1262
rect 246389 1259 246455 1262
rect 227437 1186 227503 1189
rect 229461 1186 229527 1189
rect 227437 1184 229527 1186
rect 227437 1128 227442 1184
rect 227498 1128 229466 1184
rect 229522 1128 229527 1184
rect 227437 1126 229527 1128
rect 227437 1123 227503 1126
rect 229461 1123 229527 1126
rect 243997 1186 244063 1189
rect 244641 1186 244707 1189
rect 243997 1184 244707 1186
rect 243997 1128 244002 1184
rect 244058 1128 244646 1184
rect 244702 1128 244707 1184
rect 243997 1126 244707 1128
rect 243997 1123 244063 1126
rect 244641 1123 244707 1126
rect -416 964 684344 976
rect -416 908 -404 964
rect -348 908 -324 964
rect -268 908 -244 964
rect -188 908 -164 964
rect -108 908 86171 964
rect 86227 908 86251 964
rect 86307 908 86331 964
rect 86387 908 86411 964
rect 86467 908 256601 964
rect 256657 908 256681 964
rect 256737 908 256761 964
rect 256817 908 256841 964
rect 256897 908 427031 964
rect 427087 908 427111 964
rect 427167 908 427191 964
rect 427247 908 427271 964
rect 427327 908 597461 964
rect 597517 908 597541 964
rect 597597 908 597621 964
rect 597677 908 597701 964
rect 597757 908 684036 964
rect 684092 908 684116 964
rect 684172 908 684196 964
rect 684252 908 684276 964
rect 684332 908 684344 964
rect -416 884 684344 908
rect -416 828 -404 884
rect -348 828 -324 884
rect -268 828 -244 884
rect -188 828 -164 884
rect -108 828 86171 884
rect 86227 828 86251 884
rect 86307 828 86331 884
rect 86387 828 86411 884
rect 86467 828 256601 884
rect 256657 828 256681 884
rect 256737 828 256761 884
rect 256817 828 256841 884
rect 256897 828 427031 884
rect 427087 828 427111 884
rect 427167 828 427191 884
rect 427247 828 427271 884
rect 427327 828 597461 884
rect 597517 828 597541 884
rect 597597 828 597621 884
rect 597677 828 597701 884
rect 597757 828 684036 884
rect 684092 828 684116 884
rect 684172 828 684196 884
rect 684252 828 684276 884
rect 684332 828 684344 884
rect -416 804 684344 828
rect -416 748 -404 804
rect -348 748 -324 804
rect -268 748 -244 804
rect -188 748 -164 804
rect -108 748 86171 804
rect 86227 748 86251 804
rect 86307 748 86331 804
rect 86387 748 86411 804
rect 86467 748 256601 804
rect 256657 748 256681 804
rect 256737 748 256761 804
rect 256817 748 256841 804
rect 256897 748 427031 804
rect 427087 748 427111 804
rect 427167 748 427191 804
rect 427247 748 427271 804
rect 427327 748 597461 804
rect 597517 748 597541 804
rect 597597 748 597621 804
rect 597677 748 597701 804
rect 597757 748 684036 804
rect 684092 748 684116 804
rect 684172 748 684196 804
rect 684252 748 684276 804
rect 684332 748 684344 804
rect -416 724 684344 748
rect -416 668 -404 724
rect -348 668 -324 724
rect -268 668 -244 724
rect -188 668 -164 724
rect -108 668 86171 724
rect 86227 668 86251 724
rect 86307 668 86331 724
rect 86387 668 86411 724
rect 86467 668 256601 724
rect 256657 668 256681 724
rect 256737 668 256761 724
rect 256817 668 256841 724
rect 256897 668 427031 724
rect 427087 668 427111 724
rect 427167 668 427191 724
rect 427247 668 427271 724
rect 427327 668 597461 724
rect 597517 668 597541 724
rect 597597 668 597621 724
rect 597677 668 597701 724
rect 597757 668 684036 724
rect 684092 668 684116 724
rect 684172 668 684196 724
rect 684252 668 684276 724
rect 684332 668 684344 724
rect -416 656 684344 668
rect 243629 506 243695 509
rect 244457 506 244523 509
rect 243629 504 244523 506
rect 243629 448 243634 504
rect 243690 448 244462 504
rect 244518 448 244523 504
rect 243629 446 244523 448
rect 243629 443 243695 446
rect 244457 443 244523 446
rect -1076 304 685004 316
rect -1076 248 -1064 304
rect -1008 248 -984 304
rect -928 248 -904 304
rect -848 248 -824 304
rect -768 248 86831 304
rect 86887 248 86911 304
rect 86967 248 86991 304
rect 87047 248 87071 304
rect 87127 248 257261 304
rect 257317 248 257341 304
rect 257397 248 257421 304
rect 257477 248 257501 304
rect 257557 248 427691 304
rect 427747 248 427771 304
rect 427827 248 427851 304
rect 427907 248 427931 304
rect 427987 248 598121 304
rect 598177 248 598201 304
rect 598257 248 598281 304
rect 598337 248 598361 304
rect 598417 248 684696 304
rect 684752 248 684776 304
rect 684832 248 684856 304
rect 684912 248 684936 304
rect 684992 248 685004 304
rect -1076 224 685004 248
rect -1076 168 -1064 224
rect -1008 168 -984 224
rect -928 168 -904 224
rect -848 168 -824 224
rect -768 168 86831 224
rect 86887 168 86911 224
rect 86967 168 86991 224
rect 87047 168 87071 224
rect 87127 168 257261 224
rect 257317 168 257341 224
rect 257397 168 257421 224
rect 257477 168 257501 224
rect 257557 168 427691 224
rect 427747 168 427771 224
rect 427827 168 427851 224
rect 427907 168 427931 224
rect 427987 168 598121 224
rect 598177 168 598201 224
rect 598257 168 598281 224
rect 598337 168 598361 224
rect 598417 168 684696 224
rect 684752 168 684776 224
rect 684832 168 684856 224
rect 684912 168 684936 224
rect 684992 168 685004 224
rect -1076 144 685004 168
rect -1076 88 -1064 144
rect -1008 88 -984 144
rect -928 88 -904 144
rect -848 88 -824 144
rect -768 88 86831 144
rect 86887 88 86911 144
rect 86967 88 86991 144
rect 87047 88 87071 144
rect 87127 88 257261 144
rect 257317 88 257341 144
rect 257397 88 257421 144
rect 257477 88 257501 144
rect 257557 88 427691 144
rect 427747 88 427771 144
rect 427827 88 427851 144
rect 427907 88 427931 144
rect 427987 88 598121 144
rect 598177 88 598201 144
rect 598257 88 598281 144
rect 598337 88 598361 144
rect 598417 88 684696 144
rect 684752 88 684776 144
rect 684832 88 684856 144
rect 684912 88 684936 144
rect 684992 88 685004 144
rect -1076 64 685004 88
rect -1076 8 -1064 64
rect -1008 8 -984 64
rect -928 8 -904 64
rect -848 8 -824 64
rect -768 8 86831 64
rect 86887 8 86911 64
rect 86967 8 86991 64
rect 87047 8 87071 64
rect 87127 8 257261 64
rect 257317 8 257341 64
rect 257397 8 257421 64
rect 257477 8 257501 64
rect 257557 8 427691 64
rect 427747 8 427771 64
rect 427827 8 427851 64
rect 427907 8 427931 64
rect 427987 8 598121 64
rect 598177 8 598201 64
rect 598257 8 598281 64
rect 598337 8 598361 64
rect 598417 8 684696 64
rect 684752 8 684776 64
rect 684832 8 684856 64
rect 684912 8 684936 64
rect 684992 8 685004 64
rect -1076 -4 685004 8
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[0\].u_buf_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[1\].u_buf_A
timestamp 1676037725
transform -1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[2\].u_buf_A
timestamp 1676037725
transform -1 0 33580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[3\].u_buf_A
timestamp 1676037725
transform -1 0 49036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[4\].u_buf_A
timestamp 1676037725
transform -1 0 64492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[5\].u_buf_A
timestamp 1676037725
transform 1 0 78844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[6\].u_buf_A
timestamp 1676037725
transform -1 0 95404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[7\].u_buf_A
timestamp 1676037725
transform -1 0 110860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[8\].u_buf_A
timestamp 1676037725
transform -1 0 126316 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[9\].u_buf_A
timestamp 1676037725
transform -1 0 141772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[10\].u_buf_A
timestamp 1676037725
transform -1 0 157228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[11\].u_buf_A
timestamp 1676037725
transform 1 0 171580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[12\].u_buf_A
timestamp 1676037725
transform -1 0 187772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[13\].u_buf_A
timestamp 1676037725
transform -1 0 203228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[14\].u_buf_A
timestamp 1676037725
transform 1 0 217948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[15\].u_buf_A
timestamp 1676037725
transform -1 0 234508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[16\].u_buf_A
timestamp 1676037725
transform -1 0 248216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[17\].u_buf_A
timestamp 1676037725
transform 1 0 264316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[18\].u_buf_A
timestamp 1676037725
transform -1 0 279128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[19\].u_buf_A
timestamp 1676037725
transform -1 0 294584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[20\].u_buf_A
timestamp 1676037725
transform 1 0 310684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[21\].u_buf_A
timestamp 1676037725
transform -1 0 326324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[22\].u_buf_A
timestamp 1676037725
transform -1 0 342700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[23\].u_buf_A
timestamp 1676037725
transform 1 0 357052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[24\].u_buf_A
timestamp 1676037725
transform 1 0 372508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[25\].u_buf_A
timestamp 1676037725
transform 1 0 387964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[26\].u_buf_A
timestamp 1676037725
transform 1 0 403420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[27\].u_buf_A
timestamp 1676037725
transform -1 0 419060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[28\].u_buf_A
timestamp 1676037725
transform -1 0 434516 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[29\].u_buf_A
timestamp 1676037725
transform 1 0 449788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[30\].u_buf_A
timestamp 1676037725
transform -1 0 465428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[31\].u_buf_A
timestamp 1676037725
transform -1 0 480884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[32\].u_buf_A
timestamp 1676037725
transform 1 0 496156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[33\].u_buf_A
timestamp 1676037725
transform -1 0 511796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[34\].u_buf_A
timestamp 1676037725
transform -1 0 527252 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[35\].u_buf_A
timestamp 1676037725
transform -1 0 543628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[36\].u_buf_A
timestamp 1676037725
transform 1 0 557980 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[37\].u_buf_A
timestamp 1676037725
transform 1 0 573436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[38\].u_buf_A
timestamp 1676037725
transform 1 0 588892 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[39\].u_buf_A
timestamp 1676037725
transform -1 0 604532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[40\].u_buf_A
timestamp 1676037725
transform -1 0 619988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[41\].u_buf_A
timestamp 1676037725
transform -1 0 636364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[42\].u_buf_A
timestamp 1676037725
transform -1 0 650900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[43\].u_buf_A
timestamp 1676037725
transform -1 0 666356 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[44\].u_buf_A
timestamp 1676037725
transform 1 0 681628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire2_A
timestamp 1676037725
transform -1 0 136528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire3_A
timestamp 1676037725
transform 1 0 342608 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire4_A
timestamp 1676037725
transform -1 0 436908 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire5_A
timestamp 1676037725
transform -1 0 531024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire6_A
timestamp 1676037725
transform -1 0 626152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire7_A
timestamp 1676037725
transform -1 0 339940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire8_A
timestamp 1676037725
transform 1 0 435344 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire9_A
timestamp 1676037725
transform -1 0 529184 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire11_A
timestamp 1676037725
transform -1 0 339020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire12_A
timestamp 1676037725
transform -1 0 433964 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire13_A
timestamp 1676037725
transform 1 0 528080 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire14_A
timestamp 1676037725
transform -1 0 337732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire15_A
timestamp 1676037725
transform -1 0 433412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire17_A
timestamp 1676037725
transform -1 0 335800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire18_A
timestamp 1676037725
transform -1 0 431020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire19_A
timestamp 1676037725
transform -1 0 134872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire21_A
timestamp 1676037725
transform -1 0 334972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire22_A
timestamp 1676037725
transform -1 0 429180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire23_A
timestamp 1676037725
transform -1 0 333408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire24_A
timestamp 1676037725
transform -1 0 331844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire25_A
timestamp 1676037725
transform -1 0 205068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire26_A
timestamp 1676037725
transform -1 0 189612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire27_A
timestamp 1676037725
transform -1 0 159896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire28_A
timestamp 1676037725
transform -1 0 570952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire29_A
timestamp 1676037725
transform -1 0 477480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire30_A
timestamp 1676037725
transform -1 0 382996 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire31_A
timestamp 1676037725
transform -1 0 288144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire32_A
timestamp 1676037725
transform -1 0 555496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire33_A
timestamp 1676037725
transform -1 0 462024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire34_A
timestamp 1676037725
transform -1 0 367632 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire35_A
timestamp 1676037725
transform -1 0 272688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire36_A
timestamp 1676037725
transform 1 0 525044 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire37_A
timestamp 1676037725
transform 1 0 430744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire38_A
timestamp 1676037725
transform -1 0 336352 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire39_A
timestamp 1676037725
transform -1 0 144440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire40_A
timestamp 1676037725
transform -1 0 509772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire41_A
timestamp 1676037725
transform -1 0 415656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire42_A
timestamp 1676037725
transform -1 0 321080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire43_A
timestamp 1676037725
transform 1 0 478676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire44_A
timestamp 1676037725
transform -1 0 384744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire45_A
timestamp 1676037725
transform -1 0 290260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire46_A
timestamp 1676037725
transform 1 0 463220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire47_A
timestamp 1676037725
transform -1 0 369288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire48_A
timestamp 1676037725
transform -1 0 274896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire49_A
timestamp 1676037725
transform -1 0 432860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire50_A
timestamp 1676037725
transform 1 0 338376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire51_A
timestamp 1676037725
transform -1 0 417404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire52_A
timestamp 1676037725
transform -1 0 323472 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire53_A
timestamp 1676037725
transform -1 0 386492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire54_A
timestamp 1676037725
transform -1 0 292744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire55_A
timestamp 1676037725
transform -1 0 371036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire56_A
timestamp 1676037725
transform -1 0 277380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire57_A
timestamp 1676037725
transform -1 0 340308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire58_A
timestamp 1676037725
transform -1 0 246376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire59_A
timestamp 1676037725
transform -1 0 324668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire60_A
timestamp 1676037725
transform 1 0 294400 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire61_A
timestamp 1676037725
transform 1 0 278944 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire62_A
timestamp 1676037725
transform -1 0 248860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire63_A
timestamp 1676037725
transform -1 0 113528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire64_A
timestamp 1676037725
transform -1 0 206816 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire65_A
timestamp 1676037725
transform -1 0 98072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire66_A
timestamp 1676037725
transform -1 0 191452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1676037725
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_185
timestamp 1676037725
transform 1 0 18124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_343 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1676037725
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 1676037725
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1676037725
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_429 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_437
timestamp 1676037725
transform 1 0 41308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1676037725
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1676037725
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1676037725
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_521
timestamp 1676037725
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1676037725
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1676037725
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1676037725
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1676037725
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1676037725
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1676037725
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1676037725
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1676037725
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1676037725
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1676037725
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1676037725
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1676037725
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1676037725
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1676037725
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_673
timestamp 1676037725
transform 1 0 63020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_683
timestamp 1676037725
transform 1 0 63940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_689
timestamp 1676037725
transform 1 0 64492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1676037725
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1676037725
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1676037725
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1676037725
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1676037725
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1676037725
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1676037725
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1676037725
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1676037725
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1676037725
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1676037725
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1676037725
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1676037725
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1676037725
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1676037725
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1676037725
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_841
timestamp 1676037725
transform 1 0 78476 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_851
timestamp 1676037725
transform 1 0 79396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_863
timestamp 1676037725
transform 1 0 80500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_867
timestamp 1676037725
transform 1 0 80868 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1676037725
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1676037725
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1676037725
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1676037725
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1676037725
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1676037725
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1676037725
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1676037725
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1676037725
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1676037725
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1676037725
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1676037725
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1676037725
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1676037725
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1676037725
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1009
timestamp 1676037725
transform 1 0 93932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1019
timestamp 1676037725
transform 1 0 94852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1025
timestamp 1676037725
transform 1 0 95404 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1676037725
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1037
timestamp 1676037725
transform 1 0 96508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1048
timestamp 1676037725
transform 1 0 97520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1054
timestamp 1676037725
transform 1 0 98072 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1062
timestamp 1676037725
transform 1 0 98808 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1676037725
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1676037725
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1676037725
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1676037725
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1676037725
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1676037725
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1676037725
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1676037725
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1676037725
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1676037725
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1161
timestamp 1676037725
transform 1 0 107916 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1173
timestamp 1676037725
transform 1 0 109020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1177
timestamp 1676037725
transform 1 0 109388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1187
timestamp 1676037725
transform 1 0 110308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1193
timestamp 1676037725
transform 1 0 110860 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1201
timestamp 1676037725
transform 1 0 111596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1205
timestamp 1676037725
transform 1 0 111964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1216
timestamp 1676037725
transform 1 0 112976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1222
timestamp 1676037725
transform 1 0 113528 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1230
timestamp 1676037725
transform 1 0 114264 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1233
timestamp 1676037725
transform 1 0 114540 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1245
timestamp 1676037725
transform 1 0 115644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1257
timestamp 1676037725
transform 1 0 116748 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1261
timestamp 1676037725
transform 1 0 117116 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1273
timestamp 1676037725
transform 1 0 118220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1285
timestamp 1676037725
transform 1 0 119324 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1289
timestamp 1676037725
transform 1 0 119692 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1301
timestamp 1676037725
transform 1 0 120796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1313
timestamp 1676037725
transform 1 0 121900 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1317
timestamp 1676037725
transform 1 0 122268 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1329
timestamp 1676037725
transform 1 0 123372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1341
timestamp 1676037725
transform 1 0 124476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1345
timestamp 1676037725
transform 1 0 124844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1351
timestamp 1676037725
transform 1 0 125396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1355
timestamp 1676037725
transform 1 0 125764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1361
timestamp 1676037725
transform 1 0 126316 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1369
timestamp 1676037725
transform 1 0 127052 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1373
timestamp 1676037725
transform 1 0 127420 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1385
timestamp 1676037725
transform 1 0 128524 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1397
timestamp 1676037725
transform 1 0 129628 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1401
timestamp 1676037725
transform 1 0 129996 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1413
timestamp 1676037725
transform 1 0 131100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1425
timestamp 1676037725
transform 1 0 132204 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1429
timestamp 1676037725
transform 1 0 132572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1441
timestamp 1676037725
transform 1 0 133676 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1449
timestamp 1676037725
transform 1 0 134412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1454
timestamp 1676037725
transform 1 0 134872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1457
timestamp 1676037725
transform 1 0 135148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1468
timestamp 1676037725
transform 1 0 136160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1478
timestamp 1676037725
transform 1 0 137080 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1485
timestamp 1676037725
transform 1 0 137724 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1493
timestamp 1676037725
transform 1 0 138460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1505
timestamp 1676037725
transform 1 0 139564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1511
timestamp 1676037725
transform 1 0 140116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1513
timestamp 1676037725
transform 1 0 140300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1523
timestamp 1676037725
transform 1 0 141220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1529
timestamp 1676037725
transform 1 0 141772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1537
timestamp 1676037725
transform 1 0 142508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1541
timestamp 1676037725
transform 1 0 142876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1552
timestamp 1676037725
transform 1 0 143888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1558
timestamp 1676037725
transform 1 0 144440 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1566
timestamp 1676037725
transform 1 0 145176 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1569
timestamp 1676037725
transform 1 0 145452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1581
timestamp 1676037725
transform 1 0 146556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1593
timestamp 1676037725
transform 1 0 147660 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1597
timestamp 1676037725
transform 1 0 148028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1609
timestamp 1676037725
transform 1 0 149132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1621
timestamp 1676037725
transform 1 0 150236 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1625
timestamp 1676037725
transform 1 0 150604 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1637
timestamp 1676037725
transform 1 0 151708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1649
timestamp 1676037725
transform 1 0 152812 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1653
timestamp 1676037725
transform 1 0 153180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1665
timestamp 1676037725
transform 1 0 154284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1677
timestamp 1676037725
transform 1 0 155388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1681
timestamp 1676037725
transform 1 0 155756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1691
timestamp 1676037725
transform 1 0 156676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1697
timestamp 1676037725
transform 1 0 157228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1705
timestamp 1676037725
transform 1 0 157964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1709
timestamp 1676037725
transform 1 0 158332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1720
timestamp 1676037725
transform 1 0 159344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1726
timestamp 1676037725
transform 1 0 159896 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1734
timestamp 1676037725
transform 1 0 160632 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1737
timestamp 1676037725
transform 1 0 160908 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1749
timestamp 1676037725
transform 1 0 162012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1761
timestamp 1676037725
transform 1 0 163116 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1765
timestamp 1676037725
transform 1 0 163484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1777
timestamp 1676037725
transform 1 0 164588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1789
timestamp 1676037725
transform 1 0 165692 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1793
timestamp 1676037725
transform 1 0 166060 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1805
timestamp 1676037725
transform 1 0 167164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1817
timestamp 1676037725
transform 1 0 168268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1821
timestamp 1676037725
transform 1 0 168636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1833
timestamp 1676037725
transform 1 0 169740 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1845
timestamp 1676037725
transform 1 0 170844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1849
timestamp 1676037725
transform 1 0 171212 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1859
timestamp 1676037725
transform 1 0 172132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1871
timestamp 1676037725
transform 1 0 173236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1875
timestamp 1676037725
transform 1 0 173604 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1877
timestamp 1676037725
transform 1 0 173788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1889
timestamp 1676037725
transform 1 0 174892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1901
timestamp 1676037725
transform 1 0 175996 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1905
timestamp 1676037725
transform 1 0 176364 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1917
timestamp 1676037725
transform 1 0 177468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1929
timestamp 1676037725
transform 1 0 178572 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1933
timestamp 1676037725
transform 1 0 178940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1945
timestamp 1676037725
transform 1 0 180044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1957
timestamp 1676037725
transform 1 0 181148 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1961
timestamp 1676037725
transform 1 0 181516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1973
timestamp 1676037725
transform 1 0 182620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1985
timestamp 1676037725
transform 1 0 183724 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1989
timestamp 1676037725
transform 1 0 184092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2001
timestamp 1676037725
transform 1 0 185196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2013
timestamp 1676037725
transform 1 0 186300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2017
timestamp 1676037725
transform 1 0 186668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2027
timestamp 1676037725
transform 1 0 187588 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2035
timestamp 1676037725
transform 1 0 188324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2042
timestamp 1676037725
transform 1 0 188968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2045
timestamp 1676037725
transform 1 0 189244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2049
timestamp 1676037725
transform 1 0 189612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2063
timestamp 1676037725
transform 1 0 190900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2069
timestamp 1676037725
transform 1 0 191452 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2073
timestamp 1676037725
transform 1 0 191820 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2085
timestamp 1676037725
transform 1 0 192924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2097
timestamp 1676037725
transform 1 0 194028 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2101
timestamp 1676037725
transform 1 0 194396 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2113
timestamp 1676037725
transform 1 0 195500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2125
timestamp 1676037725
transform 1 0 196604 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2129
timestamp 1676037725
transform 1 0 196972 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2141
timestamp 1676037725
transform 1 0 198076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2153
timestamp 1676037725
transform 1 0 199180 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2157
timestamp 1676037725
transform 1 0 199548 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2169
timestamp 1676037725
transform 1 0 200652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2181
timestamp 1676037725
transform 1 0 201756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2185
timestamp 1676037725
transform 1 0 202124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2195
timestamp 1676037725
transform 1 0 203044 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2201
timestamp 1676037725
transform 1 0 203596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2208
timestamp 1676037725
transform 1 0 204240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2213
timestamp 1676037725
transform 1 0 204700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2217
timestamp 1676037725
transform 1 0 205068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2223
timestamp 1676037725
transform 1 0 205620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2230
timestamp 1676037725
transform 1 0 206264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2236
timestamp 1676037725
transform 1 0 206816 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2241
timestamp 1676037725
transform 1 0 207276 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2253
timestamp 1676037725
transform 1 0 208380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2265
timestamp 1676037725
transform 1 0 209484 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2269
timestamp 1676037725
transform 1 0 209852 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2281
timestamp 1676037725
transform 1 0 210956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2293
timestamp 1676037725
transform 1 0 212060 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2297
timestamp 1676037725
transform 1 0 212428 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2309
timestamp 1676037725
transform 1 0 213532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2321
timestamp 1676037725
transform 1 0 214636 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2325
timestamp 1676037725
transform 1 0 215004 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2337
timestamp 1676037725
transform 1 0 216108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2349
timestamp 1676037725
transform 1 0 217212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2353
timestamp 1676037725
transform 1 0 217580 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2363
timestamp 1676037725
transform 1 0 218500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2375
timestamp 1676037725
transform 1 0 219604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2379
timestamp 1676037725
transform 1 0 219972 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2381
timestamp 1676037725
transform 1 0 220156 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2393
timestamp 1676037725
transform 1 0 221260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2405
timestamp 1676037725
transform 1 0 222364 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2409
timestamp 1676037725
transform 1 0 222732 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2421
timestamp 1676037725
transform 1 0 223836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2433
timestamp 1676037725
transform 1 0 224940 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2437
timestamp 1676037725
transform 1 0 225308 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2449
timestamp 1676037725
transform 1 0 226412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2461
timestamp 1676037725
transform 1 0 227516 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2465
timestamp 1676037725
transform 1 0 227884 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2477
timestamp 1676037725
transform 1 0 228988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2489
timestamp 1676037725
transform 1 0 230092 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2493
timestamp 1676037725
transform 1 0 230460 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2505
timestamp 1676037725
transform 1 0 231564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2517
timestamp 1676037725
transform 1 0 232668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2521
timestamp 1676037725
transform 1 0 233036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2531
timestamp 1676037725
transform 1 0 233956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2537
timestamp 1676037725
transform 1 0 234508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2545
timestamp 1676037725
transform 1 0 235244 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2549
timestamp 1676037725
transform 1 0 235612 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2561
timestamp 1676037725
transform 1 0 236716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2573
timestamp 1676037725
transform 1 0 237820 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2577
timestamp 1676037725
transform 1 0 238188 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2589
timestamp 1676037725
transform 1 0 239292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2601
timestamp 1676037725
transform 1 0 240396 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2605
timestamp 1676037725
transform 1 0 240764 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2617
timestamp 1676037725
transform 1 0 241868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2629
timestamp 1676037725
transform 1 0 242972 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2633
timestamp 1676037725
transform 1 0 243340 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2645
timestamp 1676037725
transform 1 0 244444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2657
timestamp 1676037725
transform 1 0 245548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2661
timestamp 1676037725
transform 1 0 245916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2666
timestamp 1676037725
transform 1 0 246376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2676
timestamp 1676037725
transform 1 0 247296 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2686
timestamp 1676037725
transform 1 0 248216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2689
timestamp 1676037725
transform 1 0 248492 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2699
timestamp 1676037725
transform 1 0 249412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2711
timestamp 1676037725
transform 1 0 250516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2715
timestamp 1676037725
transform 1 0 250884 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2717
timestamp 1676037725
transform 1 0 251068 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2729
timestamp 1676037725
transform 1 0 252172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2741
timestamp 1676037725
transform 1 0 253276 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2745
timestamp 1676037725
transform 1 0 253644 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2757
timestamp 1676037725
transform 1 0 254748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2769
timestamp 1676037725
transform 1 0 255852 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2773
timestamp 1676037725
transform 1 0 256220 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2785
timestamp 1676037725
transform 1 0 257324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2797
timestamp 1676037725
transform 1 0 258428 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2801
timestamp 1676037725
transform 1 0 258796 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2813
timestamp 1676037725
transform 1 0 259900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2825
timestamp 1676037725
transform 1 0 261004 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2829
timestamp 1676037725
transform 1 0 261372 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2841
timestamp 1676037725
transform 1 0 262476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2853
timestamp 1676037725
transform 1 0 263580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2857
timestamp 1676037725
transform 1 0 263948 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2867
timestamp 1676037725
transform 1 0 264868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2879
timestamp 1676037725
transform 1 0 265972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2883
timestamp 1676037725
transform 1 0 266340 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2885
timestamp 1676037725
transform 1 0 266524 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2897
timestamp 1676037725
transform 1 0 267628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2909
timestamp 1676037725
transform 1 0 268732 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2913
timestamp 1676037725
transform 1 0 269100 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2925
timestamp 1676037725
transform 1 0 270204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2937
timestamp 1676037725
transform 1 0 271308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2941
timestamp 1676037725
transform 1 0 271676 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2949
timestamp 1676037725
transform 1 0 272412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2952
timestamp 1676037725
transform 1 0 272688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2962
timestamp 1676037725
transform 1 0 273608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2969
timestamp 1676037725
transform 1 0 274252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2973
timestamp 1676037725
transform 1 0 274620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2976
timestamp 1676037725
transform 1 0 274896 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2986
timestamp 1676037725
transform 1 0 275816 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2994
timestamp 1676037725
transform 1 0 276552 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2997
timestamp 1676037725
transform 1 0 276828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3009
timestamp 1676037725
transform 1 0 277932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3017
timestamp 1676037725
transform 1 0 278668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3022
timestamp 1676037725
transform 1 0 279128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3025
timestamp 1676037725
transform 1 0 279404 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3035
timestamp 1676037725
transform 1 0 280324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3047
timestamp 1676037725
transform 1 0 281428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3051
timestamp 1676037725
transform 1 0 281796 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3053
timestamp 1676037725
transform 1 0 281980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3065
timestamp 1676037725
transform 1 0 283084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3077
timestamp 1676037725
transform 1 0 284188 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3081
timestamp 1676037725
transform 1 0 284556 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3093
timestamp 1676037725
transform 1 0 285660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3105
timestamp 1676037725
transform 1 0 286764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3109
timestamp 1676037725
transform 1 0 287132 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3117
timestamp 1676037725
transform 1 0 287868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3120
timestamp 1676037725
transform 1 0 288144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3130
timestamp 1676037725
transform 1 0 289064 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3137
timestamp 1676037725
transform 1 0 289708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3143
timestamp 1676037725
transform 1 0 290260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3153
timestamp 1676037725
transform 1 0 291180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3161
timestamp 1676037725
transform 1 0 291916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3165
timestamp 1676037725
transform 1 0 292284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3169
timestamp 1676037725
transform 1 0 292652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3179
timestamp 1676037725
transform 1 0 293572 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3187
timestamp 1676037725
transform 1 0 294308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3190
timestamp 1676037725
transform 1 0 294584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3193
timestamp 1676037725
transform 1 0 294860 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3203
timestamp 1676037725
transform 1 0 295780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3215
timestamp 1676037725
transform 1 0 296884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3219
timestamp 1676037725
transform 1 0 297252 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3221
timestamp 1676037725
transform 1 0 297436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3233
timestamp 1676037725
transform 1 0 298540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3245
timestamp 1676037725
transform 1 0 299644 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3249
timestamp 1676037725
transform 1 0 300012 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3261
timestamp 1676037725
transform 1 0 301116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3273
timestamp 1676037725
transform 1 0 302220 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3277
timestamp 1676037725
transform 1 0 302588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3289
timestamp 1676037725
transform 1 0 303692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3301
timestamp 1676037725
transform 1 0 304796 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3305
timestamp 1676037725
transform 1 0 305164 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3317
timestamp 1676037725
transform 1 0 306268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3329
timestamp 1676037725
transform 1 0 307372 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3333
timestamp 1676037725
transform 1 0 307740 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3345
timestamp 1676037725
transform 1 0 308844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3357
timestamp 1676037725
transform 1 0 309948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3361
timestamp 1676037725
transform 1 0 310316 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3371
timestamp 1676037725
transform 1 0 311236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3383
timestamp 1676037725
transform 1 0 312340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3387
timestamp 1676037725
transform 1 0 312708 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3389
timestamp 1676037725
transform 1 0 312892 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3401
timestamp 1676037725
transform 1 0 313996 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3413
timestamp 1676037725
transform 1 0 315100 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3417
timestamp 1676037725
transform 1 0 315468 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3429
timestamp 1676037725
transform 1 0 316572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3441
timestamp 1676037725
transform 1 0 317676 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3445
timestamp 1676037725
transform 1 0 318044 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3457
timestamp 1676037725
transform 1 0 319148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3469
timestamp 1676037725
transform 1 0 320252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3473
timestamp 1676037725
transform 1 0 320620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3478
timestamp 1676037725
transform 1 0 321080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3491
timestamp 1676037725
transform 1 0 322276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3499
timestamp 1676037725
transform 1 0 323012 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3501
timestamp 1676037725
transform 1 0 323196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3513
timestamp 1676037725
transform 1 0 324300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3526
timestamp 1676037725
transform 1 0 325496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3529
timestamp 1676037725
transform 1 0 325772 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3539
timestamp 1676037725
transform 1 0 326692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3551
timestamp 1676037725
transform 1 0 327796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3555
timestamp 1676037725
transform 1 0 328164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3557
timestamp 1676037725
transform 1 0 328348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3569
timestamp 1676037725
transform 1 0 329452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3581
timestamp 1676037725
transform 1 0 330556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3585
timestamp 1676037725
transform 1 0 330924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3593
timestamp 1676037725
transform 1 0 331660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3610
timestamp 1676037725
transform 1 0 333224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3613
timestamp 1676037725
transform 1 0 333500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3617
timestamp 1676037725
transform 1 0 333868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3627
timestamp 1676037725
transform 1 0 334788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3631
timestamp 1676037725
transform 1 0 335156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3638
timestamp 1676037725
transform 1 0 335800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3641
timestamp 1676037725
transform 1 0 336076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3653
timestamp 1676037725
transform 1 0 337180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3666
timestamp 1676037725
transform 1 0 338376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3669
timestamp 1676037725
transform 1 0 338652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3681
timestamp 1676037725
transform 1 0 339756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3694
timestamp 1676037725
transform 1 0 340952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3697
timestamp 1676037725
transform 1 0 341228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3707
timestamp 1676037725
transform 1 0 342148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3713
timestamp 1676037725
transform 1 0 342700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3721
timestamp 1676037725
transform 1 0 343436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3725
timestamp 1676037725
transform 1 0 343804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3737
timestamp 1676037725
transform 1 0 344908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3749
timestamp 1676037725
transform 1 0 346012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3753
timestamp 1676037725
transform 1 0 346380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3765
timestamp 1676037725
transform 1 0 347484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3777
timestamp 1676037725
transform 1 0 348588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3781
timestamp 1676037725
transform 1 0 348956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3793
timestamp 1676037725
transform 1 0 350060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3805
timestamp 1676037725
transform 1 0 351164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3809
timestamp 1676037725
transform 1 0 351532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3821
timestamp 1676037725
transform 1 0 352636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3833
timestamp 1676037725
transform 1 0 353740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3837
timestamp 1676037725
transform 1 0 354108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3849
timestamp 1676037725
transform 1 0 355212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3861
timestamp 1676037725
transform 1 0 356316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3865
timestamp 1676037725
transform 1 0 356684 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3875
timestamp 1676037725
transform 1 0 357604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3887
timestamp 1676037725
transform 1 0 358708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3891
timestamp 1676037725
transform 1 0 359076 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3893
timestamp 1676037725
transform 1 0 359260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3905
timestamp 1676037725
transform 1 0 360364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3917
timestamp 1676037725
transform 1 0 361468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3921
timestamp 1676037725
transform 1 0 361836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3933
timestamp 1676037725
transform 1 0 362940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3945
timestamp 1676037725
transform 1 0 364044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3949
timestamp 1676037725
transform 1 0 364412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3961
timestamp 1676037725
transform 1 0 365516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3973
timestamp 1676037725
transform 1 0 366620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3977
timestamp 1676037725
transform 1 0 366988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3983
timestamp 1676037725
transform 1 0 367540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3993
timestamp 1676037725
transform 1 0 368460 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3999
timestamp 1676037725
transform 1 0 369012 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4002
timestamp 1676037725
transform 1 0 369288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4005
timestamp 1676037725
transform 1 0 369564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4016
timestamp 1676037725
transform 1 0 370576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4020
timestamp 1676037725
transform 1 0 370944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4030
timestamp 1676037725
transform 1 0 371864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4033
timestamp 1676037725
transform 1 0 372140 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4043
timestamp 1676037725
transform 1 0 373060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4055
timestamp 1676037725
transform 1 0 374164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4059
timestamp 1676037725
transform 1 0 374532 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4061
timestamp 1676037725
transform 1 0 374716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4073
timestamp 1676037725
transform 1 0 375820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4085
timestamp 1676037725
transform 1 0 376924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4089
timestamp 1676037725
transform 1 0 377292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4101
timestamp 1676037725
transform 1 0 378396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4113
timestamp 1676037725
transform 1 0 379500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4117
timestamp 1676037725
transform 1 0 379868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4129
timestamp 1676037725
transform 1 0 380972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4141
timestamp 1676037725
transform 1 0 382076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4145
timestamp 1676037725
transform 1 0 382444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4160
timestamp 1676037725
transform 1 0 383824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4170
timestamp 1676037725
transform 1 0 384744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4173
timestamp 1676037725
transform 1 0 385020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4184
timestamp 1676037725
transform 1 0 386032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4188
timestamp 1676037725
transform 1 0 386400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4198
timestamp 1676037725
transform 1 0 387320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4201
timestamp 1676037725
transform 1 0 387596 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4211
timestamp 1676037725
transform 1 0 388516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4223
timestamp 1676037725
transform 1 0 389620 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4227
timestamp 1676037725
transform 1 0 389988 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4229
timestamp 1676037725
transform 1 0 390172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4241
timestamp 1676037725
transform 1 0 391276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4253
timestamp 1676037725
transform 1 0 392380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4257
timestamp 1676037725
transform 1 0 392748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4269
timestamp 1676037725
transform 1 0 393852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4281
timestamp 1676037725
transform 1 0 394956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4285
timestamp 1676037725
transform 1 0 395324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4297
timestamp 1676037725
transform 1 0 396428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4309
timestamp 1676037725
transform 1 0 397532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4313
timestamp 1676037725
transform 1 0 397900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4325
timestamp 1676037725
transform 1 0 399004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4337
timestamp 1676037725
transform 1 0 400108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4341
timestamp 1676037725
transform 1 0 400476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4353
timestamp 1676037725
transform 1 0 401580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4365
timestamp 1676037725
transform 1 0 402684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4369
timestamp 1676037725
transform 1 0 403052 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4379
timestamp 1676037725
transform 1 0 403972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4391
timestamp 1676037725
transform 1 0 405076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4395
timestamp 1676037725
transform 1 0 405444 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4397
timestamp 1676037725
transform 1 0 405628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4409
timestamp 1676037725
transform 1 0 406732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4421
timestamp 1676037725
transform 1 0 407836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4425
timestamp 1676037725
transform 1 0 408204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4437
timestamp 1676037725
transform 1 0 409308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4449
timestamp 1676037725
transform 1 0 410412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4453
timestamp 1676037725
transform 1 0 410780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4465
timestamp 1676037725
transform 1 0 411884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4477
timestamp 1676037725
transform 1 0 412988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4481
timestamp 1676037725
transform 1 0 413356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4493
timestamp 1676037725
transform 1 0 414460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4501
timestamp 1676037725
transform 1 0 415196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4506
timestamp 1676037725
transform 1 0 415656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4509
timestamp 1676037725
transform 1 0 415932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4520
timestamp 1676037725
transform 1 0 416944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4524
timestamp 1676037725
transform 1 0 417312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4534
timestamp 1676037725
transform 1 0 418232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4537
timestamp 1676037725
transform 1 0 418508 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4547
timestamp 1676037725
transform 1 0 419428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4559
timestamp 1676037725
transform 1 0 420532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4563
timestamp 1676037725
transform 1 0 420900 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4565
timestamp 1676037725
transform 1 0 421084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4577
timestamp 1676037725
transform 1 0 422188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4589
timestamp 1676037725
transform 1 0 423292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4593
timestamp 1676037725
transform 1 0 423660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4605
timestamp 1676037725
transform 1 0 424764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4617
timestamp 1676037725
transform 1 0 425868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4621
timestamp 1676037725
transform 1 0 426236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4633
timestamp 1676037725
transform 1 0 427340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4639
timestamp 1676037725
transform 1 0 427892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4646
timestamp 1676037725
transform 1 0 428536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4649
timestamp 1676037725
transform 1 0 428812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4653
timestamp 1676037725
transform 1 0 429180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4657
timestamp 1676037725
transform 1 0 429548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4667
timestamp 1676037725
transform 1 0 430468 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4673
timestamp 1676037725
transform 1 0 431020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4677
timestamp 1676037725
transform 1 0 431388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4688
timestamp 1676037725
transform 1 0 432400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4701
timestamp 1676037725
transform 1 0 433596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4705
timestamp 1676037725
transform 1 0 433964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4715
timestamp 1676037725
transform 1 0 434884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4728
timestamp 1676037725
transform 1 0 436080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4733
timestamp 1676037725
transform 1 0 436540 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4737
timestamp 1676037725
transform 1 0 436908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4749
timestamp 1676037725
transform 1 0 438012 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4757
timestamp 1676037725
transform 1 0 438748 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4761
timestamp 1676037725
transform 1 0 439116 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4773
timestamp 1676037725
transform 1 0 440220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4785
timestamp 1676037725
transform 1 0 441324 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4789
timestamp 1676037725
transform 1 0 441692 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4801
timestamp 1676037725
transform 1 0 442796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4813
timestamp 1676037725
transform 1 0 443900 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4817
timestamp 1676037725
transform 1 0 444268 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4829
timestamp 1676037725
transform 1 0 445372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4841
timestamp 1676037725
transform 1 0 446476 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4845
timestamp 1676037725
transform 1 0 446844 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4857
timestamp 1676037725
transform 1 0 447948 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4869
timestamp 1676037725
transform 1 0 449052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4873
timestamp 1676037725
transform 1 0 449420 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4883
timestamp 1676037725
transform 1 0 450340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4895
timestamp 1676037725
transform 1 0 451444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4899
timestamp 1676037725
transform 1 0 451812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4901
timestamp 1676037725
transform 1 0 451996 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4913
timestamp 1676037725
transform 1 0 453100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4925
timestamp 1676037725
transform 1 0 454204 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4929
timestamp 1676037725
transform 1 0 454572 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4941
timestamp 1676037725
transform 1 0 455676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4953
timestamp 1676037725
transform 1 0 456780 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4957
timestamp 1676037725
transform 1 0 457148 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4969
timestamp 1676037725
transform 1 0 458252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4981
timestamp 1676037725
transform 1 0 459356 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4985
timestamp 1676037725
transform 1 0 459724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4997
timestamp 1676037725
transform 1 0 460828 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5005
timestamp 1676037725
transform 1 0 461564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5010
timestamp 1676037725
transform 1 0 462024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5013
timestamp 1676037725
transform 1 0 462300 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5027
timestamp 1676037725
transform 1 0 463588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5039
timestamp 1676037725
transform 1 0 464692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5041
timestamp 1676037725
transform 1 0 464876 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5051
timestamp 1676037725
transform 1 0 465796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5063
timestamp 1676037725
transform 1 0 466900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5067
timestamp 1676037725
transform 1 0 467268 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5069
timestamp 1676037725
transform 1 0 467452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5081
timestamp 1676037725
transform 1 0 468556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5093
timestamp 1676037725
transform 1 0 469660 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5097
timestamp 1676037725
transform 1 0 470028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5109
timestamp 1676037725
transform 1 0 471132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5121
timestamp 1676037725
transform 1 0 472236 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5125
timestamp 1676037725
transform 1 0 472604 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5137
timestamp 1676037725
transform 1 0 473708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5149
timestamp 1676037725
transform 1 0 474812 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5153
timestamp 1676037725
transform 1 0 475180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5165
timestamp 1676037725
transform 1 0 476284 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5173
timestamp 1676037725
transform 1 0 477020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5178
timestamp 1676037725
transform 1 0 477480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5181
timestamp 1676037725
transform 1 0 477756 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5195
timestamp 1676037725
transform 1 0 479044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5207
timestamp 1676037725
transform 1 0 480148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5209
timestamp 1676037725
transform 1 0 480332 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5219
timestamp 1676037725
transform 1 0 481252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5231
timestamp 1676037725
transform 1 0 482356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5235
timestamp 1676037725
transform 1 0 482724 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5237
timestamp 1676037725
transform 1 0 482908 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5249
timestamp 1676037725
transform 1 0 484012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5261
timestamp 1676037725
transform 1 0 485116 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5265
timestamp 1676037725
transform 1 0 485484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5277
timestamp 1676037725
transform 1 0 486588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5289
timestamp 1676037725
transform 1 0 487692 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5293
timestamp 1676037725
transform 1 0 488060 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5305
timestamp 1676037725
transform 1 0 489164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5317
timestamp 1676037725
transform 1 0 490268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5321
timestamp 1676037725
transform 1 0 490636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5333
timestamp 1676037725
transform 1 0 491740 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5345
timestamp 1676037725
transform 1 0 492844 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5349
timestamp 1676037725
transform 1 0 493212 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5361
timestamp 1676037725
transform 1 0 494316 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5373
timestamp 1676037725
transform 1 0 495420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5377
timestamp 1676037725
transform 1 0 495788 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5387
timestamp 1676037725
transform 1 0 496708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5399
timestamp 1676037725
transform 1 0 497812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5403
timestamp 1676037725
transform 1 0 498180 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5405
timestamp 1676037725
transform 1 0 498364 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5417
timestamp 1676037725
transform 1 0 499468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5429
timestamp 1676037725
transform 1 0 500572 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5433
timestamp 1676037725
transform 1 0 500940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5445
timestamp 1676037725
transform 1 0 502044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5457
timestamp 1676037725
transform 1 0 503148 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5461
timestamp 1676037725
transform 1 0 503516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5473
timestamp 1676037725
transform 1 0 504620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5485
timestamp 1676037725
transform 1 0 505724 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5489
timestamp 1676037725
transform 1 0 506092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5501
timestamp 1676037725
transform 1 0 507196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5513
timestamp 1676037725
transform 1 0 508300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5517
timestamp 1676037725
transform 1 0 508668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5525
timestamp 1676037725
transform 1 0 509404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5529
timestamp 1676037725
transform 1 0 509772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5542
timestamp 1676037725
transform 1 0 510968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5545
timestamp 1676037725
transform 1 0 511244 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5555
timestamp 1676037725
transform 1 0 512164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5567
timestamp 1676037725
transform 1 0 513268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5571
timestamp 1676037725
transform 1 0 513636 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5573
timestamp 1676037725
transform 1 0 513820 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5585
timestamp 1676037725
transform 1 0 514924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5597
timestamp 1676037725
transform 1 0 516028 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5601
timestamp 1676037725
transform 1 0 516396 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5613
timestamp 1676037725
transform 1 0 517500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5625
timestamp 1676037725
transform 1 0 518604 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5629
timestamp 1676037725
transform 1 0 518972 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5641
timestamp 1676037725
transform 1 0 520076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5653
timestamp 1676037725
transform 1 0 521180 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5657
timestamp 1676037725
transform 1 0 521548 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5669
timestamp 1676037725
transform 1 0 522652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5681
timestamp 1676037725
transform 1 0 523756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5685
timestamp 1676037725
transform 1 0 524124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5693
timestamp 1676037725
transform 1 0 524860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5697
timestamp 1676037725
transform 1 0 525228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5710
timestamp 1676037725
transform 1 0 526424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5713
timestamp 1676037725
transform 1 0 526700 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5723
timestamp 1676037725
transform 1 0 527620 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5738
timestamp 1676037725
transform 1 0 529000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5741
timestamp 1676037725
transform 1 0 529276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5754
timestamp 1676037725
transform 1 0 530472 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5760
timestamp 1676037725
transform 1 0 531024 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5769
timestamp 1676037725
transform 1 0 531852 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5781
timestamp 1676037725
transform 1 0 532956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5793
timestamp 1676037725
transform 1 0 534060 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5797
timestamp 1676037725
transform 1 0 534428 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5809
timestamp 1676037725
transform 1 0 535532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5821
timestamp 1676037725
transform 1 0 536636 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5825
timestamp 1676037725
transform 1 0 537004 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5837
timestamp 1676037725
transform 1 0 538108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5849
timestamp 1676037725
transform 1 0 539212 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5853
timestamp 1676037725
transform 1 0 539580 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5865
timestamp 1676037725
transform 1 0 540684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5877
timestamp 1676037725
transform 1 0 541788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5881
timestamp 1676037725
transform 1 0 542156 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5887
timestamp 1676037725
transform 1 0 542708 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5891
timestamp 1676037725
transform 1 0 543076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5897
timestamp 1676037725
transform 1 0 543628 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5905
timestamp 1676037725
transform 1 0 544364 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5909
timestamp 1676037725
transform 1 0 544732 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5921
timestamp 1676037725
transform 1 0 545836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5933
timestamp 1676037725
transform 1 0 546940 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5937
timestamp 1676037725
transform 1 0 547308 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5949
timestamp 1676037725
transform 1 0 548412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5961
timestamp 1676037725
transform 1 0 549516 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5965
timestamp 1676037725
transform 1 0 549884 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5977
timestamp 1676037725
transform 1 0 550988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5989
timestamp 1676037725
transform 1 0 552092 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5993
timestamp 1676037725
transform 1 0 552460 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6005
timestamp 1676037725
transform 1 0 553564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6017
timestamp 1676037725
transform 1 0 554668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6021
timestamp 1676037725
transform 1 0 555036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6026
timestamp 1676037725
transform 1 0 555496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6046
timestamp 1676037725
transform 1 0 557336 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6049
timestamp 1676037725
transform 1 0 557612 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6059
timestamp 1676037725
transform 1 0 558532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6071
timestamp 1676037725
transform 1 0 559636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6075
timestamp 1676037725
transform 1 0 560004 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6077
timestamp 1676037725
transform 1 0 560188 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6089
timestamp 1676037725
transform 1 0 561292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6101
timestamp 1676037725
transform 1 0 562396 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6105
timestamp 1676037725
transform 1 0 562764 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6117
timestamp 1676037725
transform 1 0 563868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6129
timestamp 1676037725
transform 1 0 564972 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6133
timestamp 1676037725
transform 1 0 565340 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6145
timestamp 1676037725
transform 1 0 566444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6157
timestamp 1676037725
transform 1 0 567548 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6161
timestamp 1676037725
transform 1 0 567916 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6173
timestamp 1676037725
transform 1 0 569020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6185
timestamp 1676037725
transform 1 0 570124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6189
timestamp 1676037725
transform 1 0 570492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6194
timestamp 1676037725
transform 1 0 570952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6214
timestamp 1676037725
transform 1 0 572792 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6217
timestamp 1676037725
transform 1 0 573068 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6227
timestamp 1676037725
transform 1 0 573988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6239
timestamp 1676037725
transform 1 0 575092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6243
timestamp 1676037725
transform 1 0 575460 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6245
timestamp 1676037725
transform 1 0 575644 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6257
timestamp 1676037725
transform 1 0 576748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6269
timestamp 1676037725
transform 1 0 577852 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6273
timestamp 1676037725
transform 1 0 578220 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6285
timestamp 1676037725
transform 1 0 579324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6297
timestamp 1676037725
transform 1 0 580428 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6301
timestamp 1676037725
transform 1 0 580796 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6313
timestamp 1676037725
transform 1 0 581900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6325
timestamp 1676037725
transform 1 0 583004 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6329
timestamp 1676037725
transform 1 0 583372 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6341
timestamp 1676037725
transform 1 0 584476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6353
timestamp 1676037725
transform 1 0 585580 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6357
timestamp 1676037725
transform 1 0 585948 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6369
timestamp 1676037725
transform 1 0 587052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6381
timestamp 1676037725
transform 1 0 588156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6385
timestamp 1676037725
transform 1 0 588524 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6395
timestamp 1676037725
transform 1 0 589444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6407
timestamp 1676037725
transform 1 0 590548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6411
timestamp 1676037725
transform 1 0 590916 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6413
timestamp 1676037725
transform 1 0 591100 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6425
timestamp 1676037725
transform 1 0 592204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6437
timestamp 1676037725
transform 1 0 593308 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6441
timestamp 1676037725
transform 1 0 593676 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6453
timestamp 1676037725
transform 1 0 594780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6465
timestamp 1676037725
transform 1 0 595884 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6469
timestamp 1676037725
transform 1 0 596252 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6481
timestamp 1676037725
transform 1 0 597356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6493
timestamp 1676037725
transform 1 0 598460 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6497
timestamp 1676037725
transform 1 0 598828 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6509
timestamp 1676037725
transform 1 0 599932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6521
timestamp 1676037725
transform 1 0 601036 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6525
timestamp 1676037725
transform 1 0 601404 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6537
timestamp 1676037725
transform 1 0 602508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6549
timestamp 1676037725
transform 1 0 603612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6553
timestamp 1676037725
transform 1 0 603980 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6563
timestamp 1676037725
transform 1 0 604900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6575
timestamp 1676037725
transform 1 0 606004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6579
timestamp 1676037725
transform 1 0 606372 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6581
timestamp 1676037725
transform 1 0 606556 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6593
timestamp 1676037725
transform 1 0 607660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6605
timestamp 1676037725
transform 1 0 608764 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6609
timestamp 1676037725
transform 1 0 609132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6621
timestamp 1676037725
transform 1 0 610236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6633
timestamp 1676037725
transform 1 0 611340 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6637
timestamp 1676037725
transform 1 0 611708 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6649
timestamp 1676037725
transform 1 0 612812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6661
timestamp 1676037725
transform 1 0 613916 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6665
timestamp 1676037725
transform 1 0 614284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6677
timestamp 1676037725
transform 1 0 615388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6689
timestamp 1676037725
transform 1 0 616492 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6693
timestamp 1676037725
transform 1 0 616860 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6705
timestamp 1676037725
transform 1 0 617964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6717
timestamp 1676037725
transform 1 0 619068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6721
timestamp 1676037725
transform 1 0 619436 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6731
timestamp 1676037725
transform 1 0 620356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6743
timestamp 1676037725
transform 1 0 621460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6747
timestamp 1676037725
transform 1 0 621828 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6749
timestamp 1676037725
transform 1 0 622012 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6757
timestamp 1676037725
transform 1 0 622748 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6764
timestamp 1676037725
transform 1 0 623392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6777
timestamp 1676037725
transform 1 0 624588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6788
timestamp 1676037725
transform 1 0 625600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6794
timestamp 1676037725
transform 1 0 626152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6802
timestamp 1676037725
transform 1 0 626888 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6805
timestamp 1676037725
transform 1 0 627164 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6817
timestamp 1676037725
transform 1 0 628268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6829
timestamp 1676037725
transform 1 0 629372 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6833
timestamp 1676037725
transform 1 0 629740 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6845
timestamp 1676037725
transform 1 0 630844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6857
timestamp 1676037725
transform 1 0 631948 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6861
timestamp 1676037725
transform 1 0 632316 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6873
timestamp 1676037725
transform 1 0 633420 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6885
timestamp 1676037725
transform 1 0 634524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6889
timestamp 1676037725
transform 1 0 634892 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6895
timestamp 1676037725
transform 1 0 635444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6899
timestamp 1676037725
transform 1 0 635812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6905
timestamp 1676037725
transform 1 0 636364 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6913
timestamp 1676037725
transform 1 0 637100 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6917
timestamp 1676037725
transform 1 0 637468 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6929
timestamp 1676037725
transform 1 0 638572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6941
timestamp 1676037725
transform 1 0 639676 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6945
timestamp 1676037725
transform 1 0 640044 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6957
timestamp 1676037725
transform 1 0 641148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6969
timestamp 1676037725
transform 1 0 642252 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6973
timestamp 1676037725
transform 1 0 642620 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6985
timestamp 1676037725
transform 1 0 643724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6997
timestamp 1676037725
transform 1 0 644828 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7001
timestamp 1676037725
transform 1 0 645196 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7013
timestamp 1676037725
transform 1 0 646300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7025
timestamp 1676037725
transform 1 0 647404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7029
timestamp 1676037725
transform 1 0 647772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7041
timestamp 1676037725
transform 1 0 648876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7053
timestamp 1676037725
transform 1 0 649980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7057
timestamp 1676037725
transform 1 0 650348 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7067
timestamp 1676037725
transform 1 0 651268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7079
timestamp 1676037725
transform 1 0 652372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7083
timestamp 1676037725
transform 1 0 652740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7085
timestamp 1676037725
transform 1 0 652924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7097
timestamp 1676037725
transform 1 0 654028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7109
timestamp 1676037725
transform 1 0 655132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7113
timestamp 1676037725
transform 1 0 655500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7125
timestamp 1676037725
transform 1 0 656604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7137
timestamp 1676037725
transform 1 0 657708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7141
timestamp 1676037725
transform 1 0 658076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7153
timestamp 1676037725
transform 1 0 659180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7165
timestamp 1676037725
transform 1 0 660284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7169
timestamp 1676037725
transform 1 0 660652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7181
timestamp 1676037725
transform 1 0 661756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7193
timestamp 1676037725
transform 1 0 662860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7197
timestamp 1676037725
transform 1 0 663228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7209
timestamp 1676037725
transform 1 0 664332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7221
timestamp 1676037725
transform 1 0 665436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7225
timestamp 1676037725
transform 1 0 665804 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7235
timestamp 1676037725
transform 1 0 666724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7247
timestamp 1676037725
transform 1 0 667828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7251
timestamp 1676037725
transform 1 0 668196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7253
timestamp 1676037725
transform 1 0 668380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7265
timestamp 1676037725
transform 1 0 669484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7277
timestamp 1676037725
transform 1 0 670588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7281
timestamp 1676037725
transform 1 0 670956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7293
timestamp 1676037725
transform 1 0 672060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7305
timestamp 1676037725
transform 1 0 673164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7309
timestamp 1676037725
transform 1 0 673532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7321
timestamp 1676037725
transform 1 0 674636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7333
timestamp 1676037725
transform 1 0 675740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7337
timestamp 1676037725
transform 1 0 676108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7349
timestamp 1676037725
transform 1 0 677212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7361
timestamp 1676037725
transform 1 0 678316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7365
timestamp 1676037725
transform 1 0 678684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7377
timestamp 1676037725
transform 1 0 679788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7389
timestamp 1676037725
transform 1 0 680892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7393
timestamp 1676037725
transform 1 0 681260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7403
timestamp 1676037725
transform 1 0 682180 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1676037725
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1676037725
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1676037725
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1676037725
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1676037725
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1676037725
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1676037725
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1676037725
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1676037725
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1676037725
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1676037725
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1676037725
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1676037725
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1676037725
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1676037725
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1676037725
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1676037725
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1676037725
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1676037725
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1676037725
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1676037725
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1676037725
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1676037725
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1676037725
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1676037725
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1676037725
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1676037725
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1676037725
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1676037725
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1676037725
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1676037725
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1676037725
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_841
timestamp 1676037725
transform 1 0 78476 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_847
timestamp 1676037725
transform 1 0 79028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_859
timestamp 1676037725
transform 1 0 80132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_871
timestamp 1676037725
transform 1 0 81236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_883
timestamp 1676037725
transform 1 0 82340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1676037725
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1676037725
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1676037725
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1676037725
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1676037725
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1676037725
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1676037725
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1676037725
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1676037725
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1676037725
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1676037725
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1676037725
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1676037725
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1676037725
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1676037725
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1676037725
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1676037725
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1676037725
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1676037725
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1676037725
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1676037725
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1676037725
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1676037725
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1676037725
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1676037725
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1676037725
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1676037725
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1676037725
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1157
timestamp 1676037725
transform 1 0 107548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1676037725
transform 1 0 108652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1676037725
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1177
timestamp 1676037725
transform 1 0 109388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1189
timestamp 1676037725
transform 1 0 110492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1201
timestamp 1676037725
transform 1 0 111596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1213
timestamp 1676037725
transform 1 0 112700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1225
timestamp 1676037725
transform 1 0 113804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1676037725
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1233
timestamp 1676037725
transform 1 0 114540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1245
timestamp 1676037725
transform 1 0 115644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1257
timestamp 1676037725
transform 1 0 116748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1269
timestamp 1676037725
transform 1 0 117852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1281
timestamp 1676037725
transform 1 0 118956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1287
timestamp 1676037725
transform 1 0 119508 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1289
timestamp 1676037725
transform 1 0 119692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1301
timestamp 1676037725
transform 1 0 120796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1313
timestamp 1676037725
transform 1 0 121900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1325
timestamp 1676037725
transform 1 0 123004 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1337
timestamp 1676037725
transform 1 0 124108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1343
timestamp 1676037725
transform 1 0 124660 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1345
timestamp 1676037725
transform 1 0 124844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1357
timestamp 1676037725
transform 1 0 125948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1369
timestamp 1676037725
transform 1 0 127052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1381
timestamp 1676037725
transform 1 0 128156 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1393
timestamp 1676037725
transform 1 0 129260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1399
timestamp 1676037725
transform 1 0 129812 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1401
timestamp 1676037725
transform 1 0 129996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1413
timestamp 1676037725
transform 1 0 131100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1425
timestamp 1676037725
transform 1 0 132204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1437
timestamp 1676037725
transform 1 0 133308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1449
timestamp 1676037725
transform 1 0 134412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1455
timestamp 1676037725
transform 1 0 134964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1457
timestamp 1676037725
transform 1 0 135148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1469
timestamp 1676037725
transform 1 0 136252 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1472
timestamp 1676037725
transform 1 0 136528 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1484
timestamp 1676037725
transform 1 0 137632 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1496
timestamp 1676037725
transform 1 0 138736 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1508
timestamp 1676037725
transform 1 0 139840 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1513
timestamp 1676037725
transform 1 0 140300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1525
timestamp 1676037725
transform 1 0 141404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1537
timestamp 1676037725
transform 1 0 142508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1549
timestamp 1676037725
transform 1 0 143612 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1561
timestamp 1676037725
transform 1 0 144716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1567
timestamp 1676037725
transform 1 0 145268 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1569
timestamp 1676037725
transform 1 0 145452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1581
timestamp 1676037725
transform 1 0 146556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1593
timestamp 1676037725
transform 1 0 147660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1605
timestamp 1676037725
transform 1 0 148764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1617
timestamp 1676037725
transform 1 0 149868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1623
timestamp 1676037725
transform 1 0 150420 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1625
timestamp 1676037725
transform 1 0 150604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1637
timestamp 1676037725
transform 1 0 151708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1649
timestamp 1676037725
transform 1 0 152812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1661
timestamp 1676037725
transform 1 0 153916 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1673
timestamp 1676037725
transform 1 0 155020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1679
timestamp 1676037725
transform 1 0 155572 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1681
timestamp 1676037725
transform 1 0 155756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1693
timestamp 1676037725
transform 1 0 156860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1705
timestamp 1676037725
transform 1 0 157964 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1717
timestamp 1676037725
transform 1 0 159068 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1729
timestamp 1676037725
transform 1 0 160172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1735
timestamp 1676037725
transform 1 0 160724 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1737
timestamp 1676037725
transform 1 0 160908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1749
timestamp 1676037725
transform 1 0 162012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1761
timestamp 1676037725
transform 1 0 163116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1773
timestamp 1676037725
transform 1 0 164220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1785
timestamp 1676037725
transform 1 0 165324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1791
timestamp 1676037725
transform 1 0 165876 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1793
timestamp 1676037725
transform 1 0 166060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1805
timestamp 1676037725
transform 1 0 167164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1817
timestamp 1676037725
transform 1 0 168268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1829
timestamp 1676037725
transform 1 0 169372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1841
timestamp 1676037725
transform 1 0 170476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1847
timestamp 1676037725
transform 1 0 171028 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1849
timestamp 1676037725
transform 1 0 171212 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1855
timestamp 1676037725
transform 1 0 171764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1867
timestamp 1676037725
transform 1 0 172868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1879
timestamp 1676037725
transform 1 0 173972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1891
timestamp 1676037725
transform 1 0 175076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1903
timestamp 1676037725
transform 1 0 176180 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1905
timestamp 1676037725
transform 1 0 176364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1917
timestamp 1676037725
transform 1 0 177468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1929
timestamp 1676037725
transform 1 0 178572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1941
timestamp 1676037725
transform 1 0 179676 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1953
timestamp 1676037725
transform 1 0 180780 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1959
timestamp 1676037725
transform 1 0 181332 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1961
timestamp 1676037725
transform 1 0 181516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1973
timestamp 1676037725
transform 1 0 182620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1985
timestamp 1676037725
transform 1 0 183724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1997
timestamp 1676037725
transform 1 0 184828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2009
timestamp 1676037725
transform 1 0 185932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2015
timestamp 1676037725
transform 1 0 186484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2017
timestamp 1676037725
transform 1 0 186668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2025
timestamp 1676037725
transform 1 0 187404 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2029
timestamp 1676037725
transform 1 0 187772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2041
timestamp 1676037725
transform 1 0 188876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2053
timestamp 1676037725
transform 1 0 189980 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2065
timestamp 1676037725
transform 1 0 191084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2071
timestamp 1676037725
transform 1 0 191636 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2073
timestamp 1676037725
transform 1 0 191820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2085
timestamp 1676037725
transform 1 0 192924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2097
timestamp 1676037725
transform 1 0 194028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2109
timestamp 1676037725
transform 1 0 195132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2121
timestamp 1676037725
transform 1 0 196236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2127
timestamp 1676037725
transform 1 0 196788 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2129
timestamp 1676037725
transform 1 0 196972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2141
timestamp 1676037725
transform 1 0 198076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2153
timestamp 1676037725
transform 1 0 199180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2165
timestamp 1676037725
transform 1 0 200284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2177
timestamp 1676037725
transform 1 0 201388 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2183
timestamp 1676037725
transform 1 0 201940 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2185
timestamp 1676037725
transform 1 0 202124 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_2193
timestamp 1676037725
transform 1 0 202860 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2197
timestamp 1676037725
transform 1 0 203228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2209
timestamp 1676037725
transform 1 0 204332 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2221
timestamp 1676037725
transform 1 0 205436 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2233
timestamp 1676037725
transform 1 0 206540 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2239
timestamp 1676037725
transform 1 0 207092 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2241
timestamp 1676037725
transform 1 0 207276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2253
timestamp 1676037725
transform 1 0 208380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2265
timestamp 1676037725
transform 1 0 209484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2277
timestamp 1676037725
transform 1 0 210588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2289
timestamp 1676037725
transform 1 0 211692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2295
timestamp 1676037725
transform 1 0 212244 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2297
timestamp 1676037725
transform 1 0 212428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2309
timestamp 1676037725
transform 1 0 213532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2321
timestamp 1676037725
transform 1 0 214636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2333
timestamp 1676037725
transform 1 0 215740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2345
timestamp 1676037725
transform 1 0 216844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2351
timestamp 1676037725
transform 1 0 217396 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2353
timestamp 1676037725
transform 1 0 217580 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2359
timestamp 1676037725
transform 1 0 218132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2371
timestamp 1676037725
transform 1 0 219236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2383
timestamp 1676037725
transform 1 0 220340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2395
timestamp 1676037725
transform 1 0 221444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2407
timestamp 1676037725
transform 1 0 222548 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2409
timestamp 1676037725
transform 1 0 222732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2421
timestamp 1676037725
transform 1 0 223836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2433
timestamp 1676037725
transform 1 0 224940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2445
timestamp 1676037725
transform 1 0 226044 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2457
timestamp 1676037725
transform 1 0 227148 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2463
timestamp 1676037725
transform 1 0 227700 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2465
timestamp 1676037725
transform 1 0 227884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2477
timestamp 1676037725
transform 1 0 228988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2489
timestamp 1676037725
transform 1 0 230092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2501
timestamp 1676037725
transform 1 0 231196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2513
timestamp 1676037725
transform 1 0 232300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2519
timestamp 1676037725
transform 1 0 232852 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2521
timestamp 1676037725
transform 1 0 233036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2533
timestamp 1676037725
transform 1 0 234140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2545
timestamp 1676037725
transform 1 0 235244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2557
timestamp 1676037725
transform 1 0 236348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2569
timestamp 1676037725
transform 1 0 237452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2575
timestamp 1676037725
transform 1 0 238004 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2577
timestamp 1676037725
transform 1 0 238188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2589
timestamp 1676037725
transform 1 0 239292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2601
timestamp 1676037725
transform 1 0 240396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2613
timestamp 1676037725
transform 1 0 241500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2625
timestamp 1676037725
transform 1 0 242604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2631
timestamp 1676037725
transform 1 0 243156 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2633
timestamp 1676037725
transform 1 0 243340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2645
timestamp 1676037725
transform 1 0 244444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2657
timestamp 1676037725
transform 1 0 245548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2669
timestamp 1676037725
transform 1 0 246652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2681
timestamp 1676037725
transform 1 0 247756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2687
timestamp 1676037725
transform 1 0 248308 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2689
timestamp 1676037725
transform 1 0 248492 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2699
timestamp 1676037725
transform 1 0 249412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2711
timestamp 1676037725
transform 1 0 250516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2723
timestamp 1676037725
transform 1 0 251620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2735
timestamp 1676037725
transform 1 0 252724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2743
timestamp 1676037725
transform 1 0 253460 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2745
timestamp 1676037725
transform 1 0 253644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2757
timestamp 1676037725
transform 1 0 254748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2769
timestamp 1676037725
transform 1 0 255852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2781
timestamp 1676037725
transform 1 0 256956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2793
timestamp 1676037725
transform 1 0 258060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2799
timestamp 1676037725
transform 1 0 258612 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2801
timestamp 1676037725
transform 1 0 258796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2813
timestamp 1676037725
transform 1 0 259900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2825
timestamp 1676037725
transform 1 0 261004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2837
timestamp 1676037725
transform 1 0 262108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2849
timestamp 1676037725
transform 1 0 263212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2855
timestamp 1676037725
transform 1 0 263764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_2857
timestamp 1676037725
transform 1 0 263948 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2863
timestamp 1676037725
transform 1 0 264500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2875
timestamp 1676037725
transform 1 0 265604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2887
timestamp 1676037725
transform 1 0 266708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2899
timestamp 1676037725
transform 1 0 267812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2911
timestamp 1676037725
transform 1 0 268916 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2913
timestamp 1676037725
transform 1 0 269100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2925
timestamp 1676037725
transform 1 0 270204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2937
timestamp 1676037725
transform 1 0 271308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2949
timestamp 1676037725
transform 1 0 272412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2961
timestamp 1676037725
transform 1 0 273516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2967
timestamp 1676037725
transform 1 0 274068 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2969
timestamp 1676037725
transform 1 0 274252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2981
timestamp 1676037725
transform 1 0 275356 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2993
timestamp 1676037725
transform 1 0 276460 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3003
timestamp 1676037725
transform 1 0 277380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3015
timestamp 1676037725
transform 1 0 278484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3019
timestamp 1676037725
transform 1 0 278852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3022
timestamp 1676037725
transform 1 0 279128 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3025
timestamp 1676037725
transform 1 0 279404 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3033
timestamp 1676037725
transform 1 0 280140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3045
timestamp 1676037725
transform 1 0 281244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3057
timestamp 1676037725
transform 1 0 282348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3069
timestamp 1676037725
transform 1 0 283452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3077
timestamp 1676037725
transform 1 0 284188 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3081
timestamp 1676037725
transform 1 0 284556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3093
timestamp 1676037725
transform 1 0 285660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3105
timestamp 1676037725
transform 1 0 286764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3117
timestamp 1676037725
transform 1 0 287868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3129
timestamp 1676037725
transform 1 0 288972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3135
timestamp 1676037725
transform 1 0 289524 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3137
timestamp 1676037725
transform 1 0 289708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3149
timestamp 1676037725
transform 1 0 290812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3161
timestamp 1676037725
transform 1 0 291916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3167
timestamp 1676037725
transform 1 0 292468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3170
timestamp 1676037725
transform 1 0 292744 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3182
timestamp 1676037725
transform 1 0 293848 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3190
timestamp 1676037725
transform 1 0 294584 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3193
timestamp 1676037725
transform 1 0 294860 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3204
timestamp 1676037725
transform 1 0 295872 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3216
timestamp 1676037725
transform 1 0 296976 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3228
timestamp 1676037725
transform 1 0 298080 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3240
timestamp 1676037725
transform 1 0 299184 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3249
timestamp 1676037725
transform 1 0 300012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3261
timestamp 1676037725
transform 1 0 301116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3273
timestamp 1676037725
transform 1 0 302220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3285
timestamp 1676037725
transform 1 0 303324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3297
timestamp 1676037725
transform 1 0 304428 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3303
timestamp 1676037725
transform 1 0 304980 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3305
timestamp 1676037725
transform 1 0 305164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3317
timestamp 1676037725
transform 1 0 306268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3329
timestamp 1676037725
transform 1 0 307372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3341
timestamp 1676037725
transform 1 0 308476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3353
timestamp 1676037725
transform 1 0 309580 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3359
timestamp 1676037725
transform 1 0 310132 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3361
timestamp 1676037725
transform 1 0 310316 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3367
timestamp 1676037725
transform 1 0 310868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3379
timestamp 1676037725
transform 1 0 311972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3391
timestamp 1676037725
transform 1 0 313076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3403
timestamp 1676037725
transform 1 0 314180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3415
timestamp 1676037725
transform 1 0 315284 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3417
timestamp 1676037725
transform 1 0 315468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3429
timestamp 1676037725
transform 1 0 316572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3441
timestamp 1676037725
transform 1 0 317676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3453
timestamp 1676037725
transform 1 0 318780 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3465
timestamp 1676037725
transform 1 0 319884 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3471
timestamp 1676037725
transform 1 0 320436 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3473
timestamp 1676037725
transform 1 0 320620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3485
timestamp 1676037725
transform 1 0 321724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3497
timestamp 1676037725
transform 1 0 322828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3501
timestamp 1676037725
transform 1 0 323196 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3504
timestamp 1676037725
transform 1 0 323472 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3512
timestamp 1676037725
transform 1 0 324208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3517
timestamp 1676037725
transform 1 0 324668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3525
timestamp 1676037725
transform 1 0 325404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3529
timestamp 1676037725
transform 1 0 325772 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3535
timestamp 1676037725
transform 1 0 326324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3547
timestamp 1676037725
transform 1 0 327428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3559
timestamp 1676037725
transform 1 0 328532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3571
timestamp 1676037725
transform 1 0 329636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3583
timestamp 1676037725
transform 1 0 330740 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3585
timestamp 1676037725
transform 1 0 330924 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3595
timestamp 1676037725
transform 1 0 331844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3607
timestamp 1676037725
transform 1 0 332948 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3612
timestamp 1676037725
transform 1 0 333408 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3624
timestamp 1676037725
transform 1 0 334512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3629
timestamp 1676037725
transform 1 0 334972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3635
timestamp 1676037725
transform 1 0 335524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3638
timestamp 1676037725
transform 1 0 335800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3641
timestamp 1676037725
transform 1 0 336076 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3647
timestamp 1676037725
transform 1 0 336628 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3657
timestamp 1676037725
transform 1 0 337548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3665
timestamp 1676037725
transform 1 0 338284 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3668
timestamp 1676037725
transform 1 0 338560 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3681
timestamp 1676037725
transform 1 0 339756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3687
timestamp 1676037725
transform 1 0 340308 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3695
timestamp 1676037725
transform 1 0 341044 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3697
timestamp 1676037725
transform 1 0 341228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3708
timestamp 1676037725
transform 1 0 342240 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3714
timestamp 1676037725
transform 1 0 342792 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3726
timestamp 1676037725
transform 1 0 343896 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3738
timestamp 1676037725
transform 1 0 345000 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3750
timestamp 1676037725
transform 1 0 346104 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3753
timestamp 1676037725
transform 1 0 346380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3765
timestamp 1676037725
transform 1 0 347484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3777
timestamp 1676037725
transform 1 0 348588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3789
timestamp 1676037725
transform 1 0 349692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3801
timestamp 1676037725
transform 1 0 350796 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3807
timestamp 1676037725
transform 1 0 351348 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3809
timestamp 1676037725
transform 1 0 351532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3821
timestamp 1676037725
transform 1 0 352636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3833
timestamp 1676037725
transform 1 0 353740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3845
timestamp 1676037725
transform 1 0 354844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3857
timestamp 1676037725
transform 1 0 355948 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3863
timestamp 1676037725
transform 1 0 356500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3865
timestamp 1676037725
transform 1 0 356684 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3871
timestamp 1676037725
transform 1 0 357236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3883
timestamp 1676037725
transform 1 0 358340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3895
timestamp 1676037725
transform 1 0 359444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3907
timestamp 1676037725
transform 1 0 360548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3919
timestamp 1676037725
transform 1 0 361652 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3921
timestamp 1676037725
transform 1 0 361836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3933
timestamp 1676037725
transform 1 0 362940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3945
timestamp 1676037725
transform 1 0 364044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3957
timestamp 1676037725
transform 1 0 365148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3969
timestamp 1676037725
transform 1 0 366252 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3975
timestamp 1676037725
transform 1 0 366804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3977
timestamp 1676037725
transform 1 0 366988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3981
timestamp 1676037725
transform 1 0 367356 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3984
timestamp 1676037725
transform 1 0 367632 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3996
timestamp 1676037725
transform 1 0 368736 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4008
timestamp 1676037725
transform 1 0 369840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_4016
timestamp 1676037725
transform 1 0 370576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4021
timestamp 1676037725
transform 1 0 371036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_4029
timestamp 1676037725
transform 1 0 371772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4033
timestamp 1676037725
transform 1 0 372140 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4039
timestamp 1676037725
transform 1 0 372692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4051
timestamp 1676037725
transform 1 0 373796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4063
timestamp 1676037725
transform 1 0 374900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4075
timestamp 1676037725
transform 1 0 376004 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4087
timestamp 1676037725
transform 1 0 377108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4089
timestamp 1676037725
transform 1 0 377292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4101
timestamp 1676037725
transform 1 0 378396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4113
timestamp 1676037725
transform 1 0 379500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4125
timestamp 1676037725
transform 1 0 380604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4137
timestamp 1676037725
transform 1 0 381708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4143
timestamp 1676037725
transform 1 0 382260 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4145
timestamp 1676037725
transform 1 0 382444 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4151
timestamp 1676037725
transform 1 0 382996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4163
timestamp 1676037725
transform 1 0 384100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4175
timestamp 1676037725
transform 1 0 385204 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4189
timestamp 1676037725
transform 1 0 386492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_4197
timestamp 1676037725
transform 1 0 387228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4201
timestamp 1676037725
transform 1 0 387596 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4207
timestamp 1676037725
transform 1 0 388148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4219
timestamp 1676037725
transform 1 0 389252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4231
timestamp 1676037725
transform 1 0 390356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4243
timestamp 1676037725
transform 1 0 391460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4255
timestamp 1676037725
transform 1 0 392564 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4257
timestamp 1676037725
transform 1 0 392748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4269
timestamp 1676037725
transform 1 0 393852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4281
timestamp 1676037725
transform 1 0 394956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4293
timestamp 1676037725
transform 1 0 396060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4305
timestamp 1676037725
transform 1 0 397164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4311
timestamp 1676037725
transform 1 0 397716 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4313
timestamp 1676037725
transform 1 0 397900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4325
timestamp 1676037725
transform 1 0 399004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4337
timestamp 1676037725
transform 1 0 400108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4349
timestamp 1676037725
transform 1 0 401212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4361
timestamp 1676037725
transform 1 0 402316 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4367
timestamp 1676037725
transform 1 0 402868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4369
timestamp 1676037725
transform 1 0 403052 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4375
timestamp 1676037725
transform 1 0 403604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4387
timestamp 1676037725
transform 1 0 404708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4399
timestamp 1676037725
transform 1 0 405812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4411
timestamp 1676037725
transform 1 0 406916 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4423
timestamp 1676037725
transform 1 0 408020 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4425
timestamp 1676037725
transform 1 0 408204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4437
timestamp 1676037725
transform 1 0 409308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4449
timestamp 1676037725
transform 1 0 410412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4461
timestamp 1676037725
transform 1 0 411516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4473
timestamp 1676037725
transform 1 0 412620 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4479
timestamp 1676037725
transform 1 0 413172 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4481
timestamp 1676037725
transform 1 0 413356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4493
timestamp 1676037725
transform 1 0 414460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4505
timestamp 1676037725
transform 1 0 415564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4517
timestamp 1676037725
transform 1 0 416668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4525
timestamp 1676037725
transform 1 0 417404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_4533
timestamp 1676037725
transform 1 0 418140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4537
timestamp 1676037725
transform 1 0 418508 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4543
timestamp 1676037725
transform 1 0 419060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4555
timestamp 1676037725
transform 1 0 420164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4567
timestamp 1676037725
transform 1 0 421268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4579
timestamp 1676037725
transform 1 0 422372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4591
timestamp 1676037725
transform 1 0 423476 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4593
timestamp 1676037725
transform 1 0 423660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4605
timestamp 1676037725
transform 1 0 424764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4617
timestamp 1676037725
transform 1 0 425868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4629
timestamp 1676037725
transform 1 0 426972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4641
timestamp 1676037725
transform 1 0 428076 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4647
timestamp 1676037725
transform 1 0 428628 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4649
timestamp 1676037725
transform 1 0 428812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4661
timestamp 1676037725
transform 1 0 429916 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4669
timestamp 1676037725
transform 1 0 430652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4672
timestamp 1676037725
transform 1 0 430928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_4685
timestamp 1676037725
transform 1 0 432124 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4702
timestamp 1676037725
transform 1 0 433688 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4705
timestamp 1676037725
transform 1 0 433964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4716
timestamp 1676037725
transform 1 0 434976 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4722
timestamp 1676037725
transform 1 0 435528 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4734
timestamp 1676037725
transform 1 0 436632 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4746
timestamp 1676037725
transform 1 0 437736 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_4758
timestamp 1676037725
transform 1 0 438840 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4761
timestamp 1676037725
transform 1 0 439116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4773
timestamp 1676037725
transform 1 0 440220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4785
timestamp 1676037725
transform 1 0 441324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4797
timestamp 1676037725
transform 1 0 442428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4809
timestamp 1676037725
transform 1 0 443532 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4815
timestamp 1676037725
transform 1 0 444084 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4817
timestamp 1676037725
transform 1 0 444268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4829
timestamp 1676037725
transform 1 0 445372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4841
timestamp 1676037725
transform 1 0 446476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4853
timestamp 1676037725
transform 1 0 447580 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4865
timestamp 1676037725
transform 1 0 448684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4871
timestamp 1676037725
transform 1 0 449236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_4873
timestamp 1676037725
transform 1 0 449420 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4879
timestamp 1676037725
transform 1 0 449972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4891
timestamp 1676037725
transform 1 0 451076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4903
timestamp 1676037725
transform 1 0 452180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4915
timestamp 1676037725
transform 1 0 453284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4927
timestamp 1676037725
transform 1 0 454388 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4929
timestamp 1676037725
transform 1 0 454572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4941
timestamp 1676037725
transform 1 0 455676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4953
timestamp 1676037725
transform 1 0 456780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4965
timestamp 1676037725
transform 1 0 457884 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4977
timestamp 1676037725
transform 1 0 458988 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4983
timestamp 1676037725
transform 1 0 459540 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4985
timestamp 1676037725
transform 1 0 459724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4997
timestamp 1676037725
transform 1 0 460828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5009
timestamp 1676037725
transform 1 0 461932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5021
timestamp 1676037725
transform 1 0 463036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5025
timestamp 1676037725
transform 1 0 463404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5038
timestamp 1676037725
transform 1 0 464600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5041
timestamp 1676037725
transform 1 0 464876 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5047
timestamp 1676037725
transform 1 0 465428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5059
timestamp 1676037725
transform 1 0 466532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5071
timestamp 1676037725
transform 1 0 467636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5083
timestamp 1676037725
transform 1 0 468740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5095
timestamp 1676037725
transform 1 0 469844 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5097
timestamp 1676037725
transform 1 0 470028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5109
timestamp 1676037725
transform 1 0 471132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5121
timestamp 1676037725
transform 1 0 472236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5133
timestamp 1676037725
transform 1 0 473340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5145
timestamp 1676037725
transform 1 0 474444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5151
timestamp 1676037725
transform 1 0 474996 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5153
timestamp 1676037725
transform 1 0 475180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5165
timestamp 1676037725
transform 1 0 476284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5177
timestamp 1676037725
transform 1 0 477388 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5189
timestamp 1676037725
transform 1 0 478492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5193
timestamp 1676037725
transform 1 0 478860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5206
timestamp 1676037725
transform 1 0 480056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5209
timestamp 1676037725
transform 1 0 480332 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5215
timestamp 1676037725
transform 1 0 480884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5227
timestamp 1676037725
transform 1 0 481988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5239
timestamp 1676037725
transform 1 0 483092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5251
timestamp 1676037725
transform 1 0 484196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5263
timestamp 1676037725
transform 1 0 485300 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5265
timestamp 1676037725
transform 1 0 485484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5277
timestamp 1676037725
transform 1 0 486588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5289
timestamp 1676037725
transform 1 0 487692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5301
timestamp 1676037725
transform 1 0 488796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5313
timestamp 1676037725
transform 1 0 489900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5319
timestamp 1676037725
transform 1 0 490452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5321
timestamp 1676037725
transform 1 0 490636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5333
timestamp 1676037725
transform 1 0 491740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5345
timestamp 1676037725
transform 1 0 492844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5357
timestamp 1676037725
transform 1 0 493948 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5369
timestamp 1676037725
transform 1 0 495052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5375
timestamp 1676037725
transform 1 0 495604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5377
timestamp 1676037725
transform 1 0 495788 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5383
timestamp 1676037725
transform 1 0 496340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5395
timestamp 1676037725
transform 1 0 497444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5407
timestamp 1676037725
transform 1 0 498548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5419
timestamp 1676037725
transform 1 0 499652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5431
timestamp 1676037725
transform 1 0 500756 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5433
timestamp 1676037725
transform 1 0 500940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5445
timestamp 1676037725
transform 1 0 502044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5457
timestamp 1676037725
transform 1 0 503148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5469
timestamp 1676037725
transform 1 0 504252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5481
timestamp 1676037725
transform 1 0 505356 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5487
timestamp 1676037725
transform 1 0 505908 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5489
timestamp 1676037725
transform 1 0 506092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5501
timestamp 1676037725
transform 1 0 507196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5513
timestamp 1676037725
transform 1 0 508300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5525
timestamp 1676037725
transform 1 0 509404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5537
timestamp 1676037725
transform 1 0 510508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5543
timestamp 1676037725
transform 1 0 511060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5545
timestamp 1676037725
transform 1 0 511244 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5551
timestamp 1676037725
transform 1 0 511796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5563
timestamp 1676037725
transform 1 0 512900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5575
timestamp 1676037725
transform 1 0 514004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5587
timestamp 1676037725
transform 1 0 515108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5599
timestamp 1676037725
transform 1 0 516212 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5601
timestamp 1676037725
transform 1 0 516396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5613
timestamp 1676037725
transform 1 0 517500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5625
timestamp 1676037725
transform 1 0 518604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5637
timestamp 1676037725
transform 1 0 519708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5649
timestamp 1676037725
transform 1 0 520812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5655
timestamp 1676037725
transform 1 0 521364 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5657
timestamp 1676037725
transform 1 0 521548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5669
timestamp 1676037725
transform 1 0 522652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5681
timestamp 1676037725
transform 1 0 523756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5693
timestamp 1676037725
transform 1 0 524860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5705
timestamp 1676037725
transform 1 0 525964 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5711
timestamp 1676037725
transform 1 0 526516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5713
timestamp 1676037725
transform 1 0 526700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5724
timestamp 1676037725
transform 1 0 527712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5730
timestamp 1676037725
transform 1 0 528264 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5740
timestamp 1676037725
transform 1 0 529184 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5752
timestamp 1676037725
transform 1 0 530288 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5764
timestamp 1676037725
transform 1 0 531392 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5769
timestamp 1676037725
transform 1 0 531852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5781
timestamp 1676037725
transform 1 0 532956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5793
timestamp 1676037725
transform 1 0 534060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5805
timestamp 1676037725
transform 1 0 535164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5817
timestamp 1676037725
transform 1 0 536268 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5823
timestamp 1676037725
transform 1 0 536820 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5825
timestamp 1676037725
transform 1 0 537004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5837
timestamp 1676037725
transform 1 0 538108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5849
timestamp 1676037725
transform 1 0 539212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5861
timestamp 1676037725
transform 1 0 540316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5873
timestamp 1676037725
transform 1 0 541420 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5879
timestamp 1676037725
transform 1 0 541972 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5881
timestamp 1676037725
transform 1 0 542156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5893
timestamp 1676037725
transform 1 0 543260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5905
timestamp 1676037725
transform 1 0 544364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5917
timestamp 1676037725
transform 1 0 545468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5929
timestamp 1676037725
transform 1 0 546572 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5935
timestamp 1676037725
transform 1 0 547124 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5937
timestamp 1676037725
transform 1 0 547308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5949
timestamp 1676037725
transform 1 0 548412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5961
timestamp 1676037725
transform 1 0 549516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5973
timestamp 1676037725
transform 1 0 550620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5985
timestamp 1676037725
transform 1 0 551724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5991
timestamp 1676037725
transform 1 0 552276 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5993
timestamp 1676037725
transform 1 0 552460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6005
timestamp 1676037725
transform 1 0 553564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6017
timestamp 1676037725
transform 1 0 554668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6029
timestamp 1676037725
transform 1 0 555772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6041
timestamp 1676037725
transform 1 0 556876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6047
timestamp 1676037725
transform 1 0 557428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6049
timestamp 1676037725
transform 1 0 557612 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6055
timestamp 1676037725
transform 1 0 558164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6067
timestamp 1676037725
transform 1 0 559268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6079
timestamp 1676037725
transform 1 0 560372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6091
timestamp 1676037725
transform 1 0 561476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6103
timestamp 1676037725
transform 1 0 562580 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6105
timestamp 1676037725
transform 1 0 562764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6117
timestamp 1676037725
transform 1 0 563868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6129
timestamp 1676037725
transform 1 0 564972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6141
timestamp 1676037725
transform 1 0 566076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6153
timestamp 1676037725
transform 1 0 567180 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6159
timestamp 1676037725
transform 1 0 567732 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6161
timestamp 1676037725
transform 1 0 567916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6173
timestamp 1676037725
transform 1 0 569020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6185
timestamp 1676037725
transform 1 0 570124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6197
timestamp 1676037725
transform 1 0 571228 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6209
timestamp 1676037725
transform 1 0 572332 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6215
timestamp 1676037725
transform 1 0 572884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6217
timestamp 1676037725
transform 1 0 573068 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6223
timestamp 1676037725
transform 1 0 573620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6235
timestamp 1676037725
transform 1 0 574724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6247
timestamp 1676037725
transform 1 0 575828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6259
timestamp 1676037725
transform 1 0 576932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6271
timestamp 1676037725
transform 1 0 578036 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6273
timestamp 1676037725
transform 1 0 578220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6285
timestamp 1676037725
transform 1 0 579324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6297
timestamp 1676037725
transform 1 0 580428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6309
timestamp 1676037725
transform 1 0 581532 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6321
timestamp 1676037725
transform 1 0 582636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6327
timestamp 1676037725
transform 1 0 583188 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6329
timestamp 1676037725
transform 1 0 583372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6341
timestamp 1676037725
transform 1 0 584476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6353
timestamp 1676037725
transform 1 0 585580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6365
timestamp 1676037725
transform 1 0 586684 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6377
timestamp 1676037725
transform 1 0 587788 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6383
timestamp 1676037725
transform 1 0 588340 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6385
timestamp 1676037725
transform 1 0 588524 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6391
timestamp 1676037725
transform 1 0 589076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6403
timestamp 1676037725
transform 1 0 590180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6415
timestamp 1676037725
transform 1 0 591284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6427
timestamp 1676037725
transform 1 0 592388 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6439
timestamp 1676037725
transform 1 0 593492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6441
timestamp 1676037725
transform 1 0 593676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6453
timestamp 1676037725
transform 1 0 594780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6465
timestamp 1676037725
transform 1 0 595884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6477
timestamp 1676037725
transform 1 0 596988 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6489
timestamp 1676037725
transform 1 0 598092 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6495
timestamp 1676037725
transform 1 0 598644 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6497
timestamp 1676037725
transform 1 0 598828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6509
timestamp 1676037725
transform 1 0 599932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6521
timestamp 1676037725
transform 1 0 601036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6533
timestamp 1676037725
transform 1 0 602140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6545
timestamp 1676037725
transform 1 0 603244 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6551
timestamp 1676037725
transform 1 0 603796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6553
timestamp 1676037725
transform 1 0 603980 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6559
timestamp 1676037725
transform 1 0 604532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6571
timestamp 1676037725
transform 1 0 605636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6583
timestamp 1676037725
transform 1 0 606740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6595
timestamp 1676037725
transform 1 0 607844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6607
timestamp 1676037725
transform 1 0 608948 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6609
timestamp 1676037725
transform 1 0 609132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6621
timestamp 1676037725
transform 1 0 610236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6633
timestamp 1676037725
transform 1 0 611340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6645
timestamp 1676037725
transform 1 0 612444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6657
timestamp 1676037725
transform 1 0 613548 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6663
timestamp 1676037725
transform 1 0 614100 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6665
timestamp 1676037725
transform 1 0 614284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6677
timestamp 1676037725
transform 1 0 615388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6689
timestamp 1676037725
transform 1 0 616492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6701
timestamp 1676037725
transform 1 0 617596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6713
timestamp 1676037725
transform 1 0 618700 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6719
timestamp 1676037725
transform 1 0 619252 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6721
timestamp 1676037725
transform 1 0 619436 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6727
timestamp 1676037725
transform 1 0 619988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6739
timestamp 1676037725
transform 1 0 621092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6751
timestamp 1676037725
transform 1 0 622196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6763
timestamp 1676037725
transform 1 0 623300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6775
timestamp 1676037725
transform 1 0 624404 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6777
timestamp 1676037725
transform 1 0 624588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6789
timestamp 1676037725
transform 1 0 625692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6801
timestamp 1676037725
transform 1 0 626796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6813
timestamp 1676037725
transform 1 0 627900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6825
timestamp 1676037725
transform 1 0 629004 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6831
timestamp 1676037725
transform 1 0 629556 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6833
timestamp 1676037725
transform 1 0 629740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6845
timestamp 1676037725
transform 1 0 630844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6857
timestamp 1676037725
transform 1 0 631948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6869
timestamp 1676037725
transform 1 0 633052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6881
timestamp 1676037725
transform 1 0 634156 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6887
timestamp 1676037725
transform 1 0 634708 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6889
timestamp 1676037725
transform 1 0 634892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6901
timestamp 1676037725
transform 1 0 635996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6913
timestamp 1676037725
transform 1 0 637100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6925
timestamp 1676037725
transform 1 0 638204 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6937
timestamp 1676037725
transform 1 0 639308 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6943
timestamp 1676037725
transform 1 0 639860 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6945
timestamp 1676037725
transform 1 0 640044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6957
timestamp 1676037725
transform 1 0 641148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6969
timestamp 1676037725
transform 1 0 642252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6981
timestamp 1676037725
transform 1 0 643356 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6993
timestamp 1676037725
transform 1 0 644460 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6999
timestamp 1676037725
transform 1 0 645012 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7001
timestamp 1676037725
transform 1 0 645196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7013
timestamp 1676037725
transform 1 0 646300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7025
timestamp 1676037725
transform 1 0 647404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7037
timestamp 1676037725
transform 1 0 648508 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_7049
timestamp 1676037725
transform 1 0 649612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7055
timestamp 1676037725
transform 1 0 650164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7057
timestamp 1676037725
transform 1 0 650348 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7063
timestamp 1676037725
transform 1 0 650900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7075
timestamp 1676037725
transform 1 0 652004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7087
timestamp 1676037725
transform 1 0 653108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7099
timestamp 1676037725
transform 1 0 654212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7111
timestamp 1676037725
transform 1 0 655316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7113
timestamp 1676037725
transform 1 0 655500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7125
timestamp 1676037725
transform 1 0 656604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7137
timestamp 1676037725
transform 1 0 657708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7149
timestamp 1676037725
transform 1 0 658812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_7161
timestamp 1676037725
transform 1 0 659916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7167
timestamp 1676037725
transform 1 0 660468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7169
timestamp 1676037725
transform 1 0 660652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7181
timestamp 1676037725
transform 1 0 661756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7193
timestamp 1676037725
transform 1 0 662860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7205
timestamp 1676037725
transform 1 0 663964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_7217
timestamp 1676037725
transform 1 0 665068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7223
timestamp 1676037725
transform 1 0 665620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7225
timestamp 1676037725
transform 1 0 665804 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7231
timestamp 1676037725
transform 1 0 666356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7243
timestamp 1676037725
transform 1 0 667460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7255
timestamp 1676037725
transform 1 0 668564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7267
timestamp 1676037725
transform 1 0 669668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7279
timestamp 1676037725
transform 1 0 670772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7281
timestamp 1676037725
transform 1 0 670956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7293
timestamp 1676037725
transform 1 0 672060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7305
timestamp 1676037725
transform 1 0 673164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7317
timestamp 1676037725
transform 1 0 674268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_7329
timestamp 1676037725
transform 1 0 675372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7335
timestamp 1676037725
transform 1 0 675924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7337
timestamp 1676037725
transform 1 0 676108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7349
timestamp 1676037725
transform 1 0 677212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7361
timestamp 1676037725
transform 1 0 678316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7373
timestamp 1676037725
transform 1 0 679420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_7385
timestamp 1676037725
transform 1 0 680524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7391
timestamp 1676037725
transform 1 0 681076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7393
timestamp 1676037725
transform 1 0 681260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_7399
timestamp 1676037725
transform 1 0 681812 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1676037725
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1676037725
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1676037725
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1676037725
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1676037725
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1676037725
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1676037725
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1676037725
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1676037725
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1676037725
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1676037725
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1676037725
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1676037725
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1676037725
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1676037725
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1676037725
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1676037725
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1676037725
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1676037725
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1676037725
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1676037725
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1676037725
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1676037725
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1676037725
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1676037725
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1676037725
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1676037725
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1676037725
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1676037725
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1676037725
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1676037725
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1676037725
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1676037725
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1676037725
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1676037725
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1676037725
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1676037725
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1676037725
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1676037725
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1676037725
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1676037725
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1676037725
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1676037725
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1676037725
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1676037725
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1676037725
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1676037725
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1676037725
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1676037725
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1676037725
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1676037725
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1676037725
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1676037725
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1676037725
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1676037725
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1676037725
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1676037725
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1676037725
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1676037725
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1676037725
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1676037725
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1676037725
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1676037725
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1676037725
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1676037725
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1676037725
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1676037725
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1676037725
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1676037725
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1185
timestamp 1676037725
transform 1 0 110124 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1197
timestamp 1676037725
transform 1 0 111228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1676037725
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1676037725
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1217
timestamp 1676037725
transform 1 0 113068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1229
timestamp 1676037725
transform 1 0 114172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1241
timestamp 1676037725
transform 1 0 115276 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1253
timestamp 1676037725
transform 1 0 116380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1259
timestamp 1676037725
transform 1 0 116932 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1261
timestamp 1676037725
transform 1 0 117116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1273
timestamp 1676037725
transform 1 0 118220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1285
timestamp 1676037725
transform 1 0 119324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1297
timestamp 1676037725
transform 1 0 120428 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1309
timestamp 1676037725
transform 1 0 121532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1315
timestamp 1676037725
transform 1 0 122084 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1317
timestamp 1676037725
transform 1 0 122268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1329
timestamp 1676037725
transform 1 0 123372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1341
timestamp 1676037725
transform 1 0 124476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1353
timestamp 1676037725
transform 1 0 125580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1365
timestamp 1676037725
transform 1 0 126684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1371
timestamp 1676037725
transform 1 0 127236 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1373
timestamp 1676037725
transform 1 0 127420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1385
timestamp 1676037725
transform 1 0 128524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1397
timestamp 1676037725
transform 1 0 129628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1409
timestamp 1676037725
transform 1 0 130732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1421
timestamp 1676037725
transform 1 0 131836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1427
timestamp 1676037725
transform 1 0 132388 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1429
timestamp 1676037725
transform 1 0 132572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1441
timestamp 1676037725
transform 1 0 133676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1453
timestamp 1676037725
transform 1 0 134780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1465
timestamp 1676037725
transform 1 0 135884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1477
timestamp 1676037725
transform 1 0 136988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1483
timestamp 1676037725
transform 1 0 137540 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1485
timestamp 1676037725
transform 1 0 137724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1497
timestamp 1676037725
transform 1 0 138828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1509
timestamp 1676037725
transform 1 0 139932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1521
timestamp 1676037725
transform 1 0 141036 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1533
timestamp 1676037725
transform 1 0 142140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1539
timestamp 1676037725
transform 1 0 142692 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1541
timestamp 1676037725
transform 1 0 142876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1553
timestamp 1676037725
transform 1 0 143980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1565
timestamp 1676037725
transform 1 0 145084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1577
timestamp 1676037725
transform 1 0 146188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1589
timestamp 1676037725
transform 1 0 147292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1595
timestamp 1676037725
transform 1 0 147844 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1597
timestamp 1676037725
transform 1 0 148028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1609
timestamp 1676037725
transform 1 0 149132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1621
timestamp 1676037725
transform 1 0 150236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1633
timestamp 1676037725
transform 1 0 151340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1645
timestamp 1676037725
transform 1 0 152444 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1651
timestamp 1676037725
transform 1 0 152996 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1653
timestamp 1676037725
transform 1 0 153180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1665
timestamp 1676037725
transform 1 0 154284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1677
timestamp 1676037725
transform 1 0 155388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1689
timestamp 1676037725
transform 1 0 156492 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1701
timestamp 1676037725
transform 1 0 157596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1707
timestamp 1676037725
transform 1 0 158148 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1709
timestamp 1676037725
transform 1 0 158332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1721
timestamp 1676037725
transform 1 0 159436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1733
timestamp 1676037725
transform 1 0 160540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1745
timestamp 1676037725
transform 1 0 161644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1757
timestamp 1676037725
transform 1 0 162748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1763
timestamp 1676037725
transform 1 0 163300 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1765
timestamp 1676037725
transform 1 0 163484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1777
timestamp 1676037725
transform 1 0 164588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1789
timestamp 1676037725
transform 1 0 165692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1801
timestamp 1676037725
transform 1 0 166796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1813
timestamp 1676037725
transform 1 0 167900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1819
timestamp 1676037725
transform 1 0 168452 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1821
timestamp 1676037725
transform 1 0 168636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1833
timestamp 1676037725
transform 1 0 169740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1845
timestamp 1676037725
transform 1 0 170844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1857
timestamp 1676037725
transform 1 0 171948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1869
timestamp 1676037725
transform 1 0 173052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1875
timestamp 1676037725
transform 1 0 173604 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1877
timestamp 1676037725
transform 1 0 173788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1889
timestamp 1676037725
transform 1 0 174892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1901
timestamp 1676037725
transform 1 0 175996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1913
timestamp 1676037725
transform 1 0 177100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1925
timestamp 1676037725
transform 1 0 178204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1931
timestamp 1676037725
transform 1 0 178756 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1933
timestamp 1676037725
transform 1 0 178940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1945
timestamp 1676037725
transform 1 0 180044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1957
timestamp 1676037725
transform 1 0 181148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1969
timestamp 1676037725
transform 1 0 182252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1981
timestamp 1676037725
transform 1 0 183356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1987
timestamp 1676037725
transform 1 0 183908 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1989
timestamp 1676037725
transform 1 0 184092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2001
timestamp 1676037725
transform 1 0 185196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2013
timestamp 1676037725
transform 1 0 186300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2025
timestamp 1676037725
transform 1 0 187404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2037
timestamp 1676037725
transform 1 0 188508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2043
timestamp 1676037725
transform 1 0 189060 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2045
timestamp 1676037725
transform 1 0 189244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2057
timestamp 1676037725
transform 1 0 190348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2069
timestamp 1676037725
transform 1 0 191452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2081
timestamp 1676037725
transform 1 0 192556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2093
timestamp 1676037725
transform 1 0 193660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2099
timestamp 1676037725
transform 1 0 194212 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2101
timestamp 1676037725
transform 1 0 194396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2113
timestamp 1676037725
transform 1 0 195500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2125
timestamp 1676037725
transform 1 0 196604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2137
timestamp 1676037725
transform 1 0 197708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2149
timestamp 1676037725
transform 1 0 198812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2155
timestamp 1676037725
transform 1 0 199364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2157
timestamp 1676037725
transform 1 0 199548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2169
timestamp 1676037725
transform 1 0 200652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2181
timestamp 1676037725
transform 1 0 201756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2193
timestamp 1676037725
transform 1 0 202860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2205
timestamp 1676037725
transform 1 0 203964 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2211
timestamp 1676037725
transform 1 0 204516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2213
timestamp 1676037725
transform 1 0 204700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2225
timestamp 1676037725
transform 1 0 205804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2237
timestamp 1676037725
transform 1 0 206908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2249
timestamp 1676037725
transform 1 0 208012 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2261
timestamp 1676037725
transform 1 0 209116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2267
timestamp 1676037725
transform 1 0 209668 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2269
timestamp 1676037725
transform 1 0 209852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2281
timestamp 1676037725
transform 1 0 210956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2293
timestamp 1676037725
transform 1 0 212060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2305
timestamp 1676037725
transform 1 0 213164 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2317
timestamp 1676037725
transform 1 0 214268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2323
timestamp 1676037725
transform 1 0 214820 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2325
timestamp 1676037725
transform 1 0 215004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2337
timestamp 1676037725
transform 1 0 216108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2349
timestamp 1676037725
transform 1 0 217212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2361
timestamp 1676037725
transform 1 0 218316 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2373
timestamp 1676037725
transform 1 0 219420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2379
timestamp 1676037725
transform 1 0 219972 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2381
timestamp 1676037725
transform 1 0 220156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2393
timestamp 1676037725
transform 1 0 221260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2405
timestamp 1676037725
transform 1 0 222364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2417
timestamp 1676037725
transform 1 0 223468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2429
timestamp 1676037725
transform 1 0 224572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2435
timestamp 1676037725
transform 1 0 225124 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2437
timestamp 1676037725
transform 1 0 225308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2449
timestamp 1676037725
transform 1 0 226412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2461
timestamp 1676037725
transform 1 0 227516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2473
timestamp 1676037725
transform 1 0 228620 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2485
timestamp 1676037725
transform 1 0 229724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2491
timestamp 1676037725
transform 1 0 230276 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2493
timestamp 1676037725
transform 1 0 230460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2505
timestamp 1676037725
transform 1 0 231564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2517
timestamp 1676037725
transform 1 0 232668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2529
timestamp 1676037725
transform 1 0 233772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2541
timestamp 1676037725
transform 1 0 234876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2547
timestamp 1676037725
transform 1 0 235428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2549
timestamp 1676037725
transform 1 0 235612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2561
timestamp 1676037725
transform 1 0 236716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2573
timestamp 1676037725
transform 1 0 237820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2585
timestamp 1676037725
transform 1 0 238924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2597
timestamp 1676037725
transform 1 0 240028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2603
timestamp 1676037725
transform 1 0 240580 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2605
timestamp 1676037725
transform 1 0 240764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2617
timestamp 1676037725
transform 1 0 241868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2629
timestamp 1676037725
transform 1 0 242972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2641
timestamp 1676037725
transform 1 0 244076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2653
timestamp 1676037725
transform 1 0 245180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2659
timestamp 1676037725
transform 1 0 245732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2661
timestamp 1676037725
transform 1 0 245916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2673
timestamp 1676037725
transform 1 0 247020 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2685
timestamp 1676037725
transform 1 0 248124 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2693
timestamp 1676037725
transform 1 0 248860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_2705
timestamp 1676037725
transform 1 0 249964 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_2713
timestamp 1676037725
transform 1 0 250700 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2717
timestamp 1676037725
transform 1 0 251068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2729
timestamp 1676037725
transform 1 0 252172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2741
timestamp 1676037725
transform 1 0 253276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2753
timestamp 1676037725
transform 1 0 254380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2765
timestamp 1676037725
transform 1 0 255484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2771
timestamp 1676037725
transform 1 0 256036 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2773
timestamp 1676037725
transform 1 0 256220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2785
timestamp 1676037725
transform 1 0 257324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2797
timestamp 1676037725
transform 1 0 258428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2809
timestamp 1676037725
transform 1 0 259532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2821
timestamp 1676037725
transform 1 0 260636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2827
timestamp 1676037725
transform 1 0 261188 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2829
timestamp 1676037725
transform 1 0 261372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2841
timestamp 1676037725
transform 1 0 262476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2853
timestamp 1676037725
transform 1 0 263580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2865
timestamp 1676037725
transform 1 0 264684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2877
timestamp 1676037725
transform 1 0 265788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2883
timestamp 1676037725
transform 1 0 266340 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2885
timestamp 1676037725
transform 1 0 266524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2897
timestamp 1676037725
transform 1 0 267628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2909
timestamp 1676037725
transform 1 0 268732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2921
timestamp 1676037725
transform 1 0 269836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2933
timestamp 1676037725
transform 1 0 270940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2939
timestamp 1676037725
transform 1 0 271492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2941
timestamp 1676037725
transform 1 0 271676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2953
timestamp 1676037725
transform 1 0 272780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2965
timestamp 1676037725
transform 1 0 273884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2977
timestamp 1676037725
transform 1 0 274988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2989
timestamp 1676037725
transform 1 0 276092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2995
timestamp 1676037725
transform 1 0 276644 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2997
timestamp 1676037725
transform 1 0 276828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3009
timestamp 1676037725
transform 1 0 277932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3021
timestamp 1676037725
transform 1 0 279036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3033
timestamp 1676037725
transform 1 0 280140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3045
timestamp 1676037725
transform 1 0 281244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3051
timestamp 1676037725
transform 1 0 281796 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3053
timestamp 1676037725
transform 1 0 281980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3065
timestamp 1676037725
transform 1 0 283084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3077
timestamp 1676037725
transform 1 0 284188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3089
timestamp 1676037725
transform 1 0 285292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3101
timestamp 1676037725
transform 1 0 286396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3107
timestamp 1676037725
transform 1 0 286948 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3109
timestamp 1676037725
transform 1 0 287132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3121
timestamp 1676037725
transform 1 0 288236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3133
timestamp 1676037725
transform 1 0 289340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3145
timestamp 1676037725
transform 1 0 290444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3157
timestamp 1676037725
transform 1 0 291548 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3163
timestamp 1676037725
transform 1 0 292100 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3165
timestamp 1676037725
transform 1 0 292284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3177
timestamp 1676037725
transform 1 0 293388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3189
timestamp 1676037725
transform 1 0 294492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3201
timestamp 1676037725
transform 1 0 295596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3213
timestamp 1676037725
transform 1 0 296700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3219
timestamp 1676037725
transform 1 0 297252 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3221
timestamp 1676037725
transform 1 0 297436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3233
timestamp 1676037725
transform 1 0 298540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3245
timestamp 1676037725
transform 1 0 299644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3257
timestamp 1676037725
transform 1 0 300748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3269
timestamp 1676037725
transform 1 0 301852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3275
timestamp 1676037725
transform 1 0 302404 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3277
timestamp 1676037725
transform 1 0 302588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3289
timestamp 1676037725
transform 1 0 303692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3301
timestamp 1676037725
transform 1 0 304796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3313
timestamp 1676037725
transform 1 0 305900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3325
timestamp 1676037725
transform 1 0 307004 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3331
timestamp 1676037725
transform 1 0 307556 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3333
timestamp 1676037725
transform 1 0 307740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3345
timestamp 1676037725
transform 1 0 308844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3357
timestamp 1676037725
transform 1 0 309948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3369
timestamp 1676037725
transform 1 0 311052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3381
timestamp 1676037725
transform 1 0 312156 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3387
timestamp 1676037725
transform 1 0 312708 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3389
timestamp 1676037725
transform 1 0 312892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3401
timestamp 1676037725
transform 1 0 313996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3413
timestamp 1676037725
transform 1 0 315100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3425
timestamp 1676037725
transform 1 0 316204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3437
timestamp 1676037725
transform 1 0 317308 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3443
timestamp 1676037725
transform 1 0 317860 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3445
timestamp 1676037725
transform 1 0 318044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3457
timestamp 1676037725
transform 1 0 319148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3469
timestamp 1676037725
transform 1 0 320252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3481
timestamp 1676037725
transform 1 0 321356 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3493
timestamp 1676037725
transform 1 0 322460 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3499
timestamp 1676037725
transform 1 0 323012 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3501
timestamp 1676037725
transform 1 0 323196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3513
timestamp 1676037725
transform 1 0 324300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3525
timestamp 1676037725
transform 1 0 325404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3537
timestamp 1676037725
transform 1 0 326508 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3549
timestamp 1676037725
transform 1 0 327612 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3555
timestamp 1676037725
transform 1 0 328164 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3557
timestamp 1676037725
transform 1 0 328348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3569
timestamp 1676037725
transform 1 0 329452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3581
timestamp 1676037725
transform 1 0 330556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3593
timestamp 1676037725
transform 1 0 331660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3605
timestamp 1676037725
transform 1 0 332764 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3611
timestamp 1676037725
transform 1 0 333316 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3613
timestamp 1676037725
transform 1 0 333500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3625
timestamp 1676037725
transform 1 0 334604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3637
timestamp 1676037725
transform 1 0 335708 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3641
timestamp 1676037725
transform 1 0 336076 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3644
timestamp 1676037725
transform 1 0 336352 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3656
timestamp 1676037725
transform 1 0 337456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3659
timestamp 1676037725
transform 1 0 337732 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3667
timestamp 1676037725
transform 1 0 338468 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3669
timestamp 1676037725
transform 1 0 338652 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3673
timestamp 1676037725
transform 1 0 339020 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3683
timestamp 1676037725
transform 1 0 339940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3695
timestamp 1676037725
transform 1 0 341044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3707
timestamp 1676037725
transform 1 0 342148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3719
timestamp 1676037725
transform 1 0 343252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3723
timestamp 1676037725
transform 1 0 343620 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3725
timestamp 1676037725
transform 1 0 343804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3737
timestamp 1676037725
transform 1 0 344908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3749
timestamp 1676037725
transform 1 0 346012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3761
timestamp 1676037725
transform 1 0 347116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3773
timestamp 1676037725
transform 1 0 348220 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3779
timestamp 1676037725
transform 1 0 348772 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3781
timestamp 1676037725
transform 1 0 348956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3793
timestamp 1676037725
transform 1 0 350060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3805
timestamp 1676037725
transform 1 0 351164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3817
timestamp 1676037725
transform 1 0 352268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3829
timestamp 1676037725
transform 1 0 353372 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3835
timestamp 1676037725
transform 1 0 353924 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3837
timestamp 1676037725
transform 1 0 354108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3849
timestamp 1676037725
transform 1 0 355212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3861
timestamp 1676037725
transform 1 0 356316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3873
timestamp 1676037725
transform 1 0 357420 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3885
timestamp 1676037725
transform 1 0 358524 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3891
timestamp 1676037725
transform 1 0 359076 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3893
timestamp 1676037725
transform 1 0 359260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3905
timestamp 1676037725
transform 1 0 360364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3917
timestamp 1676037725
transform 1 0 361468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3929
timestamp 1676037725
transform 1 0 362572 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3941
timestamp 1676037725
transform 1 0 363676 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3947
timestamp 1676037725
transform 1 0 364228 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3949
timestamp 1676037725
transform 1 0 364412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3961
timestamp 1676037725
transform 1 0 365516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3973
timestamp 1676037725
transform 1 0 366620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3985
timestamp 1676037725
transform 1 0 367724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3997
timestamp 1676037725
transform 1 0 368828 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4003
timestamp 1676037725
transform 1 0 369380 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4005
timestamp 1676037725
transform 1 0 369564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4017
timestamp 1676037725
transform 1 0 370668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4029
timestamp 1676037725
transform 1 0 371772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4041
timestamp 1676037725
transform 1 0 372876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4053
timestamp 1676037725
transform 1 0 373980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4059
timestamp 1676037725
transform 1 0 374532 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4061
timestamp 1676037725
transform 1 0 374716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4073
timestamp 1676037725
transform 1 0 375820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4085
timestamp 1676037725
transform 1 0 376924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4097
timestamp 1676037725
transform 1 0 378028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4109
timestamp 1676037725
transform 1 0 379132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4115
timestamp 1676037725
transform 1 0 379684 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4117
timestamp 1676037725
transform 1 0 379868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4129
timestamp 1676037725
transform 1 0 380972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4141
timestamp 1676037725
transform 1 0 382076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4153
timestamp 1676037725
transform 1 0 383180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4165
timestamp 1676037725
transform 1 0 384284 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4171
timestamp 1676037725
transform 1 0 384836 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4173
timestamp 1676037725
transform 1 0 385020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4185
timestamp 1676037725
transform 1 0 386124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4197
timestamp 1676037725
transform 1 0 387228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4209
timestamp 1676037725
transform 1 0 388332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4221
timestamp 1676037725
transform 1 0 389436 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4227
timestamp 1676037725
transform 1 0 389988 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4229
timestamp 1676037725
transform 1 0 390172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4241
timestamp 1676037725
transform 1 0 391276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4253
timestamp 1676037725
transform 1 0 392380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4265
timestamp 1676037725
transform 1 0 393484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4277
timestamp 1676037725
transform 1 0 394588 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4283
timestamp 1676037725
transform 1 0 395140 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4285
timestamp 1676037725
transform 1 0 395324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4297
timestamp 1676037725
transform 1 0 396428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4309
timestamp 1676037725
transform 1 0 397532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4321
timestamp 1676037725
transform 1 0 398636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4333
timestamp 1676037725
transform 1 0 399740 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4339
timestamp 1676037725
transform 1 0 400292 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4341
timestamp 1676037725
transform 1 0 400476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4353
timestamp 1676037725
transform 1 0 401580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4365
timestamp 1676037725
transform 1 0 402684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4377
timestamp 1676037725
transform 1 0 403788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4389
timestamp 1676037725
transform 1 0 404892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4395
timestamp 1676037725
transform 1 0 405444 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4397
timestamp 1676037725
transform 1 0 405628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4409
timestamp 1676037725
transform 1 0 406732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4421
timestamp 1676037725
transform 1 0 407836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4433
timestamp 1676037725
transform 1 0 408940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4445
timestamp 1676037725
transform 1 0 410044 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4451
timestamp 1676037725
transform 1 0 410596 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4453
timestamp 1676037725
transform 1 0 410780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4465
timestamp 1676037725
transform 1 0 411884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4477
timestamp 1676037725
transform 1 0 412988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4489
timestamp 1676037725
transform 1 0 414092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4501
timestamp 1676037725
transform 1 0 415196 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4507
timestamp 1676037725
transform 1 0 415748 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4509
timestamp 1676037725
transform 1 0 415932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4521
timestamp 1676037725
transform 1 0 417036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4533
timestamp 1676037725
transform 1 0 418140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4545
timestamp 1676037725
transform 1 0 419244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4557
timestamp 1676037725
transform 1 0 420348 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4563
timestamp 1676037725
transform 1 0 420900 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4565
timestamp 1676037725
transform 1 0 421084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4577
timestamp 1676037725
transform 1 0 422188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4589
timestamp 1676037725
transform 1 0 423292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4601
timestamp 1676037725
transform 1 0 424396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4613
timestamp 1676037725
transform 1 0 425500 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4619
timestamp 1676037725
transform 1 0 426052 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4621
timestamp 1676037725
transform 1 0 426236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4633
timestamp 1676037725
transform 1 0 427340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4645
timestamp 1676037725
transform 1 0 428444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4657
timestamp 1676037725
transform 1 0 429548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4669
timestamp 1676037725
transform 1 0 430652 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4675
timestamp 1676037725
transform 1 0 431204 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4677
timestamp 1676037725
transform 1 0 431388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_4689
timestamp 1676037725
transform 1 0 432492 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_4693
timestamp 1676037725
transform 1 0 432860 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_4699
timestamp 1676037725
transform 1 0 433412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_4705
timestamp 1676037725
transform 1 0 433964 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4711
timestamp 1676037725
transform 1 0 434516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_4723
timestamp 1676037725
transform 1 0 435620 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4731
timestamp 1676037725
transform 1 0 436356 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4733
timestamp 1676037725
transform 1 0 436540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4745
timestamp 1676037725
transform 1 0 437644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4757
timestamp 1676037725
transform 1 0 438748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4769
timestamp 1676037725
transform 1 0 439852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4781
timestamp 1676037725
transform 1 0 440956 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4787
timestamp 1676037725
transform 1 0 441508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4789
timestamp 1676037725
transform 1 0 441692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4801
timestamp 1676037725
transform 1 0 442796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4813
timestamp 1676037725
transform 1 0 443900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4825
timestamp 1676037725
transform 1 0 445004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4837
timestamp 1676037725
transform 1 0 446108 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4843
timestamp 1676037725
transform 1 0 446660 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4845
timestamp 1676037725
transform 1 0 446844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4857
timestamp 1676037725
transform 1 0 447948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4869
timestamp 1676037725
transform 1 0 449052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4881
timestamp 1676037725
transform 1 0 450156 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4893
timestamp 1676037725
transform 1 0 451260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4899
timestamp 1676037725
transform 1 0 451812 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4901
timestamp 1676037725
transform 1 0 451996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4913
timestamp 1676037725
transform 1 0 453100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4925
timestamp 1676037725
transform 1 0 454204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4937
timestamp 1676037725
transform 1 0 455308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4949
timestamp 1676037725
transform 1 0 456412 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4955
timestamp 1676037725
transform 1 0 456964 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4957
timestamp 1676037725
transform 1 0 457148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4969
timestamp 1676037725
transform 1 0 458252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4981
timestamp 1676037725
transform 1 0 459356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4993
timestamp 1676037725
transform 1 0 460460 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5005
timestamp 1676037725
transform 1 0 461564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5011
timestamp 1676037725
transform 1 0 462116 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5013
timestamp 1676037725
transform 1 0 462300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5025
timestamp 1676037725
transform 1 0 463404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5037
timestamp 1676037725
transform 1 0 464508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5049
timestamp 1676037725
transform 1 0 465612 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5061
timestamp 1676037725
transform 1 0 466716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5067
timestamp 1676037725
transform 1 0 467268 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5069
timestamp 1676037725
transform 1 0 467452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5081
timestamp 1676037725
transform 1 0 468556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5093
timestamp 1676037725
transform 1 0 469660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5105
timestamp 1676037725
transform 1 0 470764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5117
timestamp 1676037725
transform 1 0 471868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5123
timestamp 1676037725
transform 1 0 472420 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5125
timestamp 1676037725
transform 1 0 472604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5137
timestamp 1676037725
transform 1 0 473708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5149
timestamp 1676037725
transform 1 0 474812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5161
timestamp 1676037725
transform 1 0 475916 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5173
timestamp 1676037725
transform 1 0 477020 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5179
timestamp 1676037725
transform 1 0 477572 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5181
timestamp 1676037725
transform 1 0 477756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5193
timestamp 1676037725
transform 1 0 478860 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5205
timestamp 1676037725
transform 1 0 479964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5217
timestamp 1676037725
transform 1 0 481068 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5229
timestamp 1676037725
transform 1 0 482172 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5235
timestamp 1676037725
transform 1 0 482724 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5237
timestamp 1676037725
transform 1 0 482908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5249
timestamp 1676037725
transform 1 0 484012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5261
timestamp 1676037725
transform 1 0 485116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5273
timestamp 1676037725
transform 1 0 486220 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5285
timestamp 1676037725
transform 1 0 487324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5291
timestamp 1676037725
transform 1 0 487876 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5293
timestamp 1676037725
transform 1 0 488060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5305
timestamp 1676037725
transform 1 0 489164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5317
timestamp 1676037725
transform 1 0 490268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5329
timestamp 1676037725
transform 1 0 491372 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5341
timestamp 1676037725
transform 1 0 492476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5347
timestamp 1676037725
transform 1 0 493028 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5349
timestamp 1676037725
transform 1 0 493212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5361
timestamp 1676037725
transform 1 0 494316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5373
timestamp 1676037725
transform 1 0 495420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5385
timestamp 1676037725
transform 1 0 496524 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5397
timestamp 1676037725
transform 1 0 497628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5403
timestamp 1676037725
transform 1 0 498180 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5405
timestamp 1676037725
transform 1 0 498364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5417
timestamp 1676037725
transform 1 0 499468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5429
timestamp 1676037725
transform 1 0 500572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5441
timestamp 1676037725
transform 1 0 501676 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5453
timestamp 1676037725
transform 1 0 502780 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5459
timestamp 1676037725
transform 1 0 503332 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5461
timestamp 1676037725
transform 1 0 503516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5473
timestamp 1676037725
transform 1 0 504620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5485
timestamp 1676037725
transform 1 0 505724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5497
timestamp 1676037725
transform 1 0 506828 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5509
timestamp 1676037725
transform 1 0 507932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5515
timestamp 1676037725
transform 1 0 508484 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5517
timestamp 1676037725
transform 1 0 508668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5529
timestamp 1676037725
transform 1 0 509772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5541
timestamp 1676037725
transform 1 0 510876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5553
timestamp 1676037725
transform 1 0 511980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5565
timestamp 1676037725
transform 1 0 513084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5571
timestamp 1676037725
transform 1 0 513636 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5573
timestamp 1676037725
transform 1 0 513820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5585
timestamp 1676037725
transform 1 0 514924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5597
timestamp 1676037725
transform 1 0 516028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5609
timestamp 1676037725
transform 1 0 517132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5621
timestamp 1676037725
transform 1 0 518236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5627
timestamp 1676037725
transform 1 0 518788 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5629
timestamp 1676037725
transform 1 0 518972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5641
timestamp 1676037725
transform 1 0 520076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5653
timestamp 1676037725
transform 1 0 521180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5665
timestamp 1676037725
transform 1 0 522284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5677
timestamp 1676037725
transform 1 0 523388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5683
timestamp 1676037725
transform 1 0 523940 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5685
timestamp 1676037725
transform 1 0 524124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5697
timestamp 1676037725
transform 1 0 525228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_5709
timestamp 1676037725
transform 1 0 526332 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5719
timestamp 1676037725
transform 1 0 527252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_5731
timestamp 1676037725
transform 1 0 528356 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5739
timestamp 1676037725
transform 1 0 529092 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5741
timestamp 1676037725
transform 1 0 529276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5753
timestamp 1676037725
transform 1 0 530380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5765
timestamp 1676037725
transform 1 0 531484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5777
timestamp 1676037725
transform 1 0 532588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5789
timestamp 1676037725
transform 1 0 533692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5795
timestamp 1676037725
transform 1 0 534244 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5797
timestamp 1676037725
transform 1 0 534428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5809
timestamp 1676037725
transform 1 0 535532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5821
timestamp 1676037725
transform 1 0 536636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5833
timestamp 1676037725
transform 1 0 537740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5845
timestamp 1676037725
transform 1 0 538844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5851
timestamp 1676037725
transform 1 0 539396 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5853
timestamp 1676037725
transform 1 0 539580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5865
timestamp 1676037725
transform 1 0 540684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5877
timestamp 1676037725
transform 1 0 541788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5889
timestamp 1676037725
transform 1 0 542892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5901
timestamp 1676037725
transform 1 0 543996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5907
timestamp 1676037725
transform 1 0 544548 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5909
timestamp 1676037725
transform 1 0 544732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5921
timestamp 1676037725
transform 1 0 545836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5933
timestamp 1676037725
transform 1 0 546940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5945
timestamp 1676037725
transform 1 0 548044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5957
timestamp 1676037725
transform 1 0 549148 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5963
timestamp 1676037725
transform 1 0 549700 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5965
timestamp 1676037725
transform 1 0 549884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5977
timestamp 1676037725
transform 1 0 550988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5989
timestamp 1676037725
transform 1 0 552092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6001
timestamp 1676037725
transform 1 0 553196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6013
timestamp 1676037725
transform 1 0 554300 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6019
timestamp 1676037725
transform 1 0 554852 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6021
timestamp 1676037725
transform 1 0 555036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6033
timestamp 1676037725
transform 1 0 556140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6045
timestamp 1676037725
transform 1 0 557244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6057
timestamp 1676037725
transform 1 0 558348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6069
timestamp 1676037725
transform 1 0 559452 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6075
timestamp 1676037725
transform 1 0 560004 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6077
timestamp 1676037725
transform 1 0 560188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6089
timestamp 1676037725
transform 1 0 561292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6101
timestamp 1676037725
transform 1 0 562396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6113
timestamp 1676037725
transform 1 0 563500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6125
timestamp 1676037725
transform 1 0 564604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6131
timestamp 1676037725
transform 1 0 565156 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6133
timestamp 1676037725
transform 1 0 565340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6145
timestamp 1676037725
transform 1 0 566444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6157
timestamp 1676037725
transform 1 0 567548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6169
timestamp 1676037725
transform 1 0 568652 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6181
timestamp 1676037725
transform 1 0 569756 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6187
timestamp 1676037725
transform 1 0 570308 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6189
timestamp 1676037725
transform 1 0 570492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6201
timestamp 1676037725
transform 1 0 571596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6213
timestamp 1676037725
transform 1 0 572700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6225
timestamp 1676037725
transform 1 0 573804 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6237
timestamp 1676037725
transform 1 0 574908 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6243
timestamp 1676037725
transform 1 0 575460 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6245
timestamp 1676037725
transform 1 0 575644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6257
timestamp 1676037725
transform 1 0 576748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6269
timestamp 1676037725
transform 1 0 577852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6281
timestamp 1676037725
transform 1 0 578956 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6293
timestamp 1676037725
transform 1 0 580060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6299
timestamp 1676037725
transform 1 0 580612 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6301
timestamp 1676037725
transform 1 0 580796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6313
timestamp 1676037725
transform 1 0 581900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6325
timestamp 1676037725
transform 1 0 583004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6337
timestamp 1676037725
transform 1 0 584108 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6349
timestamp 1676037725
transform 1 0 585212 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6355
timestamp 1676037725
transform 1 0 585764 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6357
timestamp 1676037725
transform 1 0 585948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6369
timestamp 1676037725
transform 1 0 587052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6381
timestamp 1676037725
transform 1 0 588156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6393
timestamp 1676037725
transform 1 0 589260 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6405
timestamp 1676037725
transform 1 0 590364 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6411
timestamp 1676037725
transform 1 0 590916 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6413
timestamp 1676037725
transform 1 0 591100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6425
timestamp 1676037725
transform 1 0 592204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6437
timestamp 1676037725
transform 1 0 593308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6449
timestamp 1676037725
transform 1 0 594412 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6461
timestamp 1676037725
transform 1 0 595516 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6467
timestamp 1676037725
transform 1 0 596068 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6469
timestamp 1676037725
transform 1 0 596252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6481
timestamp 1676037725
transform 1 0 597356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6493
timestamp 1676037725
transform 1 0 598460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6505
timestamp 1676037725
transform 1 0 599564 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6517
timestamp 1676037725
transform 1 0 600668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6523
timestamp 1676037725
transform 1 0 601220 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6525
timestamp 1676037725
transform 1 0 601404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6537
timestamp 1676037725
transform 1 0 602508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6549
timestamp 1676037725
transform 1 0 603612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6561
timestamp 1676037725
transform 1 0 604716 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6573
timestamp 1676037725
transform 1 0 605820 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6579
timestamp 1676037725
transform 1 0 606372 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6581
timestamp 1676037725
transform 1 0 606556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6593
timestamp 1676037725
transform 1 0 607660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6605
timestamp 1676037725
transform 1 0 608764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6617
timestamp 1676037725
transform 1 0 609868 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6629
timestamp 1676037725
transform 1 0 610972 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6635
timestamp 1676037725
transform 1 0 611524 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6637
timestamp 1676037725
transform 1 0 611708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6649
timestamp 1676037725
transform 1 0 612812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6661
timestamp 1676037725
transform 1 0 613916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6673
timestamp 1676037725
transform 1 0 615020 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6685
timestamp 1676037725
transform 1 0 616124 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6691
timestamp 1676037725
transform 1 0 616676 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6693
timestamp 1676037725
transform 1 0 616860 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6705
timestamp 1676037725
transform 1 0 617964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6717
timestamp 1676037725
transform 1 0 619068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6729
timestamp 1676037725
transform 1 0 620172 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6741
timestamp 1676037725
transform 1 0 621276 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6747
timestamp 1676037725
transform 1 0 621828 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6749
timestamp 1676037725
transform 1 0 622012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6761
timestamp 1676037725
transform 1 0 623116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6773
timestamp 1676037725
transform 1 0 624220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6785
timestamp 1676037725
transform 1 0 625324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6797
timestamp 1676037725
transform 1 0 626428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6803
timestamp 1676037725
transform 1 0 626980 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6805
timestamp 1676037725
transform 1 0 627164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6817
timestamp 1676037725
transform 1 0 628268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6829
timestamp 1676037725
transform 1 0 629372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6841
timestamp 1676037725
transform 1 0 630476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6853
timestamp 1676037725
transform 1 0 631580 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6859
timestamp 1676037725
transform 1 0 632132 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6861
timestamp 1676037725
transform 1 0 632316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6873
timestamp 1676037725
transform 1 0 633420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6885
timestamp 1676037725
transform 1 0 634524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6897
timestamp 1676037725
transform 1 0 635628 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6909
timestamp 1676037725
transform 1 0 636732 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6915
timestamp 1676037725
transform 1 0 637284 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6917
timestamp 1676037725
transform 1 0 637468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6929
timestamp 1676037725
transform 1 0 638572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6941
timestamp 1676037725
transform 1 0 639676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6953
timestamp 1676037725
transform 1 0 640780 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6965
timestamp 1676037725
transform 1 0 641884 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6971
timestamp 1676037725
transform 1 0 642436 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6973
timestamp 1676037725
transform 1 0 642620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6985
timestamp 1676037725
transform 1 0 643724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6997
timestamp 1676037725
transform 1 0 644828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7009
timestamp 1676037725
transform 1 0 645932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7021
timestamp 1676037725
transform 1 0 647036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7027
timestamp 1676037725
transform 1 0 647588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7029
timestamp 1676037725
transform 1 0 647772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7041
timestamp 1676037725
transform 1 0 648876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7053
timestamp 1676037725
transform 1 0 649980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7065
timestamp 1676037725
transform 1 0 651084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7077
timestamp 1676037725
transform 1 0 652188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7083
timestamp 1676037725
transform 1 0 652740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7085
timestamp 1676037725
transform 1 0 652924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7097
timestamp 1676037725
transform 1 0 654028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7109
timestamp 1676037725
transform 1 0 655132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7121
timestamp 1676037725
transform 1 0 656236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7133
timestamp 1676037725
transform 1 0 657340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7139
timestamp 1676037725
transform 1 0 657892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7141
timestamp 1676037725
transform 1 0 658076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7153
timestamp 1676037725
transform 1 0 659180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7165
timestamp 1676037725
transform 1 0 660284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7177
timestamp 1676037725
transform 1 0 661388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7189
timestamp 1676037725
transform 1 0 662492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7195
timestamp 1676037725
transform 1 0 663044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7197
timestamp 1676037725
transform 1 0 663228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7209
timestamp 1676037725
transform 1 0 664332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7221
timestamp 1676037725
transform 1 0 665436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7233
timestamp 1676037725
transform 1 0 666540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7245
timestamp 1676037725
transform 1 0 667644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7251
timestamp 1676037725
transform 1 0 668196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7253
timestamp 1676037725
transform 1 0 668380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7265
timestamp 1676037725
transform 1 0 669484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7277
timestamp 1676037725
transform 1 0 670588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7289
timestamp 1676037725
transform 1 0 671692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7301
timestamp 1676037725
transform 1 0 672796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7307
timestamp 1676037725
transform 1 0 673348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7309
timestamp 1676037725
transform 1 0 673532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7321
timestamp 1676037725
transform 1 0 674636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7333
timestamp 1676037725
transform 1 0 675740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7345
timestamp 1676037725
transform 1 0 676844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7357
timestamp 1676037725
transform 1 0 677948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7363
timestamp 1676037725
transform 1 0 678500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7365
timestamp 1676037725
transform 1 0 678684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7377
timestamp 1676037725
transform 1 0 679788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7389
timestamp 1676037725
transform 1 0 680892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7401
timestamp 1676037725
transform 1 0 681996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1676037725
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1676037725
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1676037725
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1676037725
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1676037725
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1676037725
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1676037725
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1676037725
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1676037725
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1676037725
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1676037725
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1676037725
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1676037725
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1676037725
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1676037725
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1676037725
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1676037725
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1676037725
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1676037725
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1676037725
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1676037725
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1676037725
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1676037725
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1676037725
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1676037725
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1676037725
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1676037725
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1676037725
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1676037725
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1676037725
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1676037725
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1676037725
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1676037725
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1676037725
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1676037725
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1676037725
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1676037725
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1676037725
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1676037725
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1676037725
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1676037725
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1676037725
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1676037725
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1676037725
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1676037725
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1676037725
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1676037725
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1676037725
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1676037725
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1676037725
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1676037725
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1676037725
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1676037725
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1676037725
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1676037725
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1676037725
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1676037725
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1676037725
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1676037725
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1676037725
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1676037725
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1676037725
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1676037725
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1676037725
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1676037725
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1676037725
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1676037725
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1676037725
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1676037725
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1676037725
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1676037725
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1676037725
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1676037725
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1676037725
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1676037725
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1676037725
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1257
timestamp 1676037725
transform 1 0 116748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1269
timestamp 1676037725
transform 1 0 117852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1281
timestamp 1676037725
transform 1 0 118956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1287
timestamp 1676037725
transform 1 0 119508 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1289
timestamp 1676037725
transform 1 0 119692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1301
timestamp 1676037725
transform 1 0 120796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1313
timestamp 1676037725
transform 1 0 121900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1325
timestamp 1676037725
transform 1 0 123004 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1337
timestamp 1676037725
transform 1 0 124108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1343
timestamp 1676037725
transform 1 0 124660 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1345
timestamp 1676037725
transform 1 0 124844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1357
timestamp 1676037725
transform 1 0 125948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1369
timestamp 1676037725
transform 1 0 127052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1381
timestamp 1676037725
transform 1 0 128156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1393
timestamp 1676037725
transform 1 0 129260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1399
timestamp 1676037725
transform 1 0 129812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1401
timestamp 1676037725
transform 1 0 129996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1413
timestamp 1676037725
transform 1 0 131100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1425
timestamp 1676037725
transform 1 0 132204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1437
timestamp 1676037725
transform 1 0 133308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1449
timestamp 1676037725
transform 1 0 134412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1455
timestamp 1676037725
transform 1 0 134964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1457
timestamp 1676037725
transform 1 0 135148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1469
timestamp 1676037725
transform 1 0 136252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1481
timestamp 1676037725
transform 1 0 137356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1493
timestamp 1676037725
transform 1 0 138460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1505
timestamp 1676037725
transform 1 0 139564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1511
timestamp 1676037725
transform 1 0 140116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1513
timestamp 1676037725
transform 1 0 140300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1525
timestamp 1676037725
transform 1 0 141404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1537
timestamp 1676037725
transform 1 0 142508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1549
timestamp 1676037725
transform 1 0 143612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1561
timestamp 1676037725
transform 1 0 144716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1567
timestamp 1676037725
transform 1 0 145268 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1569
timestamp 1676037725
transform 1 0 145452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1581
timestamp 1676037725
transform 1 0 146556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1593
timestamp 1676037725
transform 1 0 147660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1605
timestamp 1676037725
transform 1 0 148764 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1617
timestamp 1676037725
transform 1 0 149868 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1623
timestamp 1676037725
transform 1 0 150420 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1625
timestamp 1676037725
transform 1 0 150604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1637
timestamp 1676037725
transform 1 0 151708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1649
timestamp 1676037725
transform 1 0 152812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1661
timestamp 1676037725
transform 1 0 153916 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1673
timestamp 1676037725
transform 1 0 155020 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1679
timestamp 1676037725
transform 1 0 155572 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1681
timestamp 1676037725
transform 1 0 155756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1693
timestamp 1676037725
transform 1 0 156860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1705
timestamp 1676037725
transform 1 0 157964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1717
timestamp 1676037725
transform 1 0 159068 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1729
timestamp 1676037725
transform 1 0 160172 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1735
timestamp 1676037725
transform 1 0 160724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1737
timestamp 1676037725
transform 1 0 160908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1749
timestamp 1676037725
transform 1 0 162012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1761
timestamp 1676037725
transform 1 0 163116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1773
timestamp 1676037725
transform 1 0 164220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1785
timestamp 1676037725
transform 1 0 165324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1791
timestamp 1676037725
transform 1 0 165876 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1793
timestamp 1676037725
transform 1 0 166060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1805
timestamp 1676037725
transform 1 0 167164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1817
timestamp 1676037725
transform 1 0 168268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1829
timestamp 1676037725
transform 1 0 169372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1841
timestamp 1676037725
transform 1 0 170476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1847
timestamp 1676037725
transform 1 0 171028 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1849
timestamp 1676037725
transform 1 0 171212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1861
timestamp 1676037725
transform 1 0 172316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1873
timestamp 1676037725
transform 1 0 173420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1885
timestamp 1676037725
transform 1 0 174524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1897
timestamp 1676037725
transform 1 0 175628 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1903
timestamp 1676037725
transform 1 0 176180 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1905
timestamp 1676037725
transform 1 0 176364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1917
timestamp 1676037725
transform 1 0 177468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1929
timestamp 1676037725
transform 1 0 178572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1941
timestamp 1676037725
transform 1 0 179676 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1953
timestamp 1676037725
transform 1 0 180780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1959
timestamp 1676037725
transform 1 0 181332 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1961
timestamp 1676037725
transform 1 0 181516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1973
timestamp 1676037725
transform 1 0 182620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1985
timestamp 1676037725
transform 1 0 183724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1997
timestamp 1676037725
transform 1 0 184828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2009
timestamp 1676037725
transform 1 0 185932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2015
timestamp 1676037725
transform 1 0 186484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2017
timestamp 1676037725
transform 1 0 186668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2029
timestamp 1676037725
transform 1 0 187772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2041
timestamp 1676037725
transform 1 0 188876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2053
timestamp 1676037725
transform 1 0 189980 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2065
timestamp 1676037725
transform 1 0 191084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2071
timestamp 1676037725
transform 1 0 191636 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2073
timestamp 1676037725
transform 1 0 191820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2085
timestamp 1676037725
transform 1 0 192924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2097
timestamp 1676037725
transform 1 0 194028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2109
timestamp 1676037725
transform 1 0 195132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2121
timestamp 1676037725
transform 1 0 196236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2127
timestamp 1676037725
transform 1 0 196788 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2129
timestamp 1676037725
transform 1 0 196972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2141
timestamp 1676037725
transform 1 0 198076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2153
timestamp 1676037725
transform 1 0 199180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2165
timestamp 1676037725
transform 1 0 200284 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2177
timestamp 1676037725
transform 1 0 201388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2183
timestamp 1676037725
transform 1 0 201940 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2185
timestamp 1676037725
transform 1 0 202124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2197
timestamp 1676037725
transform 1 0 203228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2209
timestamp 1676037725
transform 1 0 204332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2221
timestamp 1676037725
transform 1 0 205436 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2233
timestamp 1676037725
transform 1 0 206540 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2239
timestamp 1676037725
transform 1 0 207092 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2241
timestamp 1676037725
transform 1 0 207276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2253
timestamp 1676037725
transform 1 0 208380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2265
timestamp 1676037725
transform 1 0 209484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2277
timestamp 1676037725
transform 1 0 210588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2289
timestamp 1676037725
transform 1 0 211692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2295
timestamp 1676037725
transform 1 0 212244 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2297
timestamp 1676037725
transform 1 0 212428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2309
timestamp 1676037725
transform 1 0 213532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2321
timestamp 1676037725
transform 1 0 214636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2333
timestamp 1676037725
transform 1 0 215740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2345
timestamp 1676037725
transform 1 0 216844 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2351
timestamp 1676037725
transform 1 0 217396 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2353
timestamp 1676037725
transform 1 0 217580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2365
timestamp 1676037725
transform 1 0 218684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2377
timestamp 1676037725
transform 1 0 219788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2389
timestamp 1676037725
transform 1 0 220892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2401
timestamp 1676037725
transform 1 0 221996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2407
timestamp 1676037725
transform 1 0 222548 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2409
timestamp 1676037725
transform 1 0 222732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2421
timestamp 1676037725
transform 1 0 223836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2433
timestamp 1676037725
transform 1 0 224940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2445
timestamp 1676037725
transform 1 0 226044 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2457
timestamp 1676037725
transform 1 0 227148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2463
timestamp 1676037725
transform 1 0 227700 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2465
timestamp 1676037725
transform 1 0 227884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2477
timestamp 1676037725
transform 1 0 228988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2489
timestamp 1676037725
transform 1 0 230092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2501
timestamp 1676037725
transform 1 0 231196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2513
timestamp 1676037725
transform 1 0 232300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2519
timestamp 1676037725
transform 1 0 232852 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2521
timestamp 1676037725
transform 1 0 233036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2533
timestamp 1676037725
transform 1 0 234140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2545
timestamp 1676037725
transform 1 0 235244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2557
timestamp 1676037725
transform 1 0 236348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2569
timestamp 1676037725
transform 1 0 237452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2575
timestamp 1676037725
transform 1 0 238004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2577
timestamp 1676037725
transform 1 0 238188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2589
timestamp 1676037725
transform 1 0 239292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2601
timestamp 1676037725
transform 1 0 240396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2613
timestamp 1676037725
transform 1 0 241500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2625
timestamp 1676037725
transform 1 0 242604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2631
timestamp 1676037725
transform 1 0 243156 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2633
timestamp 1676037725
transform 1 0 243340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2645
timestamp 1676037725
transform 1 0 244444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2657
timestamp 1676037725
transform 1 0 245548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2669
timestamp 1676037725
transform 1 0 246652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2681
timestamp 1676037725
transform 1 0 247756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2687
timestamp 1676037725
transform 1 0 248308 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2689
timestamp 1676037725
transform 1 0 248492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2701
timestamp 1676037725
transform 1 0 249596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2713
timestamp 1676037725
transform 1 0 250700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2725
timestamp 1676037725
transform 1 0 251804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2737
timestamp 1676037725
transform 1 0 252908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2743
timestamp 1676037725
transform 1 0 253460 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2745
timestamp 1676037725
transform 1 0 253644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2757
timestamp 1676037725
transform 1 0 254748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2769
timestamp 1676037725
transform 1 0 255852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2781
timestamp 1676037725
transform 1 0 256956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2793
timestamp 1676037725
transform 1 0 258060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2799
timestamp 1676037725
transform 1 0 258612 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2801
timestamp 1676037725
transform 1 0 258796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2813
timestamp 1676037725
transform 1 0 259900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2825
timestamp 1676037725
transform 1 0 261004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2837
timestamp 1676037725
transform 1 0 262108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2849
timestamp 1676037725
transform 1 0 263212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2855
timestamp 1676037725
transform 1 0 263764 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2857
timestamp 1676037725
transform 1 0 263948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2869
timestamp 1676037725
transform 1 0 265052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2881
timestamp 1676037725
transform 1 0 266156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2893
timestamp 1676037725
transform 1 0 267260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2905
timestamp 1676037725
transform 1 0 268364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2911
timestamp 1676037725
transform 1 0 268916 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2913
timestamp 1676037725
transform 1 0 269100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2925
timestamp 1676037725
transform 1 0 270204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2937
timestamp 1676037725
transform 1 0 271308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2949
timestamp 1676037725
transform 1 0 272412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2961
timestamp 1676037725
transform 1 0 273516 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2967
timestamp 1676037725
transform 1 0 274068 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2969
timestamp 1676037725
transform 1 0 274252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2981
timestamp 1676037725
transform 1 0 275356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2993
timestamp 1676037725
transform 1 0 276460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3005
timestamp 1676037725
transform 1 0 277564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3017
timestamp 1676037725
transform 1 0 278668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3023
timestamp 1676037725
transform 1 0 279220 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3025
timestamp 1676037725
transform 1 0 279404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3037
timestamp 1676037725
transform 1 0 280508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3049
timestamp 1676037725
transform 1 0 281612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3061
timestamp 1676037725
transform 1 0 282716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3073
timestamp 1676037725
transform 1 0 283820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3079
timestamp 1676037725
transform 1 0 284372 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3081
timestamp 1676037725
transform 1 0 284556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3093
timestamp 1676037725
transform 1 0 285660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3105
timestamp 1676037725
transform 1 0 286764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3117
timestamp 1676037725
transform 1 0 287868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3129
timestamp 1676037725
transform 1 0 288972 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3135
timestamp 1676037725
transform 1 0 289524 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3137
timestamp 1676037725
transform 1 0 289708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3149
timestamp 1676037725
transform 1 0 290812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3161
timestamp 1676037725
transform 1 0 291916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3173
timestamp 1676037725
transform 1 0 293020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3185
timestamp 1676037725
transform 1 0 294124 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3191
timestamp 1676037725
transform 1 0 294676 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3193
timestamp 1676037725
transform 1 0 294860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3205
timestamp 1676037725
transform 1 0 295964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3217
timestamp 1676037725
transform 1 0 297068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3229
timestamp 1676037725
transform 1 0 298172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3241
timestamp 1676037725
transform 1 0 299276 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3247
timestamp 1676037725
transform 1 0 299828 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3249
timestamp 1676037725
transform 1 0 300012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3261
timestamp 1676037725
transform 1 0 301116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3273
timestamp 1676037725
transform 1 0 302220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3285
timestamp 1676037725
transform 1 0 303324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3297
timestamp 1676037725
transform 1 0 304428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3303
timestamp 1676037725
transform 1 0 304980 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3305
timestamp 1676037725
transform 1 0 305164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3317
timestamp 1676037725
transform 1 0 306268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3329
timestamp 1676037725
transform 1 0 307372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3341
timestamp 1676037725
transform 1 0 308476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3353
timestamp 1676037725
transform 1 0 309580 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3359
timestamp 1676037725
transform 1 0 310132 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3361
timestamp 1676037725
transform 1 0 310316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3373
timestamp 1676037725
transform 1 0 311420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3385
timestamp 1676037725
transform 1 0 312524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3397
timestamp 1676037725
transform 1 0 313628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3409
timestamp 1676037725
transform 1 0 314732 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3415
timestamp 1676037725
transform 1 0 315284 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3417
timestamp 1676037725
transform 1 0 315468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3429
timestamp 1676037725
transform 1 0 316572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3441
timestamp 1676037725
transform 1 0 317676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3453
timestamp 1676037725
transform 1 0 318780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3465
timestamp 1676037725
transform 1 0 319884 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3471
timestamp 1676037725
transform 1 0 320436 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3473
timestamp 1676037725
transform 1 0 320620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3485
timestamp 1676037725
transform 1 0 321724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3497
timestamp 1676037725
transform 1 0 322828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3509
timestamp 1676037725
transform 1 0 323932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3521
timestamp 1676037725
transform 1 0 325036 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3527
timestamp 1676037725
transform 1 0 325588 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3529
timestamp 1676037725
transform 1 0 325772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3541
timestamp 1676037725
transform 1 0 326876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3553
timestamp 1676037725
transform 1 0 327980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3565
timestamp 1676037725
transform 1 0 329084 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3577
timestamp 1676037725
transform 1 0 330188 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3583
timestamp 1676037725
transform 1 0 330740 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3585
timestamp 1676037725
transform 1 0 330924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3597
timestamp 1676037725
transform 1 0 332028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3609
timestamp 1676037725
transform 1 0 333132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3621
timestamp 1676037725
transform 1 0 334236 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3633
timestamp 1676037725
transform 1 0 335340 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3639
timestamp 1676037725
transform 1 0 335892 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3641
timestamp 1676037725
transform 1 0 336076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3653
timestamp 1676037725
transform 1 0 337180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3665
timestamp 1676037725
transform 1 0 338284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3677
timestamp 1676037725
transform 1 0 339388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3689
timestamp 1676037725
transform 1 0 340492 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3695
timestamp 1676037725
transform 1 0 341044 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3697
timestamp 1676037725
transform 1 0 341228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3709
timestamp 1676037725
transform 1 0 342332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3721
timestamp 1676037725
transform 1 0 343436 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3733
timestamp 1676037725
transform 1 0 344540 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3745
timestamp 1676037725
transform 1 0 345644 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3751
timestamp 1676037725
transform 1 0 346196 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3753
timestamp 1676037725
transform 1 0 346380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3765
timestamp 1676037725
transform 1 0 347484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3777
timestamp 1676037725
transform 1 0 348588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3789
timestamp 1676037725
transform 1 0 349692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3801
timestamp 1676037725
transform 1 0 350796 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3807
timestamp 1676037725
transform 1 0 351348 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3809
timestamp 1676037725
transform 1 0 351532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3821
timestamp 1676037725
transform 1 0 352636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3833
timestamp 1676037725
transform 1 0 353740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3845
timestamp 1676037725
transform 1 0 354844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3857
timestamp 1676037725
transform 1 0 355948 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3863
timestamp 1676037725
transform 1 0 356500 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3865
timestamp 1676037725
transform 1 0 356684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3877
timestamp 1676037725
transform 1 0 357788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3889
timestamp 1676037725
transform 1 0 358892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3901
timestamp 1676037725
transform 1 0 359996 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3913
timestamp 1676037725
transform 1 0 361100 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3919
timestamp 1676037725
transform 1 0 361652 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3921
timestamp 1676037725
transform 1 0 361836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3933
timestamp 1676037725
transform 1 0 362940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3945
timestamp 1676037725
transform 1 0 364044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3957
timestamp 1676037725
transform 1 0 365148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3969
timestamp 1676037725
transform 1 0 366252 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3975
timestamp 1676037725
transform 1 0 366804 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3977
timestamp 1676037725
transform 1 0 366988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3989
timestamp 1676037725
transform 1 0 368092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4001
timestamp 1676037725
transform 1 0 369196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4013
timestamp 1676037725
transform 1 0 370300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4025
timestamp 1676037725
transform 1 0 371404 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4031
timestamp 1676037725
transform 1 0 371956 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4033
timestamp 1676037725
transform 1 0 372140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4045
timestamp 1676037725
transform 1 0 373244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4057
timestamp 1676037725
transform 1 0 374348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4069
timestamp 1676037725
transform 1 0 375452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4081
timestamp 1676037725
transform 1 0 376556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4087
timestamp 1676037725
transform 1 0 377108 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4089
timestamp 1676037725
transform 1 0 377292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4101
timestamp 1676037725
transform 1 0 378396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4113
timestamp 1676037725
transform 1 0 379500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4125
timestamp 1676037725
transform 1 0 380604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4137
timestamp 1676037725
transform 1 0 381708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4143
timestamp 1676037725
transform 1 0 382260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4145
timestamp 1676037725
transform 1 0 382444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4157
timestamp 1676037725
transform 1 0 383548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4169
timestamp 1676037725
transform 1 0 384652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4181
timestamp 1676037725
transform 1 0 385756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4193
timestamp 1676037725
transform 1 0 386860 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4199
timestamp 1676037725
transform 1 0 387412 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4201
timestamp 1676037725
transform 1 0 387596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4213
timestamp 1676037725
transform 1 0 388700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4225
timestamp 1676037725
transform 1 0 389804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4237
timestamp 1676037725
transform 1 0 390908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4249
timestamp 1676037725
transform 1 0 392012 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4255
timestamp 1676037725
transform 1 0 392564 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4257
timestamp 1676037725
transform 1 0 392748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4269
timestamp 1676037725
transform 1 0 393852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4281
timestamp 1676037725
transform 1 0 394956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4293
timestamp 1676037725
transform 1 0 396060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4305
timestamp 1676037725
transform 1 0 397164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4311
timestamp 1676037725
transform 1 0 397716 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4313
timestamp 1676037725
transform 1 0 397900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4325
timestamp 1676037725
transform 1 0 399004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4337
timestamp 1676037725
transform 1 0 400108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4349
timestamp 1676037725
transform 1 0 401212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4361
timestamp 1676037725
transform 1 0 402316 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4367
timestamp 1676037725
transform 1 0 402868 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4369
timestamp 1676037725
transform 1 0 403052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4381
timestamp 1676037725
transform 1 0 404156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4393
timestamp 1676037725
transform 1 0 405260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4405
timestamp 1676037725
transform 1 0 406364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4417
timestamp 1676037725
transform 1 0 407468 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4423
timestamp 1676037725
transform 1 0 408020 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4425
timestamp 1676037725
transform 1 0 408204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4437
timestamp 1676037725
transform 1 0 409308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4449
timestamp 1676037725
transform 1 0 410412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4461
timestamp 1676037725
transform 1 0 411516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4473
timestamp 1676037725
transform 1 0 412620 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4479
timestamp 1676037725
transform 1 0 413172 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4481
timestamp 1676037725
transform 1 0 413356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4493
timestamp 1676037725
transform 1 0 414460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4505
timestamp 1676037725
transform 1 0 415564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4517
timestamp 1676037725
transform 1 0 416668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4529
timestamp 1676037725
transform 1 0 417772 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4535
timestamp 1676037725
transform 1 0 418324 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4537
timestamp 1676037725
transform 1 0 418508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4549
timestamp 1676037725
transform 1 0 419612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4561
timestamp 1676037725
transform 1 0 420716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4573
timestamp 1676037725
transform 1 0 421820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4585
timestamp 1676037725
transform 1 0 422924 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4591
timestamp 1676037725
transform 1 0 423476 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4593
timestamp 1676037725
transform 1 0 423660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4605
timestamp 1676037725
transform 1 0 424764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4617
timestamp 1676037725
transform 1 0 425868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4629
timestamp 1676037725
transform 1 0 426972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4641
timestamp 1676037725
transform 1 0 428076 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4647
timestamp 1676037725
transform 1 0 428628 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4649
timestamp 1676037725
transform 1 0 428812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4661
timestamp 1676037725
transform 1 0 429916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4673
timestamp 1676037725
transform 1 0 431020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4685
timestamp 1676037725
transform 1 0 432124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4697
timestamp 1676037725
transform 1 0 433228 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4703
timestamp 1676037725
transform 1 0 433780 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4705
timestamp 1676037725
transform 1 0 433964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4717
timestamp 1676037725
transform 1 0 435068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4729
timestamp 1676037725
transform 1 0 436172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4741
timestamp 1676037725
transform 1 0 437276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4753
timestamp 1676037725
transform 1 0 438380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4759
timestamp 1676037725
transform 1 0 438932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4761
timestamp 1676037725
transform 1 0 439116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4773
timestamp 1676037725
transform 1 0 440220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4785
timestamp 1676037725
transform 1 0 441324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4797
timestamp 1676037725
transform 1 0 442428 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4809
timestamp 1676037725
transform 1 0 443532 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4815
timestamp 1676037725
transform 1 0 444084 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4817
timestamp 1676037725
transform 1 0 444268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4829
timestamp 1676037725
transform 1 0 445372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4841
timestamp 1676037725
transform 1 0 446476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4853
timestamp 1676037725
transform 1 0 447580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4865
timestamp 1676037725
transform 1 0 448684 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4871
timestamp 1676037725
transform 1 0 449236 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4873
timestamp 1676037725
transform 1 0 449420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4885
timestamp 1676037725
transform 1 0 450524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4897
timestamp 1676037725
transform 1 0 451628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4909
timestamp 1676037725
transform 1 0 452732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4921
timestamp 1676037725
transform 1 0 453836 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4927
timestamp 1676037725
transform 1 0 454388 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4929
timestamp 1676037725
transform 1 0 454572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4941
timestamp 1676037725
transform 1 0 455676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4953
timestamp 1676037725
transform 1 0 456780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4965
timestamp 1676037725
transform 1 0 457884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4977
timestamp 1676037725
transform 1 0 458988 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4983
timestamp 1676037725
transform 1 0 459540 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4985
timestamp 1676037725
transform 1 0 459724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4997
timestamp 1676037725
transform 1 0 460828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5009
timestamp 1676037725
transform 1 0 461932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5021
timestamp 1676037725
transform 1 0 463036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5033
timestamp 1676037725
transform 1 0 464140 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5039
timestamp 1676037725
transform 1 0 464692 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5041
timestamp 1676037725
transform 1 0 464876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5053
timestamp 1676037725
transform 1 0 465980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5065
timestamp 1676037725
transform 1 0 467084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5077
timestamp 1676037725
transform 1 0 468188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5089
timestamp 1676037725
transform 1 0 469292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5095
timestamp 1676037725
transform 1 0 469844 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5097
timestamp 1676037725
transform 1 0 470028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5109
timestamp 1676037725
transform 1 0 471132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5121
timestamp 1676037725
transform 1 0 472236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5133
timestamp 1676037725
transform 1 0 473340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5145
timestamp 1676037725
transform 1 0 474444 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5151
timestamp 1676037725
transform 1 0 474996 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5153
timestamp 1676037725
transform 1 0 475180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5165
timestamp 1676037725
transform 1 0 476284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5177
timestamp 1676037725
transform 1 0 477388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5189
timestamp 1676037725
transform 1 0 478492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5201
timestamp 1676037725
transform 1 0 479596 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5207
timestamp 1676037725
transform 1 0 480148 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5209
timestamp 1676037725
transform 1 0 480332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5221
timestamp 1676037725
transform 1 0 481436 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5233
timestamp 1676037725
transform 1 0 482540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5245
timestamp 1676037725
transform 1 0 483644 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5257
timestamp 1676037725
transform 1 0 484748 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5263
timestamp 1676037725
transform 1 0 485300 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5265
timestamp 1676037725
transform 1 0 485484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5277
timestamp 1676037725
transform 1 0 486588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5289
timestamp 1676037725
transform 1 0 487692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5301
timestamp 1676037725
transform 1 0 488796 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5313
timestamp 1676037725
transform 1 0 489900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5319
timestamp 1676037725
transform 1 0 490452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5321
timestamp 1676037725
transform 1 0 490636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5333
timestamp 1676037725
transform 1 0 491740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5345
timestamp 1676037725
transform 1 0 492844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5357
timestamp 1676037725
transform 1 0 493948 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5369
timestamp 1676037725
transform 1 0 495052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5375
timestamp 1676037725
transform 1 0 495604 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5377
timestamp 1676037725
transform 1 0 495788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5389
timestamp 1676037725
transform 1 0 496892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5401
timestamp 1676037725
transform 1 0 497996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5413
timestamp 1676037725
transform 1 0 499100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5425
timestamp 1676037725
transform 1 0 500204 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5431
timestamp 1676037725
transform 1 0 500756 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5433
timestamp 1676037725
transform 1 0 500940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5445
timestamp 1676037725
transform 1 0 502044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5457
timestamp 1676037725
transform 1 0 503148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5469
timestamp 1676037725
transform 1 0 504252 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5481
timestamp 1676037725
transform 1 0 505356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5487
timestamp 1676037725
transform 1 0 505908 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5489
timestamp 1676037725
transform 1 0 506092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5501
timestamp 1676037725
transform 1 0 507196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5513
timestamp 1676037725
transform 1 0 508300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5525
timestamp 1676037725
transform 1 0 509404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5537
timestamp 1676037725
transform 1 0 510508 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5543
timestamp 1676037725
transform 1 0 511060 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5545
timestamp 1676037725
transform 1 0 511244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5557
timestamp 1676037725
transform 1 0 512348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5569
timestamp 1676037725
transform 1 0 513452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5581
timestamp 1676037725
transform 1 0 514556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5593
timestamp 1676037725
transform 1 0 515660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5599
timestamp 1676037725
transform 1 0 516212 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5601
timestamp 1676037725
transform 1 0 516396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5613
timestamp 1676037725
transform 1 0 517500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5625
timestamp 1676037725
transform 1 0 518604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5637
timestamp 1676037725
transform 1 0 519708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5649
timestamp 1676037725
transform 1 0 520812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5655
timestamp 1676037725
transform 1 0 521364 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5657
timestamp 1676037725
transform 1 0 521548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5669
timestamp 1676037725
transform 1 0 522652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5681
timestamp 1676037725
transform 1 0 523756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5693
timestamp 1676037725
transform 1 0 524860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5705
timestamp 1676037725
transform 1 0 525964 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5711
timestamp 1676037725
transform 1 0 526516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5713
timestamp 1676037725
transform 1 0 526700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5725
timestamp 1676037725
transform 1 0 527804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5737
timestamp 1676037725
transform 1 0 528908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5749
timestamp 1676037725
transform 1 0 530012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5761
timestamp 1676037725
transform 1 0 531116 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5767
timestamp 1676037725
transform 1 0 531668 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5769
timestamp 1676037725
transform 1 0 531852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5781
timestamp 1676037725
transform 1 0 532956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5793
timestamp 1676037725
transform 1 0 534060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5805
timestamp 1676037725
transform 1 0 535164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5817
timestamp 1676037725
transform 1 0 536268 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5823
timestamp 1676037725
transform 1 0 536820 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5825
timestamp 1676037725
transform 1 0 537004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5837
timestamp 1676037725
transform 1 0 538108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5849
timestamp 1676037725
transform 1 0 539212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5861
timestamp 1676037725
transform 1 0 540316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5873
timestamp 1676037725
transform 1 0 541420 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5879
timestamp 1676037725
transform 1 0 541972 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5881
timestamp 1676037725
transform 1 0 542156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5893
timestamp 1676037725
transform 1 0 543260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5905
timestamp 1676037725
transform 1 0 544364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5917
timestamp 1676037725
transform 1 0 545468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5929
timestamp 1676037725
transform 1 0 546572 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5935
timestamp 1676037725
transform 1 0 547124 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5937
timestamp 1676037725
transform 1 0 547308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5949
timestamp 1676037725
transform 1 0 548412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5961
timestamp 1676037725
transform 1 0 549516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5973
timestamp 1676037725
transform 1 0 550620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5985
timestamp 1676037725
transform 1 0 551724 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5991
timestamp 1676037725
transform 1 0 552276 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5993
timestamp 1676037725
transform 1 0 552460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6005
timestamp 1676037725
transform 1 0 553564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6017
timestamp 1676037725
transform 1 0 554668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6029
timestamp 1676037725
transform 1 0 555772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6041
timestamp 1676037725
transform 1 0 556876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6047
timestamp 1676037725
transform 1 0 557428 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6049
timestamp 1676037725
transform 1 0 557612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6061
timestamp 1676037725
transform 1 0 558716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6073
timestamp 1676037725
transform 1 0 559820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6085
timestamp 1676037725
transform 1 0 560924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6097
timestamp 1676037725
transform 1 0 562028 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6103
timestamp 1676037725
transform 1 0 562580 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6105
timestamp 1676037725
transform 1 0 562764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6117
timestamp 1676037725
transform 1 0 563868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6129
timestamp 1676037725
transform 1 0 564972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6141
timestamp 1676037725
transform 1 0 566076 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6153
timestamp 1676037725
transform 1 0 567180 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6159
timestamp 1676037725
transform 1 0 567732 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6161
timestamp 1676037725
transform 1 0 567916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6173
timestamp 1676037725
transform 1 0 569020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6185
timestamp 1676037725
transform 1 0 570124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6197
timestamp 1676037725
transform 1 0 571228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6209
timestamp 1676037725
transform 1 0 572332 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6215
timestamp 1676037725
transform 1 0 572884 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6217
timestamp 1676037725
transform 1 0 573068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6229
timestamp 1676037725
transform 1 0 574172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6241
timestamp 1676037725
transform 1 0 575276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6253
timestamp 1676037725
transform 1 0 576380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6265
timestamp 1676037725
transform 1 0 577484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6271
timestamp 1676037725
transform 1 0 578036 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6273
timestamp 1676037725
transform 1 0 578220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6285
timestamp 1676037725
transform 1 0 579324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6297
timestamp 1676037725
transform 1 0 580428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6309
timestamp 1676037725
transform 1 0 581532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6321
timestamp 1676037725
transform 1 0 582636 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6327
timestamp 1676037725
transform 1 0 583188 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6329
timestamp 1676037725
transform 1 0 583372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6341
timestamp 1676037725
transform 1 0 584476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6353
timestamp 1676037725
transform 1 0 585580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6365
timestamp 1676037725
transform 1 0 586684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6377
timestamp 1676037725
transform 1 0 587788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6383
timestamp 1676037725
transform 1 0 588340 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6385
timestamp 1676037725
transform 1 0 588524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6397
timestamp 1676037725
transform 1 0 589628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6409
timestamp 1676037725
transform 1 0 590732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6421
timestamp 1676037725
transform 1 0 591836 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6433
timestamp 1676037725
transform 1 0 592940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6439
timestamp 1676037725
transform 1 0 593492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6441
timestamp 1676037725
transform 1 0 593676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6453
timestamp 1676037725
transform 1 0 594780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6465
timestamp 1676037725
transform 1 0 595884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6477
timestamp 1676037725
transform 1 0 596988 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6489
timestamp 1676037725
transform 1 0 598092 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6495
timestamp 1676037725
transform 1 0 598644 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6497
timestamp 1676037725
transform 1 0 598828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6509
timestamp 1676037725
transform 1 0 599932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6521
timestamp 1676037725
transform 1 0 601036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6533
timestamp 1676037725
transform 1 0 602140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6545
timestamp 1676037725
transform 1 0 603244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6551
timestamp 1676037725
transform 1 0 603796 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6553
timestamp 1676037725
transform 1 0 603980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6565
timestamp 1676037725
transform 1 0 605084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6577
timestamp 1676037725
transform 1 0 606188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6589
timestamp 1676037725
transform 1 0 607292 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6601
timestamp 1676037725
transform 1 0 608396 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6607
timestamp 1676037725
transform 1 0 608948 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6609
timestamp 1676037725
transform 1 0 609132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6621
timestamp 1676037725
transform 1 0 610236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6633
timestamp 1676037725
transform 1 0 611340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6645
timestamp 1676037725
transform 1 0 612444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6657
timestamp 1676037725
transform 1 0 613548 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6663
timestamp 1676037725
transform 1 0 614100 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6665
timestamp 1676037725
transform 1 0 614284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6677
timestamp 1676037725
transform 1 0 615388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6689
timestamp 1676037725
transform 1 0 616492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6701
timestamp 1676037725
transform 1 0 617596 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6713
timestamp 1676037725
transform 1 0 618700 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6719
timestamp 1676037725
transform 1 0 619252 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6721
timestamp 1676037725
transform 1 0 619436 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6733
timestamp 1676037725
transform 1 0 620540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6745
timestamp 1676037725
transform 1 0 621644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6757
timestamp 1676037725
transform 1 0 622748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6769
timestamp 1676037725
transform 1 0 623852 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6775
timestamp 1676037725
transform 1 0 624404 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6777
timestamp 1676037725
transform 1 0 624588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6789
timestamp 1676037725
transform 1 0 625692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6801
timestamp 1676037725
transform 1 0 626796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6813
timestamp 1676037725
transform 1 0 627900 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6825
timestamp 1676037725
transform 1 0 629004 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6831
timestamp 1676037725
transform 1 0 629556 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6833
timestamp 1676037725
transform 1 0 629740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6845
timestamp 1676037725
transform 1 0 630844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6857
timestamp 1676037725
transform 1 0 631948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6869
timestamp 1676037725
transform 1 0 633052 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6881
timestamp 1676037725
transform 1 0 634156 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6887
timestamp 1676037725
transform 1 0 634708 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6889
timestamp 1676037725
transform 1 0 634892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6901
timestamp 1676037725
transform 1 0 635996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6913
timestamp 1676037725
transform 1 0 637100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6925
timestamp 1676037725
transform 1 0 638204 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6937
timestamp 1676037725
transform 1 0 639308 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6943
timestamp 1676037725
transform 1 0 639860 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6945
timestamp 1676037725
transform 1 0 640044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6957
timestamp 1676037725
transform 1 0 641148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6969
timestamp 1676037725
transform 1 0 642252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_6981
timestamp 1676037725
transform 1 0 643356 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_6993
timestamp 1676037725
transform 1 0 644460 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6999
timestamp 1676037725
transform 1 0 645012 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7001
timestamp 1676037725
transform 1 0 645196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7013
timestamp 1676037725
transform 1 0 646300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7025
timestamp 1676037725
transform 1 0 647404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7037
timestamp 1676037725
transform 1 0 648508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_7049
timestamp 1676037725
transform 1 0 649612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7055
timestamp 1676037725
transform 1 0 650164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7057
timestamp 1676037725
transform 1 0 650348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7069
timestamp 1676037725
transform 1 0 651452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7081
timestamp 1676037725
transform 1 0 652556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7093
timestamp 1676037725
transform 1 0 653660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_7105
timestamp 1676037725
transform 1 0 654764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7111
timestamp 1676037725
transform 1 0 655316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7113
timestamp 1676037725
transform 1 0 655500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7125
timestamp 1676037725
transform 1 0 656604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7137
timestamp 1676037725
transform 1 0 657708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7149
timestamp 1676037725
transform 1 0 658812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_7161
timestamp 1676037725
transform 1 0 659916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7167
timestamp 1676037725
transform 1 0 660468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7169
timestamp 1676037725
transform 1 0 660652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7181
timestamp 1676037725
transform 1 0 661756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7193
timestamp 1676037725
transform 1 0 662860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7205
timestamp 1676037725
transform 1 0 663964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_7217
timestamp 1676037725
transform 1 0 665068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7223
timestamp 1676037725
transform 1 0 665620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7225
timestamp 1676037725
transform 1 0 665804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7237
timestamp 1676037725
transform 1 0 666908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7249
timestamp 1676037725
transform 1 0 668012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7261
timestamp 1676037725
transform 1 0 669116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_7273
timestamp 1676037725
transform 1 0 670220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7279
timestamp 1676037725
transform 1 0 670772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7281
timestamp 1676037725
transform 1 0 670956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7293
timestamp 1676037725
transform 1 0 672060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7305
timestamp 1676037725
transform 1 0 673164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7317
timestamp 1676037725
transform 1 0 674268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_7329
timestamp 1676037725
transform 1 0 675372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7335
timestamp 1676037725
transform 1 0 675924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7337
timestamp 1676037725
transform 1 0 676108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7349
timestamp 1676037725
transform 1 0 677212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7361
timestamp 1676037725
transform 1 0 678316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7373
timestamp 1676037725
transform 1 0 679420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_7385
timestamp 1676037725
transform 1 0 680524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7391
timestamp 1676037725
transform 1 0 681076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_7393
timestamp 1676037725
transform 1 0 681260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7405
timestamp 1676037725
transform 1 0 682364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1676037725
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1676037725
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1676037725
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1676037725
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1676037725
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1676037725
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1676037725
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1676037725
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1676037725
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1676037725
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1676037725
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1676037725
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1676037725
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1676037725
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1676037725
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1676037725
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1676037725
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1676037725
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1676037725
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1676037725
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1676037725
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1676037725
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1676037725
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1676037725
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1676037725
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1676037725
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1676037725
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1676037725
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1676037725
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1676037725
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1676037725
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1676037725
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1676037725
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1676037725
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1676037725
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1676037725
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1676037725
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1676037725
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1676037725
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1676037725
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1676037725
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1676037725
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1676037725
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1676037725
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1676037725
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1676037725
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1676037725
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1676037725
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1676037725
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1676037725
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1676037725
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1676037725
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1676037725
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1676037725
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1676037725
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1676037725
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1676037725
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1676037725
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1676037725
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1676037725
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1676037725
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1676037725
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1676037725
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1676037725
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1676037725
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1676037725
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1676037725
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1676037725
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1676037725
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1217
timestamp 1676037725
transform 1 0 113068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1229
timestamp 1676037725
transform 1 0 114172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1241
timestamp 1676037725
transform 1 0 115276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1253
timestamp 1676037725
transform 1 0 116380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1676037725
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1261
timestamp 1676037725
transform 1 0 117116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1273
timestamp 1676037725
transform 1 0 118220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1285
timestamp 1676037725
transform 1 0 119324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1297
timestamp 1676037725
transform 1 0 120428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1309
timestamp 1676037725
transform 1 0 121532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1315
timestamp 1676037725
transform 1 0 122084 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1317
timestamp 1676037725
transform 1 0 122268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1329
timestamp 1676037725
transform 1 0 123372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1341
timestamp 1676037725
transform 1 0 124476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1353
timestamp 1676037725
transform 1 0 125580 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1365
timestamp 1676037725
transform 1 0 126684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1371
timestamp 1676037725
transform 1 0 127236 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1373
timestamp 1676037725
transform 1 0 127420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1385
timestamp 1676037725
transform 1 0 128524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1397
timestamp 1676037725
transform 1 0 129628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1409
timestamp 1676037725
transform 1 0 130732 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1421
timestamp 1676037725
transform 1 0 131836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1427
timestamp 1676037725
transform 1 0 132388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1429
timestamp 1676037725
transform 1 0 132572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1441
timestamp 1676037725
transform 1 0 133676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1453
timestamp 1676037725
transform 1 0 134780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1465
timestamp 1676037725
transform 1 0 135884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1477
timestamp 1676037725
transform 1 0 136988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1483
timestamp 1676037725
transform 1 0 137540 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1485
timestamp 1676037725
transform 1 0 137724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1497
timestamp 1676037725
transform 1 0 138828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1509
timestamp 1676037725
transform 1 0 139932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1521
timestamp 1676037725
transform 1 0 141036 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1533
timestamp 1676037725
transform 1 0 142140 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1539
timestamp 1676037725
transform 1 0 142692 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1541
timestamp 1676037725
transform 1 0 142876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1553
timestamp 1676037725
transform 1 0 143980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1565
timestamp 1676037725
transform 1 0 145084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1577
timestamp 1676037725
transform 1 0 146188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1589
timestamp 1676037725
transform 1 0 147292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1595
timestamp 1676037725
transform 1 0 147844 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1597
timestamp 1676037725
transform 1 0 148028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1609
timestamp 1676037725
transform 1 0 149132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1621
timestamp 1676037725
transform 1 0 150236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1633
timestamp 1676037725
transform 1 0 151340 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1645
timestamp 1676037725
transform 1 0 152444 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1651
timestamp 1676037725
transform 1 0 152996 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1653
timestamp 1676037725
transform 1 0 153180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1665
timestamp 1676037725
transform 1 0 154284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1677
timestamp 1676037725
transform 1 0 155388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1689
timestamp 1676037725
transform 1 0 156492 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1701
timestamp 1676037725
transform 1 0 157596 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1707
timestamp 1676037725
transform 1 0 158148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1709
timestamp 1676037725
transform 1 0 158332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1721
timestamp 1676037725
transform 1 0 159436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1733
timestamp 1676037725
transform 1 0 160540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1745
timestamp 1676037725
transform 1 0 161644 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1757
timestamp 1676037725
transform 1 0 162748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1763
timestamp 1676037725
transform 1 0 163300 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1765
timestamp 1676037725
transform 1 0 163484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1777
timestamp 1676037725
transform 1 0 164588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1789
timestamp 1676037725
transform 1 0 165692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1801
timestamp 1676037725
transform 1 0 166796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1813
timestamp 1676037725
transform 1 0 167900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1819
timestamp 1676037725
transform 1 0 168452 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1821
timestamp 1676037725
transform 1 0 168636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1833
timestamp 1676037725
transform 1 0 169740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1845
timestamp 1676037725
transform 1 0 170844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1857
timestamp 1676037725
transform 1 0 171948 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1869
timestamp 1676037725
transform 1 0 173052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1875
timestamp 1676037725
transform 1 0 173604 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1877
timestamp 1676037725
transform 1 0 173788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1889
timestamp 1676037725
transform 1 0 174892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1901
timestamp 1676037725
transform 1 0 175996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1913
timestamp 1676037725
transform 1 0 177100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1925
timestamp 1676037725
transform 1 0 178204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1931
timestamp 1676037725
transform 1 0 178756 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1933
timestamp 1676037725
transform 1 0 178940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1945
timestamp 1676037725
transform 1 0 180044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1957
timestamp 1676037725
transform 1 0 181148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1969
timestamp 1676037725
transform 1 0 182252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1981
timestamp 1676037725
transform 1 0 183356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1987
timestamp 1676037725
transform 1 0 183908 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1989
timestamp 1676037725
transform 1 0 184092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2001
timestamp 1676037725
transform 1 0 185196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2013
timestamp 1676037725
transform 1 0 186300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2025
timestamp 1676037725
transform 1 0 187404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2037
timestamp 1676037725
transform 1 0 188508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2043
timestamp 1676037725
transform 1 0 189060 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2045
timestamp 1676037725
transform 1 0 189244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2057
timestamp 1676037725
transform 1 0 190348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2069
timestamp 1676037725
transform 1 0 191452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2081
timestamp 1676037725
transform 1 0 192556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2093
timestamp 1676037725
transform 1 0 193660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2099
timestamp 1676037725
transform 1 0 194212 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2101
timestamp 1676037725
transform 1 0 194396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2113
timestamp 1676037725
transform 1 0 195500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2125
timestamp 1676037725
transform 1 0 196604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2137
timestamp 1676037725
transform 1 0 197708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2149
timestamp 1676037725
transform 1 0 198812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2155
timestamp 1676037725
transform 1 0 199364 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2157
timestamp 1676037725
transform 1 0 199548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2169
timestamp 1676037725
transform 1 0 200652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2181
timestamp 1676037725
transform 1 0 201756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2193
timestamp 1676037725
transform 1 0 202860 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2205
timestamp 1676037725
transform 1 0 203964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2211
timestamp 1676037725
transform 1 0 204516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2213
timestamp 1676037725
transform 1 0 204700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2225
timestamp 1676037725
transform 1 0 205804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2237
timestamp 1676037725
transform 1 0 206908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2249
timestamp 1676037725
transform 1 0 208012 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2261
timestamp 1676037725
transform 1 0 209116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2267
timestamp 1676037725
transform 1 0 209668 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2269
timestamp 1676037725
transform 1 0 209852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2281
timestamp 1676037725
transform 1 0 210956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2293
timestamp 1676037725
transform 1 0 212060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2305
timestamp 1676037725
transform 1 0 213164 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2317
timestamp 1676037725
transform 1 0 214268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2323
timestamp 1676037725
transform 1 0 214820 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2325
timestamp 1676037725
transform 1 0 215004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2337
timestamp 1676037725
transform 1 0 216108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2349
timestamp 1676037725
transform 1 0 217212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2361
timestamp 1676037725
transform 1 0 218316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2373
timestamp 1676037725
transform 1 0 219420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2379
timestamp 1676037725
transform 1 0 219972 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2381
timestamp 1676037725
transform 1 0 220156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2393
timestamp 1676037725
transform 1 0 221260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2405
timestamp 1676037725
transform 1 0 222364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2417
timestamp 1676037725
transform 1 0 223468 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2429
timestamp 1676037725
transform 1 0 224572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2435
timestamp 1676037725
transform 1 0 225124 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2437
timestamp 1676037725
transform 1 0 225308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2449
timestamp 1676037725
transform 1 0 226412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2461
timestamp 1676037725
transform 1 0 227516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2473
timestamp 1676037725
transform 1 0 228620 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2485
timestamp 1676037725
transform 1 0 229724 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2491
timestamp 1676037725
transform 1 0 230276 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2493
timestamp 1676037725
transform 1 0 230460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2505
timestamp 1676037725
transform 1 0 231564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2517
timestamp 1676037725
transform 1 0 232668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2529
timestamp 1676037725
transform 1 0 233772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2541
timestamp 1676037725
transform 1 0 234876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2547
timestamp 1676037725
transform 1 0 235428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2549
timestamp 1676037725
transform 1 0 235612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2561
timestamp 1676037725
transform 1 0 236716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2573
timestamp 1676037725
transform 1 0 237820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2585
timestamp 1676037725
transform 1 0 238924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2597
timestamp 1676037725
transform 1 0 240028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2603
timestamp 1676037725
transform 1 0 240580 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2605
timestamp 1676037725
transform 1 0 240764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2617
timestamp 1676037725
transform 1 0 241868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2629
timestamp 1676037725
transform 1 0 242972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2641
timestamp 1676037725
transform 1 0 244076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2653
timestamp 1676037725
transform 1 0 245180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2659
timestamp 1676037725
transform 1 0 245732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2661
timestamp 1676037725
transform 1 0 245916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2673
timestamp 1676037725
transform 1 0 247020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2685
timestamp 1676037725
transform 1 0 248124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2697
timestamp 1676037725
transform 1 0 249228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2709
timestamp 1676037725
transform 1 0 250332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2715
timestamp 1676037725
transform 1 0 250884 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2717
timestamp 1676037725
transform 1 0 251068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2729
timestamp 1676037725
transform 1 0 252172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2741
timestamp 1676037725
transform 1 0 253276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2753
timestamp 1676037725
transform 1 0 254380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2765
timestamp 1676037725
transform 1 0 255484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2771
timestamp 1676037725
transform 1 0 256036 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2773
timestamp 1676037725
transform 1 0 256220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2785
timestamp 1676037725
transform 1 0 257324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2797
timestamp 1676037725
transform 1 0 258428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2809
timestamp 1676037725
transform 1 0 259532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2821
timestamp 1676037725
transform 1 0 260636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2827
timestamp 1676037725
transform 1 0 261188 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2829
timestamp 1676037725
transform 1 0 261372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2841
timestamp 1676037725
transform 1 0 262476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2853
timestamp 1676037725
transform 1 0 263580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2865
timestamp 1676037725
transform 1 0 264684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2877
timestamp 1676037725
transform 1 0 265788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2883
timestamp 1676037725
transform 1 0 266340 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2885
timestamp 1676037725
transform 1 0 266524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2897
timestamp 1676037725
transform 1 0 267628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2909
timestamp 1676037725
transform 1 0 268732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2921
timestamp 1676037725
transform 1 0 269836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2933
timestamp 1676037725
transform 1 0 270940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2939
timestamp 1676037725
transform 1 0 271492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2941
timestamp 1676037725
transform 1 0 271676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2953
timestamp 1676037725
transform 1 0 272780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2965
timestamp 1676037725
transform 1 0 273884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2977
timestamp 1676037725
transform 1 0 274988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2989
timestamp 1676037725
transform 1 0 276092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2995
timestamp 1676037725
transform 1 0 276644 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2997
timestamp 1676037725
transform 1 0 276828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3009
timestamp 1676037725
transform 1 0 277932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3021
timestamp 1676037725
transform 1 0 279036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3033
timestamp 1676037725
transform 1 0 280140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3045
timestamp 1676037725
transform 1 0 281244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3051
timestamp 1676037725
transform 1 0 281796 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3053
timestamp 1676037725
transform 1 0 281980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3065
timestamp 1676037725
transform 1 0 283084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3077
timestamp 1676037725
transform 1 0 284188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3089
timestamp 1676037725
transform 1 0 285292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3101
timestamp 1676037725
transform 1 0 286396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3107
timestamp 1676037725
transform 1 0 286948 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3109
timestamp 1676037725
transform 1 0 287132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3121
timestamp 1676037725
transform 1 0 288236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3133
timestamp 1676037725
transform 1 0 289340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3145
timestamp 1676037725
transform 1 0 290444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3157
timestamp 1676037725
transform 1 0 291548 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3163
timestamp 1676037725
transform 1 0 292100 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3165
timestamp 1676037725
transform 1 0 292284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3177
timestamp 1676037725
transform 1 0 293388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3189
timestamp 1676037725
transform 1 0 294492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3201
timestamp 1676037725
transform 1 0 295596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3213
timestamp 1676037725
transform 1 0 296700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3219
timestamp 1676037725
transform 1 0 297252 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3221
timestamp 1676037725
transform 1 0 297436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3233
timestamp 1676037725
transform 1 0 298540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3245
timestamp 1676037725
transform 1 0 299644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3257
timestamp 1676037725
transform 1 0 300748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3269
timestamp 1676037725
transform 1 0 301852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3275
timestamp 1676037725
transform 1 0 302404 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3277
timestamp 1676037725
transform 1 0 302588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3289
timestamp 1676037725
transform 1 0 303692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3301
timestamp 1676037725
transform 1 0 304796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3313
timestamp 1676037725
transform 1 0 305900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3325
timestamp 1676037725
transform 1 0 307004 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3331
timestamp 1676037725
transform 1 0 307556 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3333
timestamp 1676037725
transform 1 0 307740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3345
timestamp 1676037725
transform 1 0 308844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3357
timestamp 1676037725
transform 1 0 309948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3369
timestamp 1676037725
transform 1 0 311052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3381
timestamp 1676037725
transform 1 0 312156 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3387
timestamp 1676037725
transform 1 0 312708 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3389
timestamp 1676037725
transform 1 0 312892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3401
timestamp 1676037725
transform 1 0 313996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3413
timestamp 1676037725
transform 1 0 315100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3425
timestamp 1676037725
transform 1 0 316204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3437
timestamp 1676037725
transform 1 0 317308 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3443
timestamp 1676037725
transform 1 0 317860 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3445
timestamp 1676037725
transform 1 0 318044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3457
timestamp 1676037725
transform 1 0 319148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3469
timestamp 1676037725
transform 1 0 320252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3481
timestamp 1676037725
transform 1 0 321356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3493
timestamp 1676037725
transform 1 0 322460 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3499
timestamp 1676037725
transform 1 0 323012 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3501
timestamp 1676037725
transform 1 0 323196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3513
timestamp 1676037725
transform 1 0 324300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3525
timestamp 1676037725
transform 1 0 325404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3537
timestamp 1676037725
transform 1 0 326508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3549
timestamp 1676037725
transform 1 0 327612 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3555
timestamp 1676037725
transform 1 0 328164 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3557
timestamp 1676037725
transform 1 0 328348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3569
timestamp 1676037725
transform 1 0 329452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3581
timestamp 1676037725
transform 1 0 330556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3593
timestamp 1676037725
transform 1 0 331660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3605
timestamp 1676037725
transform 1 0 332764 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3611
timestamp 1676037725
transform 1 0 333316 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3613
timestamp 1676037725
transform 1 0 333500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3625
timestamp 1676037725
transform 1 0 334604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3637
timestamp 1676037725
transform 1 0 335708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3649
timestamp 1676037725
transform 1 0 336812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3661
timestamp 1676037725
transform 1 0 337916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3667
timestamp 1676037725
transform 1 0 338468 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3669
timestamp 1676037725
transform 1 0 338652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3681
timestamp 1676037725
transform 1 0 339756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3693
timestamp 1676037725
transform 1 0 340860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3705
timestamp 1676037725
transform 1 0 341964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3717
timestamp 1676037725
transform 1 0 343068 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3723
timestamp 1676037725
transform 1 0 343620 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3725
timestamp 1676037725
transform 1 0 343804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3737
timestamp 1676037725
transform 1 0 344908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3749
timestamp 1676037725
transform 1 0 346012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3761
timestamp 1676037725
transform 1 0 347116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3773
timestamp 1676037725
transform 1 0 348220 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3779
timestamp 1676037725
transform 1 0 348772 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3781
timestamp 1676037725
transform 1 0 348956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3793
timestamp 1676037725
transform 1 0 350060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3805
timestamp 1676037725
transform 1 0 351164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3817
timestamp 1676037725
transform 1 0 352268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3829
timestamp 1676037725
transform 1 0 353372 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3835
timestamp 1676037725
transform 1 0 353924 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3837
timestamp 1676037725
transform 1 0 354108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3849
timestamp 1676037725
transform 1 0 355212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3861
timestamp 1676037725
transform 1 0 356316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3873
timestamp 1676037725
transform 1 0 357420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3885
timestamp 1676037725
transform 1 0 358524 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3891
timestamp 1676037725
transform 1 0 359076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3893
timestamp 1676037725
transform 1 0 359260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3905
timestamp 1676037725
transform 1 0 360364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3917
timestamp 1676037725
transform 1 0 361468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3929
timestamp 1676037725
transform 1 0 362572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3941
timestamp 1676037725
transform 1 0 363676 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3947
timestamp 1676037725
transform 1 0 364228 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3949
timestamp 1676037725
transform 1 0 364412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3961
timestamp 1676037725
transform 1 0 365516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3973
timestamp 1676037725
transform 1 0 366620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3985
timestamp 1676037725
transform 1 0 367724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3997
timestamp 1676037725
transform 1 0 368828 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4003
timestamp 1676037725
transform 1 0 369380 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4005
timestamp 1676037725
transform 1 0 369564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4017
timestamp 1676037725
transform 1 0 370668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4029
timestamp 1676037725
transform 1 0 371772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4041
timestamp 1676037725
transform 1 0 372876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4053
timestamp 1676037725
transform 1 0 373980 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4059
timestamp 1676037725
transform 1 0 374532 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4061
timestamp 1676037725
transform 1 0 374716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4073
timestamp 1676037725
transform 1 0 375820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4085
timestamp 1676037725
transform 1 0 376924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4097
timestamp 1676037725
transform 1 0 378028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4109
timestamp 1676037725
transform 1 0 379132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4115
timestamp 1676037725
transform 1 0 379684 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4117
timestamp 1676037725
transform 1 0 379868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4129
timestamp 1676037725
transform 1 0 380972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4141
timestamp 1676037725
transform 1 0 382076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4153
timestamp 1676037725
transform 1 0 383180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4165
timestamp 1676037725
transform 1 0 384284 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4171
timestamp 1676037725
transform 1 0 384836 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4173
timestamp 1676037725
transform 1 0 385020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4185
timestamp 1676037725
transform 1 0 386124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4197
timestamp 1676037725
transform 1 0 387228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4209
timestamp 1676037725
transform 1 0 388332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4221
timestamp 1676037725
transform 1 0 389436 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4227
timestamp 1676037725
transform 1 0 389988 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4229
timestamp 1676037725
transform 1 0 390172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4241
timestamp 1676037725
transform 1 0 391276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4253
timestamp 1676037725
transform 1 0 392380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4265
timestamp 1676037725
transform 1 0 393484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4277
timestamp 1676037725
transform 1 0 394588 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4283
timestamp 1676037725
transform 1 0 395140 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4285
timestamp 1676037725
transform 1 0 395324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4297
timestamp 1676037725
transform 1 0 396428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4309
timestamp 1676037725
transform 1 0 397532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4321
timestamp 1676037725
transform 1 0 398636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4333
timestamp 1676037725
transform 1 0 399740 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4339
timestamp 1676037725
transform 1 0 400292 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4341
timestamp 1676037725
transform 1 0 400476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4353
timestamp 1676037725
transform 1 0 401580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4365
timestamp 1676037725
transform 1 0 402684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4377
timestamp 1676037725
transform 1 0 403788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4389
timestamp 1676037725
transform 1 0 404892 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4395
timestamp 1676037725
transform 1 0 405444 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4397
timestamp 1676037725
transform 1 0 405628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4409
timestamp 1676037725
transform 1 0 406732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4421
timestamp 1676037725
transform 1 0 407836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4433
timestamp 1676037725
transform 1 0 408940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4445
timestamp 1676037725
transform 1 0 410044 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4451
timestamp 1676037725
transform 1 0 410596 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4453
timestamp 1676037725
transform 1 0 410780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4465
timestamp 1676037725
transform 1 0 411884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4477
timestamp 1676037725
transform 1 0 412988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4489
timestamp 1676037725
transform 1 0 414092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4501
timestamp 1676037725
transform 1 0 415196 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4507
timestamp 1676037725
transform 1 0 415748 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4509
timestamp 1676037725
transform 1 0 415932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4521
timestamp 1676037725
transform 1 0 417036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4533
timestamp 1676037725
transform 1 0 418140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4545
timestamp 1676037725
transform 1 0 419244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4557
timestamp 1676037725
transform 1 0 420348 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4563
timestamp 1676037725
transform 1 0 420900 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4565
timestamp 1676037725
transform 1 0 421084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4577
timestamp 1676037725
transform 1 0 422188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4589
timestamp 1676037725
transform 1 0 423292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4601
timestamp 1676037725
transform 1 0 424396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4613
timestamp 1676037725
transform 1 0 425500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4619
timestamp 1676037725
transform 1 0 426052 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4621
timestamp 1676037725
transform 1 0 426236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4633
timestamp 1676037725
transform 1 0 427340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4645
timestamp 1676037725
transform 1 0 428444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4657
timestamp 1676037725
transform 1 0 429548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4669
timestamp 1676037725
transform 1 0 430652 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4675
timestamp 1676037725
transform 1 0 431204 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4677
timestamp 1676037725
transform 1 0 431388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4689
timestamp 1676037725
transform 1 0 432492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4701
timestamp 1676037725
transform 1 0 433596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4713
timestamp 1676037725
transform 1 0 434700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4725
timestamp 1676037725
transform 1 0 435804 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4731
timestamp 1676037725
transform 1 0 436356 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4733
timestamp 1676037725
transform 1 0 436540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4745
timestamp 1676037725
transform 1 0 437644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4757
timestamp 1676037725
transform 1 0 438748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4769
timestamp 1676037725
transform 1 0 439852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4781
timestamp 1676037725
transform 1 0 440956 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4787
timestamp 1676037725
transform 1 0 441508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4789
timestamp 1676037725
transform 1 0 441692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4801
timestamp 1676037725
transform 1 0 442796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4813
timestamp 1676037725
transform 1 0 443900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4825
timestamp 1676037725
transform 1 0 445004 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4837
timestamp 1676037725
transform 1 0 446108 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4843
timestamp 1676037725
transform 1 0 446660 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4845
timestamp 1676037725
transform 1 0 446844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4857
timestamp 1676037725
transform 1 0 447948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4869
timestamp 1676037725
transform 1 0 449052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4881
timestamp 1676037725
transform 1 0 450156 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4893
timestamp 1676037725
transform 1 0 451260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4899
timestamp 1676037725
transform 1 0 451812 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4901
timestamp 1676037725
transform 1 0 451996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4913
timestamp 1676037725
transform 1 0 453100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4925
timestamp 1676037725
transform 1 0 454204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4937
timestamp 1676037725
transform 1 0 455308 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4949
timestamp 1676037725
transform 1 0 456412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4955
timestamp 1676037725
transform 1 0 456964 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4957
timestamp 1676037725
transform 1 0 457148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4969
timestamp 1676037725
transform 1 0 458252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4981
timestamp 1676037725
transform 1 0 459356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4993
timestamp 1676037725
transform 1 0 460460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5005
timestamp 1676037725
transform 1 0 461564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5011
timestamp 1676037725
transform 1 0 462116 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5013
timestamp 1676037725
transform 1 0 462300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5025
timestamp 1676037725
transform 1 0 463404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5037
timestamp 1676037725
transform 1 0 464508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5049
timestamp 1676037725
transform 1 0 465612 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5061
timestamp 1676037725
transform 1 0 466716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5067
timestamp 1676037725
transform 1 0 467268 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5069
timestamp 1676037725
transform 1 0 467452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5081
timestamp 1676037725
transform 1 0 468556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5093
timestamp 1676037725
transform 1 0 469660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5105
timestamp 1676037725
transform 1 0 470764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5117
timestamp 1676037725
transform 1 0 471868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5123
timestamp 1676037725
transform 1 0 472420 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5125
timestamp 1676037725
transform 1 0 472604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5137
timestamp 1676037725
transform 1 0 473708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5149
timestamp 1676037725
transform 1 0 474812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5161
timestamp 1676037725
transform 1 0 475916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5173
timestamp 1676037725
transform 1 0 477020 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5179
timestamp 1676037725
transform 1 0 477572 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5181
timestamp 1676037725
transform 1 0 477756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5193
timestamp 1676037725
transform 1 0 478860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5205
timestamp 1676037725
transform 1 0 479964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5217
timestamp 1676037725
transform 1 0 481068 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5229
timestamp 1676037725
transform 1 0 482172 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5235
timestamp 1676037725
transform 1 0 482724 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5237
timestamp 1676037725
transform 1 0 482908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5249
timestamp 1676037725
transform 1 0 484012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5261
timestamp 1676037725
transform 1 0 485116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5273
timestamp 1676037725
transform 1 0 486220 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5285
timestamp 1676037725
transform 1 0 487324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5291
timestamp 1676037725
transform 1 0 487876 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5293
timestamp 1676037725
transform 1 0 488060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5305
timestamp 1676037725
transform 1 0 489164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5317
timestamp 1676037725
transform 1 0 490268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5329
timestamp 1676037725
transform 1 0 491372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5341
timestamp 1676037725
transform 1 0 492476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5347
timestamp 1676037725
transform 1 0 493028 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5349
timestamp 1676037725
transform 1 0 493212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5361
timestamp 1676037725
transform 1 0 494316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5373
timestamp 1676037725
transform 1 0 495420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5385
timestamp 1676037725
transform 1 0 496524 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5397
timestamp 1676037725
transform 1 0 497628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5403
timestamp 1676037725
transform 1 0 498180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5405
timestamp 1676037725
transform 1 0 498364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5417
timestamp 1676037725
transform 1 0 499468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5429
timestamp 1676037725
transform 1 0 500572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5441
timestamp 1676037725
transform 1 0 501676 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5453
timestamp 1676037725
transform 1 0 502780 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5459
timestamp 1676037725
transform 1 0 503332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5461
timestamp 1676037725
transform 1 0 503516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5473
timestamp 1676037725
transform 1 0 504620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5485
timestamp 1676037725
transform 1 0 505724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5497
timestamp 1676037725
transform 1 0 506828 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5509
timestamp 1676037725
transform 1 0 507932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5515
timestamp 1676037725
transform 1 0 508484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5517
timestamp 1676037725
transform 1 0 508668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5529
timestamp 1676037725
transform 1 0 509772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5541
timestamp 1676037725
transform 1 0 510876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5553
timestamp 1676037725
transform 1 0 511980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5565
timestamp 1676037725
transform 1 0 513084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5571
timestamp 1676037725
transform 1 0 513636 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5573
timestamp 1676037725
transform 1 0 513820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5585
timestamp 1676037725
transform 1 0 514924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5597
timestamp 1676037725
transform 1 0 516028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5609
timestamp 1676037725
transform 1 0 517132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5621
timestamp 1676037725
transform 1 0 518236 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5627
timestamp 1676037725
transform 1 0 518788 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5629
timestamp 1676037725
transform 1 0 518972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5641
timestamp 1676037725
transform 1 0 520076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5653
timestamp 1676037725
transform 1 0 521180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5665
timestamp 1676037725
transform 1 0 522284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5677
timestamp 1676037725
transform 1 0 523388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5683
timestamp 1676037725
transform 1 0 523940 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5685
timestamp 1676037725
transform 1 0 524124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5697
timestamp 1676037725
transform 1 0 525228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5709
timestamp 1676037725
transform 1 0 526332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5721
timestamp 1676037725
transform 1 0 527436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5733
timestamp 1676037725
transform 1 0 528540 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5739
timestamp 1676037725
transform 1 0 529092 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5741
timestamp 1676037725
transform 1 0 529276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5753
timestamp 1676037725
transform 1 0 530380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5765
timestamp 1676037725
transform 1 0 531484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5777
timestamp 1676037725
transform 1 0 532588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5789
timestamp 1676037725
transform 1 0 533692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5795
timestamp 1676037725
transform 1 0 534244 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5797
timestamp 1676037725
transform 1 0 534428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5809
timestamp 1676037725
transform 1 0 535532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5821
timestamp 1676037725
transform 1 0 536636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5833
timestamp 1676037725
transform 1 0 537740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5845
timestamp 1676037725
transform 1 0 538844 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5851
timestamp 1676037725
transform 1 0 539396 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5853
timestamp 1676037725
transform 1 0 539580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5865
timestamp 1676037725
transform 1 0 540684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5877
timestamp 1676037725
transform 1 0 541788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5889
timestamp 1676037725
transform 1 0 542892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5901
timestamp 1676037725
transform 1 0 543996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5907
timestamp 1676037725
transform 1 0 544548 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5909
timestamp 1676037725
transform 1 0 544732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5921
timestamp 1676037725
transform 1 0 545836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5933
timestamp 1676037725
transform 1 0 546940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5945
timestamp 1676037725
transform 1 0 548044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5957
timestamp 1676037725
transform 1 0 549148 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5963
timestamp 1676037725
transform 1 0 549700 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5965
timestamp 1676037725
transform 1 0 549884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5977
timestamp 1676037725
transform 1 0 550988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5989
timestamp 1676037725
transform 1 0 552092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6001
timestamp 1676037725
transform 1 0 553196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6013
timestamp 1676037725
transform 1 0 554300 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6019
timestamp 1676037725
transform 1 0 554852 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6021
timestamp 1676037725
transform 1 0 555036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6033
timestamp 1676037725
transform 1 0 556140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6045
timestamp 1676037725
transform 1 0 557244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6057
timestamp 1676037725
transform 1 0 558348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6069
timestamp 1676037725
transform 1 0 559452 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6075
timestamp 1676037725
transform 1 0 560004 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6077
timestamp 1676037725
transform 1 0 560188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6089
timestamp 1676037725
transform 1 0 561292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6101
timestamp 1676037725
transform 1 0 562396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6113
timestamp 1676037725
transform 1 0 563500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6125
timestamp 1676037725
transform 1 0 564604 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6131
timestamp 1676037725
transform 1 0 565156 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6133
timestamp 1676037725
transform 1 0 565340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6145
timestamp 1676037725
transform 1 0 566444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6157
timestamp 1676037725
transform 1 0 567548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6169
timestamp 1676037725
transform 1 0 568652 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6181
timestamp 1676037725
transform 1 0 569756 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6187
timestamp 1676037725
transform 1 0 570308 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6189
timestamp 1676037725
transform 1 0 570492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6201
timestamp 1676037725
transform 1 0 571596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6213
timestamp 1676037725
transform 1 0 572700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6225
timestamp 1676037725
transform 1 0 573804 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6237
timestamp 1676037725
transform 1 0 574908 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6243
timestamp 1676037725
transform 1 0 575460 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6245
timestamp 1676037725
transform 1 0 575644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6257
timestamp 1676037725
transform 1 0 576748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6269
timestamp 1676037725
transform 1 0 577852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6281
timestamp 1676037725
transform 1 0 578956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6293
timestamp 1676037725
transform 1 0 580060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6299
timestamp 1676037725
transform 1 0 580612 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6301
timestamp 1676037725
transform 1 0 580796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6313
timestamp 1676037725
transform 1 0 581900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6325
timestamp 1676037725
transform 1 0 583004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6337
timestamp 1676037725
transform 1 0 584108 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6349
timestamp 1676037725
transform 1 0 585212 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6355
timestamp 1676037725
transform 1 0 585764 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6357
timestamp 1676037725
transform 1 0 585948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6369
timestamp 1676037725
transform 1 0 587052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6381
timestamp 1676037725
transform 1 0 588156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6393
timestamp 1676037725
transform 1 0 589260 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6405
timestamp 1676037725
transform 1 0 590364 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6411
timestamp 1676037725
transform 1 0 590916 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6413
timestamp 1676037725
transform 1 0 591100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6425
timestamp 1676037725
transform 1 0 592204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6437
timestamp 1676037725
transform 1 0 593308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6449
timestamp 1676037725
transform 1 0 594412 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6461
timestamp 1676037725
transform 1 0 595516 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6467
timestamp 1676037725
transform 1 0 596068 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6469
timestamp 1676037725
transform 1 0 596252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6481
timestamp 1676037725
transform 1 0 597356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6493
timestamp 1676037725
transform 1 0 598460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6505
timestamp 1676037725
transform 1 0 599564 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6517
timestamp 1676037725
transform 1 0 600668 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6523
timestamp 1676037725
transform 1 0 601220 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6525
timestamp 1676037725
transform 1 0 601404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6537
timestamp 1676037725
transform 1 0 602508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6549
timestamp 1676037725
transform 1 0 603612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6561
timestamp 1676037725
transform 1 0 604716 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6573
timestamp 1676037725
transform 1 0 605820 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6579
timestamp 1676037725
transform 1 0 606372 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6581
timestamp 1676037725
transform 1 0 606556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6593
timestamp 1676037725
transform 1 0 607660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6605
timestamp 1676037725
transform 1 0 608764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6617
timestamp 1676037725
transform 1 0 609868 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6629
timestamp 1676037725
transform 1 0 610972 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6635
timestamp 1676037725
transform 1 0 611524 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6637
timestamp 1676037725
transform 1 0 611708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6649
timestamp 1676037725
transform 1 0 612812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6661
timestamp 1676037725
transform 1 0 613916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6673
timestamp 1676037725
transform 1 0 615020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6685
timestamp 1676037725
transform 1 0 616124 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6691
timestamp 1676037725
transform 1 0 616676 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6693
timestamp 1676037725
transform 1 0 616860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6705
timestamp 1676037725
transform 1 0 617964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6717
timestamp 1676037725
transform 1 0 619068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6729
timestamp 1676037725
transform 1 0 620172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6741
timestamp 1676037725
transform 1 0 621276 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6747
timestamp 1676037725
transform 1 0 621828 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6749
timestamp 1676037725
transform 1 0 622012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6761
timestamp 1676037725
transform 1 0 623116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6773
timestamp 1676037725
transform 1 0 624220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6785
timestamp 1676037725
transform 1 0 625324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6797
timestamp 1676037725
transform 1 0 626428 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6803
timestamp 1676037725
transform 1 0 626980 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6805
timestamp 1676037725
transform 1 0 627164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6817
timestamp 1676037725
transform 1 0 628268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6829
timestamp 1676037725
transform 1 0 629372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6841
timestamp 1676037725
transform 1 0 630476 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6853
timestamp 1676037725
transform 1 0 631580 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6859
timestamp 1676037725
transform 1 0 632132 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6861
timestamp 1676037725
transform 1 0 632316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6873
timestamp 1676037725
transform 1 0 633420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6885
timestamp 1676037725
transform 1 0 634524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6897
timestamp 1676037725
transform 1 0 635628 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6909
timestamp 1676037725
transform 1 0 636732 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6915
timestamp 1676037725
transform 1 0 637284 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6917
timestamp 1676037725
transform 1 0 637468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6929
timestamp 1676037725
transform 1 0 638572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6941
timestamp 1676037725
transform 1 0 639676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6953
timestamp 1676037725
transform 1 0 640780 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6965
timestamp 1676037725
transform 1 0 641884 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6971
timestamp 1676037725
transform 1 0 642436 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6973
timestamp 1676037725
transform 1 0 642620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6985
timestamp 1676037725
transform 1 0 643724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6997
timestamp 1676037725
transform 1 0 644828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7009
timestamp 1676037725
transform 1 0 645932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7021
timestamp 1676037725
transform 1 0 647036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7027
timestamp 1676037725
transform 1 0 647588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7029
timestamp 1676037725
transform 1 0 647772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7041
timestamp 1676037725
transform 1 0 648876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7053
timestamp 1676037725
transform 1 0 649980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7065
timestamp 1676037725
transform 1 0 651084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7077
timestamp 1676037725
transform 1 0 652188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7083
timestamp 1676037725
transform 1 0 652740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7085
timestamp 1676037725
transform 1 0 652924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7097
timestamp 1676037725
transform 1 0 654028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7109
timestamp 1676037725
transform 1 0 655132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7121
timestamp 1676037725
transform 1 0 656236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7133
timestamp 1676037725
transform 1 0 657340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7139
timestamp 1676037725
transform 1 0 657892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7141
timestamp 1676037725
transform 1 0 658076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7153
timestamp 1676037725
transform 1 0 659180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7165
timestamp 1676037725
transform 1 0 660284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7177
timestamp 1676037725
transform 1 0 661388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7189
timestamp 1676037725
transform 1 0 662492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7195
timestamp 1676037725
transform 1 0 663044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7197
timestamp 1676037725
transform 1 0 663228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7209
timestamp 1676037725
transform 1 0 664332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7221
timestamp 1676037725
transform 1 0 665436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7233
timestamp 1676037725
transform 1 0 666540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7245
timestamp 1676037725
transform 1 0 667644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7251
timestamp 1676037725
transform 1 0 668196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7253
timestamp 1676037725
transform 1 0 668380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7265
timestamp 1676037725
transform 1 0 669484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7277
timestamp 1676037725
transform 1 0 670588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7289
timestamp 1676037725
transform 1 0 671692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7301
timestamp 1676037725
transform 1 0 672796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7307
timestamp 1676037725
transform 1 0 673348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7309
timestamp 1676037725
transform 1 0 673532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7321
timestamp 1676037725
transform 1 0 674636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7333
timestamp 1676037725
transform 1 0 675740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7345
timestamp 1676037725
transform 1 0 676844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7357
timestamp 1676037725
transform 1 0 677948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7363
timestamp 1676037725
transform 1 0 678500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7365
timestamp 1676037725
transform 1 0 678684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7377
timestamp 1676037725
transform 1 0 679788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7389
timestamp 1676037725
transform 1 0 680892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7401
timestamp 1676037725
transform 1 0 681996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1676037725
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1676037725
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1676037725
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1676037725
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1676037725
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1676037725
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1676037725
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1676037725
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1676037725
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1676037725
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1676037725
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1676037725
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1676037725
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1676037725
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1676037725
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1676037725
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1676037725
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1676037725
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1676037725
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1676037725
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1676037725
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1676037725
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1676037725
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1676037725
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1676037725
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1676037725
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1676037725
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1676037725
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1676037725
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1676037725
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1676037725
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1676037725
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1676037725
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1676037725
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1676037725
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1676037725
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1676037725
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1676037725
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1676037725
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1676037725
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1676037725
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1676037725
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1676037725
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1676037725
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1676037725
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1676037725
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1676037725
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1676037725
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1676037725
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1676037725
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1676037725
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1676037725
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1676037725
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1676037725
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1676037725
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1676037725
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1676037725
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1676037725
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1676037725
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1676037725
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1676037725
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1676037725
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1676037725
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1676037725
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1676037725
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1676037725
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1676037725
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1676037725
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1676037725
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1676037725
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1676037725
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1676037725
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1676037725
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1245
timestamp 1676037725
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1257
timestamp 1676037725
transform 1 0 116748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1269
timestamp 1676037725
transform 1 0 117852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1281
timestamp 1676037725
transform 1 0 118956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1287
timestamp 1676037725
transform 1 0 119508 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1289
timestamp 1676037725
transform 1 0 119692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1301
timestamp 1676037725
transform 1 0 120796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1313
timestamp 1676037725
transform 1 0 121900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1325
timestamp 1676037725
transform 1 0 123004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1337
timestamp 1676037725
transform 1 0 124108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1343
timestamp 1676037725
transform 1 0 124660 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1345
timestamp 1676037725
transform 1 0 124844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1357
timestamp 1676037725
transform 1 0 125948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1369
timestamp 1676037725
transform 1 0 127052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1381
timestamp 1676037725
transform 1 0 128156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1393
timestamp 1676037725
transform 1 0 129260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1399
timestamp 1676037725
transform 1 0 129812 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1401
timestamp 1676037725
transform 1 0 129996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1413
timestamp 1676037725
transform 1 0 131100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1425
timestamp 1676037725
transform 1 0 132204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1437
timestamp 1676037725
transform 1 0 133308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1449
timestamp 1676037725
transform 1 0 134412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1455
timestamp 1676037725
transform 1 0 134964 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1457
timestamp 1676037725
transform 1 0 135148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1469
timestamp 1676037725
transform 1 0 136252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1481
timestamp 1676037725
transform 1 0 137356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1493
timestamp 1676037725
transform 1 0 138460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1505
timestamp 1676037725
transform 1 0 139564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1511
timestamp 1676037725
transform 1 0 140116 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1513
timestamp 1676037725
transform 1 0 140300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1525
timestamp 1676037725
transform 1 0 141404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1537
timestamp 1676037725
transform 1 0 142508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1549
timestamp 1676037725
transform 1 0 143612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1561
timestamp 1676037725
transform 1 0 144716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1567
timestamp 1676037725
transform 1 0 145268 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1569
timestamp 1676037725
transform 1 0 145452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1581
timestamp 1676037725
transform 1 0 146556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1593
timestamp 1676037725
transform 1 0 147660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1605
timestamp 1676037725
transform 1 0 148764 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1617
timestamp 1676037725
transform 1 0 149868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1623
timestamp 1676037725
transform 1 0 150420 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1625
timestamp 1676037725
transform 1 0 150604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1637
timestamp 1676037725
transform 1 0 151708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1649
timestamp 1676037725
transform 1 0 152812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1661
timestamp 1676037725
transform 1 0 153916 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1673
timestamp 1676037725
transform 1 0 155020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1679
timestamp 1676037725
transform 1 0 155572 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1681
timestamp 1676037725
transform 1 0 155756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1693
timestamp 1676037725
transform 1 0 156860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1705
timestamp 1676037725
transform 1 0 157964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1717
timestamp 1676037725
transform 1 0 159068 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1729
timestamp 1676037725
transform 1 0 160172 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1735
timestamp 1676037725
transform 1 0 160724 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1737
timestamp 1676037725
transform 1 0 160908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1749
timestamp 1676037725
transform 1 0 162012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1761
timestamp 1676037725
transform 1 0 163116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1773
timestamp 1676037725
transform 1 0 164220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1785
timestamp 1676037725
transform 1 0 165324 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1791
timestamp 1676037725
transform 1 0 165876 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1793
timestamp 1676037725
transform 1 0 166060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1805
timestamp 1676037725
transform 1 0 167164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1817
timestamp 1676037725
transform 1 0 168268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1829
timestamp 1676037725
transform 1 0 169372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1841
timestamp 1676037725
transform 1 0 170476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1847
timestamp 1676037725
transform 1 0 171028 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1849
timestamp 1676037725
transform 1 0 171212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1861
timestamp 1676037725
transform 1 0 172316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1873
timestamp 1676037725
transform 1 0 173420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1885
timestamp 1676037725
transform 1 0 174524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1897
timestamp 1676037725
transform 1 0 175628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1903
timestamp 1676037725
transform 1 0 176180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1905
timestamp 1676037725
transform 1 0 176364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1917
timestamp 1676037725
transform 1 0 177468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1929
timestamp 1676037725
transform 1 0 178572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1941
timestamp 1676037725
transform 1 0 179676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1953
timestamp 1676037725
transform 1 0 180780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1959
timestamp 1676037725
transform 1 0 181332 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1961
timestamp 1676037725
transform 1 0 181516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1973
timestamp 1676037725
transform 1 0 182620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1985
timestamp 1676037725
transform 1 0 183724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1997
timestamp 1676037725
transform 1 0 184828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2009
timestamp 1676037725
transform 1 0 185932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2015
timestamp 1676037725
transform 1 0 186484 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2017
timestamp 1676037725
transform 1 0 186668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2029
timestamp 1676037725
transform 1 0 187772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2041
timestamp 1676037725
transform 1 0 188876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2053
timestamp 1676037725
transform 1 0 189980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2065
timestamp 1676037725
transform 1 0 191084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2071
timestamp 1676037725
transform 1 0 191636 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2073
timestamp 1676037725
transform 1 0 191820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2085
timestamp 1676037725
transform 1 0 192924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2097
timestamp 1676037725
transform 1 0 194028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2109
timestamp 1676037725
transform 1 0 195132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2121
timestamp 1676037725
transform 1 0 196236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2127
timestamp 1676037725
transform 1 0 196788 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2129
timestamp 1676037725
transform 1 0 196972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2141
timestamp 1676037725
transform 1 0 198076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2153
timestamp 1676037725
transform 1 0 199180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2165
timestamp 1676037725
transform 1 0 200284 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2177
timestamp 1676037725
transform 1 0 201388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2183
timestamp 1676037725
transform 1 0 201940 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2185
timestamp 1676037725
transform 1 0 202124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2197
timestamp 1676037725
transform 1 0 203228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2209
timestamp 1676037725
transform 1 0 204332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2221
timestamp 1676037725
transform 1 0 205436 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2233
timestamp 1676037725
transform 1 0 206540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2239
timestamp 1676037725
transform 1 0 207092 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2241
timestamp 1676037725
transform 1 0 207276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2253
timestamp 1676037725
transform 1 0 208380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2265
timestamp 1676037725
transform 1 0 209484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2277
timestamp 1676037725
transform 1 0 210588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2289
timestamp 1676037725
transform 1 0 211692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2295
timestamp 1676037725
transform 1 0 212244 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2297
timestamp 1676037725
transform 1 0 212428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2309
timestamp 1676037725
transform 1 0 213532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2321
timestamp 1676037725
transform 1 0 214636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2333
timestamp 1676037725
transform 1 0 215740 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2345
timestamp 1676037725
transform 1 0 216844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2351
timestamp 1676037725
transform 1 0 217396 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2353
timestamp 1676037725
transform 1 0 217580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2365
timestamp 1676037725
transform 1 0 218684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2377
timestamp 1676037725
transform 1 0 219788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2389
timestamp 1676037725
transform 1 0 220892 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2401
timestamp 1676037725
transform 1 0 221996 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2407
timestamp 1676037725
transform 1 0 222548 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2409
timestamp 1676037725
transform 1 0 222732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2421
timestamp 1676037725
transform 1 0 223836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2433
timestamp 1676037725
transform 1 0 224940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2445
timestamp 1676037725
transform 1 0 226044 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2457
timestamp 1676037725
transform 1 0 227148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2463
timestamp 1676037725
transform 1 0 227700 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2465
timestamp 1676037725
transform 1 0 227884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2477
timestamp 1676037725
transform 1 0 228988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2489
timestamp 1676037725
transform 1 0 230092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2501
timestamp 1676037725
transform 1 0 231196 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2513
timestamp 1676037725
transform 1 0 232300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2519
timestamp 1676037725
transform 1 0 232852 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2521
timestamp 1676037725
transform 1 0 233036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2533
timestamp 1676037725
transform 1 0 234140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2545
timestamp 1676037725
transform 1 0 235244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2557
timestamp 1676037725
transform 1 0 236348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2569
timestamp 1676037725
transform 1 0 237452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2575
timestamp 1676037725
transform 1 0 238004 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2577
timestamp 1676037725
transform 1 0 238188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2589
timestamp 1676037725
transform 1 0 239292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2601
timestamp 1676037725
transform 1 0 240396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2613
timestamp 1676037725
transform 1 0 241500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2625
timestamp 1676037725
transform 1 0 242604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2631
timestamp 1676037725
transform 1 0 243156 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2633
timestamp 1676037725
transform 1 0 243340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2645
timestamp 1676037725
transform 1 0 244444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2657
timestamp 1676037725
transform 1 0 245548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2669
timestamp 1676037725
transform 1 0 246652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2681
timestamp 1676037725
transform 1 0 247756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2687
timestamp 1676037725
transform 1 0 248308 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2689
timestamp 1676037725
transform 1 0 248492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2701
timestamp 1676037725
transform 1 0 249596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2713
timestamp 1676037725
transform 1 0 250700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2725
timestamp 1676037725
transform 1 0 251804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2737
timestamp 1676037725
transform 1 0 252908 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2743
timestamp 1676037725
transform 1 0 253460 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2745
timestamp 1676037725
transform 1 0 253644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2757
timestamp 1676037725
transform 1 0 254748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2769
timestamp 1676037725
transform 1 0 255852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2781
timestamp 1676037725
transform 1 0 256956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2793
timestamp 1676037725
transform 1 0 258060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2799
timestamp 1676037725
transform 1 0 258612 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2801
timestamp 1676037725
transform 1 0 258796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2813
timestamp 1676037725
transform 1 0 259900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2825
timestamp 1676037725
transform 1 0 261004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2837
timestamp 1676037725
transform 1 0 262108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2849
timestamp 1676037725
transform 1 0 263212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2855
timestamp 1676037725
transform 1 0 263764 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2857
timestamp 1676037725
transform 1 0 263948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2869
timestamp 1676037725
transform 1 0 265052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2881
timestamp 1676037725
transform 1 0 266156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2893
timestamp 1676037725
transform 1 0 267260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2905
timestamp 1676037725
transform 1 0 268364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2911
timestamp 1676037725
transform 1 0 268916 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2913
timestamp 1676037725
transform 1 0 269100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2925
timestamp 1676037725
transform 1 0 270204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2937
timestamp 1676037725
transform 1 0 271308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2949
timestamp 1676037725
transform 1 0 272412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2961
timestamp 1676037725
transform 1 0 273516 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2967
timestamp 1676037725
transform 1 0 274068 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2969
timestamp 1676037725
transform 1 0 274252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2981
timestamp 1676037725
transform 1 0 275356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2993
timestamp 1676037725
transform 1 0 276460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3005
timestamp 1676037725
transform 1 0 277564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3017
timestamp 1676037725
transform 1 0 278668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3023
timestamp 1676037725
transform 1 0 279220 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3025
timestamp 1676037725
transform 1 0 279404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3037
timestamp 1676037725
transform 1 0 280508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3049
timestamp 1676037725
transform 1 0 281612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3061
timestamp 1676037725
transform 1 0 282716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3073
timestamp 1676037725
transform 1 0 283820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3079
timestamp 1676037725
transform 1 0 284372 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3081
timestamp 1676037725
transform 1 0 284556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3093
timestamp 1676037725
transform 1 0 285660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3105
timestamp 1676037725
transform 1 0 286764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3117
timestamp 1676037725
transform 1 0 287868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3129
timestamp 1676037725
transform 1 0 288972 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3135
timestamp 1676037725
transform 1 0 289524 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3137
timestamp 1676037725
transform 1 0 289708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3149
timestamp 1676037725
transform 1 0 290812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3161
timestamp 1676037725
transform 1 0 291916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3173
timestamp 1676037725
transform 1 0 293020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3185
timestamp 1676037725
transform 1 0 294124 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3191
timestamp 1676037725
transform 1 0 294676 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3193
timestamp 1676037725
transform 1 0 294860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3205
timestamp 1676037725
transform 1 0 295964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3217
timestamp 1676037725
transform 1 0 297068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3229
timestamp 1676037725
transform 1 0 298172 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3241
timestamp 1676037725
transform 1 0 299276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3247
timestamp 1676037725
transform 1 0 299828 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3249
timestamp 1676037725
transform 1 0 300012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3261
timestamp 1676037725
transform 1 0 301116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3273
timestamp 1676037725
transform 1 0 302220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3285
timestamp 1676037725
transform 1 0 303324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3297
timestamp 1676037725
transform 1 0 304428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3303
timestamp 1676037725
transform 1 0 304980 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3305
timestamp 1676037725
transform 1 0 305164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3317
timestamp 1676037725
transform 1 0 306268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3329
timestamp 1676037725
transform 1 0 307372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3341
timestamp 1676037725
transform 1 0 308476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3353
timestamp 1676037725
transform 1 0 309580 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3359
timestamp 1676037725
transform 1 0 310132 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3361
timestamp 1676037725
transform 1 0 310316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3373
timestamp 1676037725
transform 1 0 311420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3385
timestamp 1676037725
transform 1 0 312524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3397
timestamp 1676037725
transform 1 0 313628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3409
timestamp 1676037725
transform 1 0 314732 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3415
timestamp 1676037725
transform 1 0 315284 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3417
timestamp 1676037725
transform 1 0 315468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3429
timestamp 1676037725
transform 1 0 316572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3441
timestamp 1676037725
transform 1 0 317676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3453
timestamp 1676037725
transform 1 0 318780 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3465
timestamp 1676037725
transform 1 0 319884 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3471
timestamp 1676037725
transform 1 0 320436 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3473
timestamp 1676037725
transform 1 0 320620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3485
timestamp 1676037725
transform 1 0 321724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3497
timestamp 1676037725
transform 1 0 322828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3509
timestamp 1676037725
transform 1 0 323932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3521
timestamp 1676037725
transform 1 0 325036 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3527
timestamp 1676037725
transform 1 0 325588 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3529
timestamp 1676037725
transform 1 0 325772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3541
timestamp 1676037725
transform 1 0 326876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3553
timestamp 1676037725
transform 1 0 327980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3565
timestamp 1676037725
transform 1 0 329084 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3577
timestamp 1676037725
transform 1 0 330188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3583
timestamp 1676037725
transform 1 0 330740 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3585
timestamp 1676037725
transform 1 0 330924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3597
timestamp 1676037725
transform 1 0 332028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3609
timestamp 1676037725
transform 1 0 333132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3621
timestamp 1676037725
transform 1 0 334236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3633
timestamp 1676037725
transform 1 0 335340 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3639
timestamp 1676037725
transform 1 0 335892 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3641
timestamp 1676037725
transform 1 0 336076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3653
timestamp 1676037725
transform 1 0 337180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3665
timestamp 1676037725
transform 1 0 338284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3677
timestamp 1676037725
transform 1 0 339388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3689
timestamp 1676037725
transform 1 0 340492 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3695
timestamp 1676037725
transform 1 0 341044 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3697
timestamp 1676037725
transform 1 0 341228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3709
timestamp 1676037725
transform 1 0 342332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3721
timestamp 1676037725
transform 1 0 343436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3733
timestamp 1676037725
transform 1 0 344540 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3745
timestamp 1676037725
transform 1 0 345644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3751
timestamp 1676037725
transform 1 0 346196 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3753
timestamp 1676037725
transform 1 0 346380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3765
timestamp 1676037725
transform 1 0 347484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3777
timestamp 1676037725
transform 1 0 348588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3789
timestamp 1676037725
transform 1 0 349692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3801
timestamp 1676037725
transform 1 0 350796 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3807
timestamp 1676037725
transform 1 0 351348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3809
timestamp 1676037725
transform 1 0 351532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3821
timestamp 1676037725
transform 1 0 352636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3833
timestamp 1676037725
transform 1 0 353740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3845
timestamp 1676037725
transform 1 0 354844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3857
timestamp 1676037725
transform 1 0 355948 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3863
timestamp 1676037725
transform 1 0 356500 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3865
timestamp 1676037725
transform 1 0 356684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3877
timestamp 1676037725
transform 1 0 357788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3889
timestamp 1676037725
transform 1 0 358892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3901
timestamp 1676037725
transform 1 0 359996 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3913
timestamp 1676037725
transform 1 0 361100 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3919
timestamp 1676037725
transform 1 0 361652 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3921
timestamp 1676037725
transform 1 0 361836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3933
timestamp 1676037725
transform 1 0 362940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3945
timestamp 1676037725
transform 1 0 364044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3957
timestamp 1676037725
transform 1 0 365148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3969
timestamp 1676037725
transform 1 0 366252 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3975
timestamp 1676037725
transform 1 0 366804 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3977
timestamp 1676037725
transform 1 0 366988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3989
timestamp 1676037725
transform 1 0 368092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4001
timestamp 1676037725
transform 1 0 369196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4013
timestamp 1676037725
transform 1 0 370300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4025
timestamp 1676037725
transform 1 0 371404 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4031
timestamp 1676037725
transform 1 0 371956 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4033
timestamp 1676037725
transform 1 0 372140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4045
timestamp 1676037725
transform 1 0 373244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4057
timestamp 1676037725
transform 1 0 374348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4069
timestamp 1676037725
transform 1 0 375452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4081
timestamp 1676037725
transform 1 0 376556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4087
timestamp 1676037725
transform 1 0 377108 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4089
timestamp 1676037725
transform 1 0 377292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4101
timestamp 1676037725
transform 1 0 378396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4113
timestamp 1676037725
transform 1 0 379500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4125
timestamp 1676037725
transform 1 0 380604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4137
timestamp 1676037725
transform 1 0 381708 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4143
timestamp 1676037725
transform 1 0 382260 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4145
timestamp 1676037725
transform 1 0 382444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4157
timestamp 1676037725
transform 1 0 383548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4169
timestamp 1676037725
transform 1 0 384652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4181
timestamp 1676037725
transform 1 0 385756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4193
timestamp 1676037725
transform 1 0 386860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4199
timestamp 1676037725
transform 1 0 387412 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4201
timestamp 1676037725
transform 1 0 387596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4213
timestamp 1676037725
transform 1 0 388700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4225
timestamp 1676037725
transform 1 0 389804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4237
timestamp 1676037725
transform 1 0 390908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4249
timestamp 1676037725
transform 1 0 392012 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4255
timestamp 1676037725
transform 1 0 392564 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4257
timestamp 1676037725
transform 1 0 392748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4269
timestamp 1676037725
transform 1 0 393852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4281
timestamp 1676037725
transform 1 0 394956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4293
timestamp 1676037725
transform 1 0 396060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4305
timestamp 1676037725
transform 1 0 397164 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4311
timestamp 1676037725
transform 1 0 397716 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4313
timestamp 1676037725
transform 1 0 397900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4325
timestamp 1676037725
transform 1 0 399004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4337
timestamp 1676037725
transform 1 0 400108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4349
timestamp 1676037725
transform 1 0 401212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4361
timestamp 1676037725
transform 1 0 402316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4367
timestamp 1676037725
transform 1 0 402868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4369
timestamp 1676037725
transform 1 0 403052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4381
timestamp 1676037725
transform 1 0 404156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4393
timestamp 1676037725
transform 1 0 405260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4405
timestamp 1676037725
transform 1 0 406364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4417
timestamp 1676037725
transform 1 0 407468 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4423
timestamp 1676037725
transform 1 0 408020 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4425
timestamp 1676037725
transform 1 0 408204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4437
timestamp 1676037725
transform 1 0 409308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4449
timestamp 1676037725
transform 1 0 410412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4461
timestamp 1676037725
transform 1 0 411516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4473
timestamp 1676037725
transform 1 0 412620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4479
timestamp 1676037725
transform 1 0 413172 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4481
timestamp 1676037725
transform 1 0 413356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4493
timestamp 1676037725
transform 1 0 414460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4505
timestamp 1676037725
transform 1 0 415564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4517
timestamp 1676037725
transform 1 0 416668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4529
timestamp 1676037725
transform 1 0 417772 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4535
timestamp 1676037725
transform 1 0 418324 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4537
timestamp 1676037725
transform 1 0 418508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4549
timestamp 1676037725
transform 1 0 419612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4561
timestamp 1676037725
transform 1 0 420716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4573
timestamp 1676037725
transform 1 0 421820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4585
timestamp 1676037725
transform 1 0 422924 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4591
timestamp 1676037725
transform 1 0 423476 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4593
timestamp 1676037725
transform 1 0 423660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4605
timestamp 1676037725
transform 1 0 424764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4617
timestamp 1676037725
transform 1 0 425868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4629
timestamp 1676037725
transform 1 0 426972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4641
timestamp 1676037725
transform 1 0 428076 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4647
timestamp 1676037725
transform 1 0 428628 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4649
timestamp 1676037725
transform 1 0 428812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4661
timestamp 1676037725
transform 1 0 429916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4673
timestamp 1676037725
transform 1 0 431020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4685
timestamp 1676037725
transform 1 0 432124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4697
timestamp 1676037725
transform 1 0 433228 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4703
timestamp 1676037725
transform 1 0 433780 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4705
timestamp 1676037725
transform 1 0 433964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4717
timestamp 1676037725
transform 1 0 435068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4729
timestamp 1676037725
transform 1 0 436172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4741
timestamp 1676037725
transform 1 0 437276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4753
timestamp 1676037725
transform 1 0 438380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4759
timestamp 1676037725
transform 1 0 438932 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4761
timestamp 1676037725
transform 1 0 439116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4773
timestamp 1676037725
transform 1 0 440220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4785
timestamp 1676037725
transform 1 0 441324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4797
timestamp 1676037725
transform 1 0 442428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4809
timestamp 1676037725
transform 1 0 443532 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4815
timestamp 1676037725
transform 1 0 444084 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4817
timestamp 1676037725
transform 1 0 444268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4829
timestamp 1676037725
transform 1 0 445372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4841
timestamp 1676037725
transform 1 0 446476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4853
timestamp 1676037725
transform 1 0 447580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4865
timestamp 1676037725
transform 1 0 448684 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4871
timestamp 1676037725
transform 1 0 449236 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4873
timestamp 1676037725
transform 1 0 449420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4885
timestamp 1676037725
transform 1 0 450524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4897
timestamp 1676037725
transform 1 0 451628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4909
timestamp 1676037725
transform 1 0 452732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4921
timestamp 1676037725
transform 1 0 453836 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4927
timestamp 1676037725
transform 1 0 454388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4929
timestamp 1676037725
transform 1 0 454572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4941
timestamp 1676037725
transform 1 0 455676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4953
timestamp 1676037725
transform 1 0 456780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4965
timestamp 1676037725
transform 1 0 457884 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4977
timestamp 1676037725
transform 1 0 458988 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4983
timestamp 1676037725
transform 1 0 459540 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4985
timestamp 1676037725
transform 1 0 459724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4997
timestamp 1676037725
transform 1 0 460828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5009
timestamp 1676037725
transform 1 0 461932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5021
timestamp 1676037725
transform 1 0 463036 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5033
timestamp 1676037725
transform 1 0 464140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5039
timestamp 1676037725
transform 1 0 464692 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5041
timestamp 1676037725
transform 1 0 464876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5053
timestamp 1676037725
transform 1 0 465980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5065
timestamp 1676037725
transform 1 0 467084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5077
timestamp 1676037725
transform 1 0 468188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5089
timestamp 1676037725
transform 1 0 469292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5095
timestamp 1676037725
transform 1 0 469844 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5097
timestamp 1676037725
transform 1 0 470028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5109
timestamp 1676037725
transform 1 0 471132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5121
timestamp 1676037725
transform 1 0 472236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5133
timestamp 1676037725
transform 1 0 473340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5145
timestamp 1676037725
transform 1 0 474444 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5151
timestamp 1676037725
transform 1 0 474996 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5153
timestamp 1676037725
transform 1 0 475180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5165
timestamp 1676037725
transform 1 0 476284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5177
timestamp 1676037725
transform 1 0 477388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5189
timestamp 1676037725
transform 1 0 478492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5201
timestamp 1676037725
transform 1 0 479596 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5207
timestamp 1676037725
transform 1 0 480148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5209
timestamp 1676037725
transform 1 0 480332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5221
timestamp 1676037725
transform 1 0 481436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5233
timestamp 1676037725
transform 1 0 482540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5245
timestamp 1676037725
transform 1 0 483644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5257
timestamp 1676037725
transform 1 0 484748 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5263
timestamp 1676037725
transform 1 0 485300 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5265
timestamp 1676037725
transform 1 0 485484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5277
timestamp 1676037725
transform 1 0 486588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5289
timestamp 1676037725
transform 1 0 487692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5301
timestamp 1676037725
transform 1 0 488796 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5313
timestamp 1676037725
transform 1 0 489900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5319
timestamp 1676037725
transform 1 0 490452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5321
timestamp 1676037725
transform 1 0 490636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5333
timestamp 1676037725
transform 1 0 491740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5345
timestamp 1676037725
transform 1 0 492844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5357
timestamp 1676037725
transform 1 0 493948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5369
timestamp 1676037725
transform 1 0 495052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5375
timestamp 1676037725
transform 1 0 495604 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5377
timestamp 1676037725
transform 1 0 495788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5389
timestamp 1676037725
transform 1 0 496892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5401
timestamp 1676037725
transform 1 0 497996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5413
timestamp 1676037725
transform 1 0 499100 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5425
timestamp 1676037725
transform 1 0 500204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5431
timestamp 1676037725
transform 1 0 500756 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5433
timestamp 1676037725
transform 1 0 500940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5445
timestamp 1676037725
transform 1 0 502044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5457
timestamp 1676037725
transform 1 0 503148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5469
timestamp 1676037725
transform 1 0 504252 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5481
timestamp 1676037725
transform 1 0 505356 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5487
timestamp 1676037725
transform 1 0 505908 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5489
timestamp 1676037725
transform 1 0 506092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5501
timestamp 1676037725
transform 1 0 507196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5513
timestamp 1676037725
transform 1 0 508300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5525
timestamp 1676037725
transform 1 0 509404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5537
timestamp 1676037725
transform 1 0 510508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5543
timestamp 1676037725
transform 1 0 511060 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5545
timestamp 1676037725
transform 1 0 511244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5557
timestamp 1676037725
transform 1 0 512348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5569
timestamp 1676037725
transform 1 0 513452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5581
timestamp 1676037725
transform 1 0 514556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5593
timestamp 1676037725
transform 1 0 515660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5599
timestamp 1676037725
transform 1 0 516212 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5601
timestamp 1676037725
transform 1 0 516396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5613
timestamp 1676037725
transform 1 0 517500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5625
timestamp 1676037725
transform 1 0 518604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5637
timestamp 1676037725
transform 1 0 519708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5649
timestamp 1676037725
transform 1 0 520812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5655
timestamp 1676037725
transform 1 0 521364 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5657
timestamp 1676037725
transform 1 0 521548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5669
timestamp 1676037725
transform 1 0 522652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5681
timestamp 1676037725
transform 1 0 523756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5693
timestamp 1676037725
transform 1 0 524860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5705
timestamp 1676037725
transform 1 0 525964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5711
timestamp 1676037725
transform 1 0 526516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5713
timestamp 1676037725
transform 1 0 526700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5725
timestamp 1676037725
transform 1 0 527804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5737
timestamp 1676037725
transform 1 0 528908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5749
timestamp 1676037725
transform 1 0 530012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5761
timestamp 1676037725
transform 1 0 531116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5767
timestamp 1676037725
transform 1 0 531668 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5769
timestamp 1676037725
transform 1 0 531852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5781
timestamp 1676037725
transform 1 0 532956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5793
timestamp 1676037725
transform 1 0 534060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5805
timestamp 1676037725
transform 1 0 535164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5817
timestamp 1676037725
transform 1 0 536268 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5823
timestamp 1676037725
transform 1 0 536820 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5825
timestamp 1676037725
transform 1 0 537004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5837
timestamp 1676037725
transform 1 0 538108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5849
timestamp 1676037725
transform 1 0 539212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5861
timestamp 1676037725
transform 1 0 540316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5873
timestamp 1676037725
transform 1 0 541420 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5879
timestamp 1676037725
transform 1 0 541972 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5881
timestamp 1676037725
transform 1 0 542156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5893
timestamp 1676037725
transform 1 0 543260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5905
timestamp 1676037725
transform 1 0 544364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5917
timestamp 1676037725
transform 1 0 545468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5929
timestamp 1676037725
transform 1 0 546572 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5935
timestamp 1676037725
transform 1 0 547124 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5937
timestamp 1676037725
transform 1 0 547308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5949
timestamp 1676037725
transform 1 0 548412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5961
timestamp 1676037725
transform 1 0 549516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5973
timestamp 1676037725
transform 1 0 550620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5985
timestamp 1676037725
transform 1 0 551724 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5991
timestamp 1676037725
transform 1 0 552276 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5993
timestamp 1676037725
transform 1 0 552460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6005
timestamp 1676037725
transform 1 0 553564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6017
timestamp 1676037725
transform 1 0 554668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6029
timestamp 1676037725
transform 1 0 555772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6041
timestamp 1676037725
transform 1 0 556876 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6047
timestamp 1676037725
transform 1 0 557428 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6049
timestamp 1676037725
transform 1 0 557612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6061
timestamp 1676037725
transform 1 0 558716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6073
timestamp 1676037725
transform 1 0 559820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6085
timestamp 1676037725
transform 1 0 560924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6097
timestamp 1676037725
transform 1 0 562028 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6103
timestamp 1676037725
transform 1 0 562580 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6105
timestamp 1676037725
transform 1 0 562764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6117
timestamp 1676037725
transform 1 0 563868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6129
timestamp 1676037725
transform 1 0 564972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6141
timestamp 1676037725
transform 1 0 566076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6153
timestamp 1676037725
transform 1 0 567180 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6159
timestamp 1676037725
transform 1 0 567732 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6161
timestamp 1676037725
transform 1 0 567916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6173
timestamp 1676037725
transform 1 0 569020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6185
timestamp 1676037725
transform 1 0 570124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6197
timestamp 1676037725
transform 1 0 571228 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6209
timestamp 1676037725
transform 1 0 572332 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6215
timestamp 1676037725
transform 1 0 572884 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6217
timestamp 1676037725
transform 1 0 573068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6229
timestamp 1676037725
transform 1 0 574172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6241
timestamp 1676037725
transform 1 0 575276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6253
timestamp 1676037725
transform 1 0 576380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6265
timestamp 1676037725
transform 1 0 577484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6271
timestamp 1676037725
transform 1 0 578036 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6273
timestamp 1676037725
transform 1 0 578220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6285
timestamp 1676037725
transform 1 0 579324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6297
timestamp 1676037725
transform 1 0 580428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6309
timestamp 1676037725
transform 1 0 581532 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6321
timestamp 1676037725
transform 1 0 582636 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6327
timestamp 1676037725
transform 1 0 583188 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6329
timestamp 1676037725
transform 1 0 583372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6341
timestamp 1676037725
transform 1 0 584476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6353
timestamp 1676037725
transform 1 0 585580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6365
timestamp 1676037725
transform 1 0 586684 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6377
timestamp 1676037725
transform 1 0 587788 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6383
timestamp 1676037725
transform 1 0 588340 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6385
timestamp 1676037725
transform 1 0 588524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6397
timestamp 1676037725
transform 1 0 589628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6409
timestamp 1676037725
transform 1 0 590732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6421
timestamp 1676037725
transform 1 0 591836 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6433
timestamp 1676037725
transform 1 0 592940 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6439
timestamp 1676037725
transform 1 0 593492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6441
timestamp 1676037725
transform 1 0 593676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6453
timestamp 1676037725
transform 1 0 594780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6465
timestamp 1676037725
transform 1 0 595884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6477
timestamp 1676037725
transform 1 0 596988 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6489
timestamp 1676037725
transform 1 0 598092 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6495
timestamp 1676037725
transform 1 0 598644 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6497
timestamp 1676037725
transform 1 0 598828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6509
timestamp 1676037725
transform 1 0 599932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6521
timestamp 1676037725
transform 1 0 601036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6533
timestamp 1676037725
transform 1 0 602140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6545
timestamp 1676037725
transform 1 0 603244 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6551
timestamp 1676037725
transform 1 0 603796 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6553
timestamp 1676037725
transform 1 0 603980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6565
timestamp 1676037725
transform 1 0 605084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6577
timestamp 1676037725
transform 1 0 606188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6589
timestamp 1676037725
transform 1 0 607292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6601
timestamp 1676037725
transform 1 0 608396 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6607
timestamp 1676037725
transform 1 0 608948 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6609
timestamp 1676037725
transform 1 0 609132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6621
timestamp 1676037725
transform 1 0 610236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6633
timestamp 1676037725
transform 1 0 611340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6645
timestamp 1676037725
transform 1 0 612444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6657
timestamp 1676037725
transform 1 0 613548 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6663
timestamp 1676037725
transform 1 0 614100 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6665
timestamp 1676037725
transform 1 0 614284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6677
timestamp 1676037725
transform 1 0 615388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6689
timestamp 1676037725
transform 1 0 616492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6701
timestamp 1676037725
transform 1 0 617596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6713
timestamp 1676037725
transform 1 0 618700 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6719
timestamp 1676037725
transform 1 0 619252 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6721
timestamp 1676037725
transform 1 0 619436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6733
timestamp 1676037725
transform 1 0 620540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6745
timestamp 1676037725
transform 1 0 621644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6757
timestamp 1676037725
transform 1 0 622748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6769
timestamp 1676037725
transform 1 0 623852 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6775
timestamp 1676037725
transform 1 0 624404 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6777
timestamp 1676037725
transform 1 0 624588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6789
timestamp 1676037725
transform 1 0 625692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6801
timestamp 1676037725
transform 1 0 626796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6813
timestamp 1676037725
transform 1 0 627900 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6825
timestamp 1676037725
transform 1 0 629004 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6831
timestamp 1676037725
transform 1 0 629556 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6833
timestamp 1676037725
transform 1 0 629740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6845
timestamp 1676037725
transform 1 0 630844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6857
timestamp 1676037725
transform 1 0 631948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6869
timestamp 1676037725
transform 1 0 633052 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6881
timestamp 1676037725
transform 1 0 634156 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6887
timestamp 1676037725
transform 1 0 634708 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6889
timestamp 1676037725
transform 1 0 634892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6901
timestamp 1676037725
transform 1 0 635996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6913
timestamp 1676037725
transform 1 0 637100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6925
timestamp 1676037725
transform 1 0 638204 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6937
timestamp 1676037725
transform 1 0 639308 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6943
timestamp 1676037725
transform 1 0 639860 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6945
timestamp 1676037725
transform 1 0 640044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6957
timestamp 1676037725
transform 1 0 641148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6969
timestamp 1676037725
transform 1 0 642252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6981
timestamp 1676037725
transform 1 0 643356 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6993
timestamp 1676037725
transform 1 0 644460 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6999
timestamp 1676037725
transform 1 0 645012 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7001
timestamp 1676037725
transform 1 0 645196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7013
timestamp 1676037725
transform 1 0 646300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7025
timestamp 1676037725
transform 1 0 647404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7037
timestamp 1676037725
transform 1 0 648508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_7049
timestamp 1676037725
transform 1 0 649612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7055
timestamp 1676037725
transform 1 0 650164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7057
timestamp 1676037725
transform 1 0 650348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7069
timestamp 1676037725
transform 1 0 651452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7081
timestamp 1676037725
transform 1 0 652556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7093
timestamp 1676037725
transform 1 0 653660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_7105
timestamp 1676037725
transform 1 0 654764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7111
timestamp 1676037725
transform 1 0 655316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7113
timestamp 1676037725
transform 1 0 655500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7125
timestamp 1676037725
transform 1 0 656604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7137
timestamp 1676037725
transform 1 0 657708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7149
timestamp 1676037725
transform 1 0 658812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_7161
timestamp 1676037725
transform 1 0 659916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7167
timestamp 1676037725
transform 1 0 660468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7169
timestamp 1676037725
transform 1 0 660652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7181
timestamp 1676037725
transform 1 0 661756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7193
timestamp 1676037725
transform 1 0 662860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7205
timestamp 1676037725
transform 1 0 663964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_7217
timestamp 1676037725
transform 1 0 665068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7223
timestamp 1676037725
transform 1 0 665620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7225
timestamp 1676037725
transform 1 0 665804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7237
timestamp 1676037725
transform 1 0 666908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7249
timestamp 1676037725
transform 1 0 668012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7261
timestamp 1676037725
transform 1 0 669116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_7273
timestamp 1676037725
transform 1 0 670220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7279
timestamp 1676037725
transform 1 0 670772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7281
timestamp 1676037725
transform 1 0 670956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7293
timestamp 1676037725
transform 1 0 672060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7305
timestamp 1676037725
transform 1 0 673164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7317
timestamp 1676037725
transform 1 0 674268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_7329
timestamp 1676037725
transform 1 0 675372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7335
timestamp 1676037725
transform 1 0 675924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7337
timestamp 1676037725
transform 1 0 676108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7349
timestamp 1676037725
transform 1 0 677212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7361
timestamp 1676037725
transform 1 0 678316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7373
timestamp 1676037725
transform 1 0 679420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_7385
timestamp 1676037725
transform 1 0 680524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7391
timestamp 1676037725
transform 1 0 681076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7393
timestamp 1676037725
transform 1 0 681260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7405
timestamp 1676037725
transform 1 0 682364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1676037725
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1676037725
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1676037725
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1676037725
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1676037725
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1676037725
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1676037725
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1676037725
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1676037725
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1676037725
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1676037725
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1676037725
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1676037725
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1676037725
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1676037725
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1676037725
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1676037725
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1676037725
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1676037725
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1676037725
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1676037725
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1676037725
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1676037725
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1676037725
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1676037725
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1676037725
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1676037725
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1676037725
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1676037725
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1676037725
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1676037725
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1676037725
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1676037725
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1676037725
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1676037725
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1676037725
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1676037725
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1676037725
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1676037725
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1676037725
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1676037725
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1676037725
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1676037725
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1676037725
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1676037725
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1676037725
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1676037725
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1676037725
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1676037725
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1676037725
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1676037725
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1676037725
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1676037725
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1676037725
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1676037725
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1676037725
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1676037725
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1676037725
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1676037725
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1676037725
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1676037725
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1676037725
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1676037725
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1676037725
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1676037725
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1676037725
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1676037725
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1676037725
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1229
timestamp 1676037725
transform 1 0 114172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1241
timestamp 1676037725
transform 1 0 115276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1676037725
transform 1 0 116380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1676037725
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1261
timestamp 1676037725
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1273
timestamp 1676037725
transform 1 0 118220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1285
timestamp 1676037725
transform 1 0 119324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1297
timestamp 1676037725
transform 1 0 120428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1309
timestamp 1676037725
transform 1 0 121532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1315
timestamp 1676037725
transform 1 0 122084 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1317
timestamp 1676037725
transform 1 0 122268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1329
timestamp 1676037725
transform 1 0 123372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1341
timestamp 1676037725
transform 1 0 124476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1353
timestamp 1676037725
transform 1 0 125580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1365
timestamp 1676037725
transform 1 0 126684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1371
timestamp 1676037725
transform 1 0 127236 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1373
timestamp 1676037725
transform 1 0 127420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1385
timestamp 1676037725
transform 1 0 128524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1397
timestamp 1676037725
transform 1 0 129628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1409
timestamp 1676037725
transform 1 0 130732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1421
timestamp 1676037725
transform 1 0 131836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1427
timestamp 1676037725
transform 1 0 132388 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1429
timestamp 1676037725
transform 1 0 132572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1441
timestamp 1676037725
transform 1 0 133676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1453
timestamp 1676037725
transform 1 0 134780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1465
timestamp 1676037725
transform 1 0 135884 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1477
timestamp 1676037725
transform 1 0 136988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1483
timestamp 1676037725
transform 1 0 137540 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1485
timestamp 1676037725
transform 1 0 137724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1497
timestamp 1676037725
transform 1 0 138828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1509
timestamp 1676037725
transform 1 0 139932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1521
timestamp 1676037725
transform 1 0 141036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1533
timestamp 1676037725
transform 1 0 142140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1539
timestamp 1676037725
transform 1 0 142692 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1541
timestamp 1676037725
transform 1 0 142876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1553
timestamp 1676037725
transform 1 0 143980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1565
timestamp 1676037725
transform 1 0 145084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1577
timestamp 1676037725
transform 1 0 146188 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1589
timestamp 1676037725
transform 1 0 147292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1595
timestamp 1676037725
transform 1 0 147844 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1597
timestamp 1676037725
transform 1 0 148028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1609
timestamp 1676037725
transform 1 0 149132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1621
timestamp 1676037725
transform 1 0 150236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1633
timestamp 1676037725
transform 1 0 151340 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1645
timestamp 1676037725
transform 1 0 152444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1651
timestamp 1676037725
transform 1 0 152996 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1653
timestamp 1676037725
transform 1 0 153180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1665
timestamp 1676037725
transform 1 0 154284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1677
timestamp 1676037725
transform 1 0 155388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1689
timestamp 1676037725
transform 1 0 156492 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1701
timestamp 1676037725
transform 1 0 157596 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1707
timestamp 1676037725
transform 1 0 158148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1709
timestamp 1676037725
transform 1 0 158332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1721
timestamp 1676037725
transform 1 0 159436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1733
timestamp 1676037725
transform 1 0 160540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1745
timestamp 1676037725
transform 1 0 161644 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1757
timestamp 1676037725
transform 1 0 162748 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1763
timestamp 1676037725
transform 1 0 163300 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1765
timestamp 1676037725
transform 1 0 163484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1777
timestamp 1676037725
transform 1 0 164588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1789
timestamp 1676037725
transform 1 0 165692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1801
timestamp 1676037725
transform 1 0 166796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1813
timestamp 1676037725
transform 1 0 167900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1819
timestamp 1676037725
transform 1 0 168452 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1821
timestamp 1676037725
transform 1 0 168636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1833
timestamp 1676037725
transform 1 0 169740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1845
timestamp 1676037725
transform 1 0 170844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1857
timestamp 1676037725
transform 1 0 171948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1869
timestamp 1676037725
transform 1 0 173052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1875
timestamp 1676037725
transform 1 0 173604 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1877
timestamp 1676037725
transform 1 0 173788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1889
timestamp 1676037725
transform 1 0 174892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1901
timestamp 1676037725
transform 1 0 175996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1913
timestamp 1676037725
transform 1 0 177100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1925
timestamp 1676037725
transform 1 0 178204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1931
timestamp 1676037725
transform 1 0 178756 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1933
timestamp 1676037725
transform 1 0 178940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1945
timestamp 1676037725
transform 1 0 180044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1957
timestamp 1676037725
transform 1 0 181148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1969
timestamp 1676037725
transform 1 0 182252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1981
timestamp 1676037725
transform 1 0 183356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1987
timestamp 1676037725
transform 1 0 183908 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1989
timestamp 1676037725
transform 1 0 184092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2001
timestamp 1676037725
transform 1 0 185196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2013
timestamp 1676037725
transform 1 0 186300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2025
timestamp 1676037725
transform 1 0 187404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2037
timestamp 1676037725
transform 1 0 188508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2043
timestamp 1676037725
transform 1 0 189060 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2045
timestamp 1676037725
transform 1 0 189244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2057
timestamp 1676037725
transform 1 0 190348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2069
timestamp 1676037725
transform 1 0 191452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2081
timestamp 1676037725
transform 1 0 192556 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2093
timestamp 1676037725
transform 1 0 193660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2099
timestamp 1676037725
transform 1 0 194212 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2101
timestamp 1676037725
transform 1 0 194396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2113
timestamp 1676037725
transform 1 0 195500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2125
timestamp 1676037725
transform 1 0 196604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2137
timestamp 1676037725
transform 1 0 197708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2149
timestamp 1676037725
transform 1 0 198812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2155
timestamp 1676037725
transform 1 0 199364 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2157
timestamp 1676037725
transform 1 0 199548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2169
timestamp 1676037725
transform 1 0 200652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2181
timestamp 1676037725
transform 1 0 201756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2193
timestamp 1676037725
transform 1 0 202860 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2205
timestamp 1676037725
transform 1 0 203964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2211
timestamp 1676037725
transform 1 0 204516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2213
timestamp 1676037725
transform 1 0 204700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2225
timestamp 1676037725
transform 1 0 205804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2237
timestamp 1676037725
transform 1 0 206908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2249
timestamp 1676037725
transform 1 0 208012 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2261
timestamp 1676037725
transform 1 0 209116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2267
timestamp 1676037725
transform 1 0 209668 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2269
timestamp 1676037725
transform 1 0 209852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2281
timestamp 1676037725
transform 1 0 210956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2293
timestamp 1676037725
transform 1 0 212060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2305
timestamp 1676037725
transform 1 0 213164 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2317
timestamp 1676037725
transform 1 0 214268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2323
timestamp 1676037725
transform 1 0 214820 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2325
timestamp 1676037725
transform 1 0 215004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2337
timestamp 1676037725
transform 1 0 216108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2349
timestamp 1676037725
transform 1 0 217212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2361
timestamp 1676037725
transform 1 0 218316 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2373
timestamp 1676037725
transform 1 0 219420 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2379
timestamp 1676037725
transform 1 0 219972 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2381
timestamp 1676037725
transform 1 0 220156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2393
timestamp 1676037725
transform 1 0 221260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2405
timestamp 1676037725
transform 1 0 222364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2417
timestamp 1676037725
transform 1 0 223468 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2429
timestamp 1676037725
transform 1 0 224572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2435
timestamp 1676037725
transform 1 0 225124 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2437
timestamp 1676037725
transform 1 0 225308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2449
timestamp 1676037725
transform 1 0 226412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2461
timestamp 1676037725
transform 1 0 227516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2473
timestamp 1676037725
transform 1 0 228620 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2485
timestamp 1676037725
transform 1 0 229724 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2491
timestamp 1676037725
transform 1 0 230276 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2493
timestamp 1676037725
transform 1 0 230460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2505
timestamp 1676037725
transform 1 0 231564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2517
timestamp 1676037725
transform 1 0 232668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2529
timestamp 1676037725
transform 1 0 233772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2541
timestamp 1676037725
transform 1 0 234876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2547
timestamp 1676037725
transform 1 0 235428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2549
timestamp 1676037725
transform 1 0 235612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2561
timestamp 1676037725
transform 1 0 236716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2573
timestamp 1676037725
transform 1 0 237820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2585
timestamp 1676037725
transform 1 0 238924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2597
timestamp 1676037725
transform 1 0 240028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2603
timestamp 1676037725
transform 1 0 240580 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2605
timestamp 1676037725
transform 1 0 240764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2617
timestamp 1676037725
transform 1 0 241868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2629
timestamp 1676037725
transform 1 0 242972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2641
timestamp 1676037725
transform 1 0 244076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2653
timestamp 1676037725
transform 1 0 245180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2659
timestamp 1676037725
transform 1 0 245732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2661
timestamp 1676037725
transform 1 0 245916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2673
timestamp 1676037725
transform 1 0 247020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2685
timestamp 1676037725
transform 1 0 248124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2697
timestamp 1676037725
transform 1 0 249228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2709
timestamp 1676037725
transform 1 0 250332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2715
timestamp 1676037725
transform 1 0 250884 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2717
timestamp 1676037725
transform 1 0 251068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2729
timestamp 1676037725
transform 1 0 252172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2741
timestamp 1676037725
transform 1 0 253276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2753
timestamp 1676037725
transform 1 0 254380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2765
timestamp 1676037725
transform 1 0 255484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2771
timestamp 1676037725
transform 1 0 256036 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2773
timestamp 1676037725
transform 1 0 256220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2785
timestamp 1676037725
transform 1 0 257324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2797
timestamp 1676037725
transform 1 0 258428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2809
timestamp 1676037725
transform 1 0 259532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2821
timestamp 1676037725
transform 1 0 260636 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2827
timestamp 1676037725
transform 1 0 261188 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2829
timestamp 1676037725
transform 1 0 261372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2841
timestamp 1676037725
transform 1 0 262476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2853
timestamp 1676037725
transform 1 0 263580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2865
timestamp 1676037725
transform 1 0 264684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2877
timestamp 1676037725
transform 1 0 265788 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2883
timestamp 1676037725
transform 1 0 266340 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2885
timestamp 1676037725
transform 1 0 266524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2897
timestamp 1676037725
transform 1 0 267628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2909
timestamp 1676037725
transform 1 0 268732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2921
timestamp 1676037725
transform 1 0 269836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2933
timestamp 1676037725
transform 1 0 270940 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2939
timestamp 1676037725
transform 1 0 271492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2941
timestamp 1676037725
transform 1 0 271676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2953
timestamp 1676037725
transform 1 0 272780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2965
timestamp 1676037725
transform 1 0 273884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2977
timestamp 1676037725
transform 1 0 274988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2989
timestamp 1676037725
transform 1 0 276092 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2995
timestamp 1676037725
transform 1 0 276644 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2997
timestamp 1676037725
transform 1 0 276828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3009
timestamp 1676037725
transform 1 0 277932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3021
timestamp 1676037725
transform 1 0 279036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3033
timestamp 1676037725
transform 1 0 280140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3045
timestamp 1676037725
transform 1 0 281244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3051
timestamp 1676037725
transform 1 0 281796 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3053
timestamp 1676037725
transform 1 0 281980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3065
timestamp 1676037725
transform 1 0 283084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3077
timestamp 1676037725
transform 1 0 284188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3089
timestamp 1676037725
transform 1 0 285292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3101
timestamp 1676037725
transform 1 0 286396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3107
timestamp 1676037725
transform 1 0 286948 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3109
timestamp 1676037725
transform 1 0 287132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3121
timestamp 1676037725
transform 1 0 288236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3133
timestamp 1676037725
transform 1 0 289340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3145
timestamp 1676037725
transform 1 0 290444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3157
timestamp 1676037725
transform 1 0 291548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3163
timestamp 1676037725
transform 1 0 292100 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3165
timestamp 1676037725
transform 1 0 292284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3177
timestamp 1676037725
transform 1 0 293388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3189
timestamp 1676037725
transform 1 0 294492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3201
timestamp 1676037725
transform 1 0 295596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3213
timestamp 1676037725
transform 1 0 296700 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3219
timestamp 1676037725
transform 1 0 297252 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3221
timestamp 1676037725
transform 1 0 297436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3233
timestamp 1676037725
transform 1 0 298540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3245
timestamp 1676037725
transform 1 0 299644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3257
timestamp 1676037725
transform 1 0 300748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3269
timestamp 1676037725
transform 1 0 301852 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3275
timestamp 1676037725
transform 1 0 302404 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3277
timestamp 1676037725
transform 1 0 302588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3289
timestamp 1676037725
transform 1 0 303692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3301
timestamp 1676037725
transform 1 0 304796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3313
timestamp 1676037725
transform 1 0 305900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3325
timestamp 1676037725
transform 1 0 307004 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3331
timestamp 1676037725
transform 1 0 307556 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3333
timestamp 1676037725
transform 1 0 307740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3345
timestamp 1676037725
transform 1 0 308844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3357
timestamp 1676037725
transform 1 0 309948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3369
timestamp 1676037725
transform 1 0 311052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3381
timestamp 1676037725
transform 1 0 312156 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3387
timestamp 1676037725
transform 1 0 312708 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3389
timestamp 1676037725
transform 1 0 312892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3401
timestamp 1676037725
transform 1 0 313996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3413
timestamp 1676037725
transform 1 0 315100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3425
timestamp 1676037725
transform 1 0 316204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3437
timestamp 1676037725
transform 1 0 317308 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3443
timestamp 1676037725
transform 1 0 317860 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3445
timestamp 1676037725
transform 1 0 318044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3457
timestamp 1676037725
transform 1 0 319148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3469
timestamp 1676037725
transform 1 0 320252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3481
timestamp 1676037725
transform 1 0 321356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3493
timestamp 1676037725
transform 1 0 322460 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3499
timestamp 1676037725
transform 1 0 323012 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3501
timestamp 1676037725
transform 1 0 323196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3513
timestamp 1676037725
transform 1 0 324300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3525
timestamp 1676037725
transform 1 0 325404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3537
timestamp 1676037725
transform 1 0 326508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3549
timestamp 1676037725
transform 1 0 327612 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3555
timestamp 1676037725
transform 1 0 328164 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3557
timestamp 1676037725
transform 1 0 328348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3569
timestamp 1676037725
transform 1 0 329452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3581
timestamp 1676037725
transform 1 0 330556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3593
timestamp 1676037725
transform 1 0 331660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3605
timestamp 1676037725
transform 1 0 332764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3611
timestamp 1676037725
transform 1 0 333316 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3613
timestamp 1676037725
transform 1 0 333500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3625
timestamp 1676037725
transform 1 0 334604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3637
timestamp 1676037725
transform 1 0 335708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3649
timestamp 1676037725
transform 1 0 336812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3661
timestamp 1676037725
transform 1 0 337916 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3667
timestamp 1676037725
transform 1 0 338468 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3669
timestamp 1676037725
transform 1 0 338652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3681
timestamp 1676037725
transform 1 0 339756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3693
timestamp 1676037725
transform 1 0 340860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3705
timestamp 1676037725
transform 1 0 341964 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3717
timestamp 1676037725
transform 1 0 343068 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3723
timestamp 1676037725
transform 1 0 343620 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3725
timestamp 1676037725
transform 1 0 343804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3737
timestamp 1676037725
transform 1 0 344908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3749
timestamp 1676037725
transform 1 0 346012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3761
timestamp 1676037725
transform 1 0 347116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3773
timestamp 1676037725
transform 1 0 348220 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3779
timestamp 1676037725
transform 1 0 348772 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3781
timestamp 1676037725
transform 1 0 348956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3793
timestamp 1676037725
transform 1 0 350060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3805
timestamp 1676037725
transform 1 0 351164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3817
timestamp 1676037725
transform 1 0 352268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3829
timestamp 1676037725
transform 1 0 353372 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3835
timestamp 1676037725
transform 1 0 353924 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3837
timestamp 1676037725
transform 1 0 354108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3849
timestamp 1676037725
transform 1 0 355212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3861
timestamp 1676037725
transform 1 0 356316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3873
timestamp 1676037725
transform 1 0 357420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3885
timestamp 1676037725
transform 1 0 358524 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3891
timestamp 1676037725
transform 1 0 359076 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3893
timestamp 1676037725
transform 1 0 359260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3905
timestamp 1676037725
transform 1 0 360364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3917
timestamp 1676037725
transform 1 0 361468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3929
timestamp 1676037725
transform 1 0 362572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3941
timestamp 1676037725
transform 1 0 363676 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3947
timestamp 1676037725
transform 1 0 364228 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3949
timestamp 1676037725
transform 1 0 364412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3961
timestamp 1676037725
transform 1 0 365516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3973
timestamp 1676037725
transform 1 0 366620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3985
timestamp 1676037725
transform 1 0 367724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3997
timestamp 1676037725
transform 1 0 368828 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4003
timestamp 1676037725
transform 1 0 369380 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4005
timestamp 1676037725
transform 1 0 369564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4017
timestamp 1676037725
transform 1 0 370668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4029
timestamp 1676037725
transform 1 0 371772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4041
timestamp 1676037725
transform 1 0 372876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4053
timestamp 1676037725
transform 1 0 373980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4059
timestamp 1676037725
transform 1 0 374532 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4061
timestamp 1676037725
transform 1 0 374716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4073
timestamp 1676037725
transform 1 0 375820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4085
timestamp 1676037725
transform 1 0 376924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4097
timestamp 1676037725
transform 1 0 378028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4109
timestamp 1676037725
transform 1 0 379132 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4115
timestamp 1676037725
transform 1 0 379684 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4117
timestamp 1676037725
transform 1 0 379868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4129
timestamp 1676037725
transform 1 0 380972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4141
timestamp 1676037725
transform 1 0 382076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4153
timestamp 1676037725
transform 1 0 383180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4165
timestamp 1676037725
transform 1 0 384284 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4171
timestamp 1676037725
transform 1 0 384836 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4173
timestamp 1676037725
transform 1 0 385020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4185
timestamp 1676037725
transform 1 0 386124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4197
timestamp 1676037725
transform 1 0 387228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4209
timestamp 1676037725
transform 1 0 388332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4221
timestamp 1676037725
transform 1 0 389436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4227
timestamp 1676037725
transform 1 0 389988 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4229
timestamp 1676037725
transform 1 0 390172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4241
timestamp 1676037725
transform 1 0 391276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4253
timestamp 1676037725
transform 1 0 392380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4265
timestamp 1676037725
transform 1 0 393484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4277
timestamp 1676037725
transform 1 0 394588 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4283
timestamp 1676037725
transform 1 0 395140 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4285
timestamp 1676037725
transform 1 0 395324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4297
timestamp 1676037725
transform 1 0 396428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4309
timestamp 1676037725
transform 1 0 397532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4321
timestamp 1676037725
transform 1 0 398636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4333
timestamp 1676037725
transform 1 0 399740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4339
timestamp 1676037725
transform 1 0 400292 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4341
timestamp 1676037725
transform 1 0 400476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4353
timestamp 1676037725
transform 1 0 401580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4365
timestamp 1676037725
transform 1 0 402684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4377
timestamp 1676037725
transform 1 0 403788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4389
timestamp 1676037725
transform 1 0 404892 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4395
timestamp 1676037725
transform 1 0 405444 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4397
timestamp 1676037725
transform 1 0 405628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4409
timestamp 1676037725
transform 1 0 406732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4421
timestamp 1676037725
transform 1 0 407836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4433
timestamp 1676037725
transform 1 0 408940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4445
timestamp 1676037725
transform 1 0 410044 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4451
timestamp 1676037725
transform 1 0 410596 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4453
timestamp 1676037725
transform 1 0 410780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4465
timestamp 1676037725
transform 1 0 411884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4477
timestamp 1676037725
transform 1 0 412988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4489
timestamp 1676037725
transform 1 0 414092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4501
timestamp 1676037725
transform 1 0 415196 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4507
timestamp 1676037725
transform 1 0 415748 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4509
timestamp 1676037725
transform 1 0 415932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4521
timestamp 1676037725
transform 1 0 417036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4533
timestamp 1676037725
transform 1 0 418140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4545
timestamp 1676037725
transform 1 0 419244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4557
timestamp 1676037725
transform 1 0 420348 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4563
timestamp 1676037725
transform 1 0 420900 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4565
timestamp 1676037725
transform 1 0 421084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4577
timestamp 1676037725
transform 1 0 422188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4589
timestamp 1676037725
transform 1 0 423292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4601
timestamp 1676037725
transform 1 0 424396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4613
timestamp 1676037725
transform 1 0 425500 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4619
timestamp 1676037725
transform 1 0 426052 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4621
timestamp 1676037725
transform 1 0 426236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4633
timestamp 1676037725
transform 1 0 427340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4645
timestamp 1676037725
transform 1 0 428444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4657
timestamp 1676037725
transform 1 0 429548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4669
timestamp 1676037725
transform 1 0 430652 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4675
timestamp 1676037725
transform 1 0 431204 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4677
timestamp 1676037725
transform 1 0 431388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4689
timestamp 1676037725
transform 1 0 432492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4701
timestamp 1676037725
transform 1 0 433596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4713
timestamp 1676037725
transform 1 0 434700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4725
timestamp 1676037725
transform 1 0 435804 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4731
timestamp 1676037725
transform 1 0 436356 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4733
timestamp 1676037725
transform 1 0 436540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4745
timestamp 1676037725
transform 1 0 437644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4757
timestamp 1676037725
transform 1 0 438748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4769
timestamp 1676037725
transform 1 0 439852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4781
timestamp 1676037725
transform 1 0 440956 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4787
timestamp 1676037725
transform 1 0 441508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4789
timestamp 1676037725
transform 1 0 441692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4801
timestamp 1676037725
transform 1 0 442796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4813
timestamp 1676037725
transform 1 0 443900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4825
timestamp 1676037725
transform 1 0 445004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4837
timestamp 1676037725
transform 1 0 446108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4843
timestamp 1676037725
transform 1 0 446660 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4845
timestamp 1676037725
transform 1 0 446844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4857
timestamp 1676037725
transform 1 0 447948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4869
timestamp 1676037725
transform 1 0 449052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4881
timestamp 1676037725
transform 1 0 450156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4893
timestamp 1676037725
transform 1 0 451260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4899
timestamp 1676037725
transform 1 0 451812 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4901
timestamp 1676037725
transform 1 0 451996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4913
timestamp 1676037725
transform 1 0 453100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4925
timestamp 1676037725
transform 1 0 454204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4937
timestamp 1676037725
transform 1 0 455308 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4949
timestamp 1676037725
transform 1 0 456412 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4955
timestamp 1676037725
transform 1 0 456964 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4957
timestamp 1676037725
transform 1 0 457148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4969
timestamp 1676037725
transform 1 0 458252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4981
timestamp 1676037725
transform 1 0 459356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4993
timestamp 1676037725
transform 1 0 460460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5005
timestamp 1676037725
transform 1 0 461564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5011
timestamp 1676037725
transform 1 0 462116 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5013
timestamp 1676037725
transform 1 0 462300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5025
timestamp 1676037725
transform 1 0 463404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5037
timestamp 1676037725
transform 1 0 464508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5049
timestamp 1676037725
transform 1 0 465612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5061
timestamp 1676037725
transform 1 0 466716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5067
timestamp 1676037725
transform 1 0 467268 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5069
timestamp 1676037725
transform 1 0 467452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5081
timestamp 1676037725
transform 1 0 468556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5093
timestamp 1676037725
transform 1 0 469660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5105
timestamp 1676037725
transform 1 0 470764 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5117
timestamp 1676037725
transform 1 0 471868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5123
timestamp 1676037725
transform 1 0 472420 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5125
timestamp 1676037725
transform 1 0 472604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5137
timestamp 1676037725
transform 1 0 473708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5149
timestamp 1676037725
transform 1 0 474812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5161
timestamp 1676037725
transform 1 0 475916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5173
timestamp 1676037725
transform 1 0 477020 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5179
timestamp 1676037725
transform 1 0 477572 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5181
timestamp 1676037725
transform 1 0 477756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5193
timestamp 1676037725
transform 1 0 478860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5205
timestamp 1676037725
transform 1 0 479964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5217
timestamp 1676037725
transform 1 0 481068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5229
timestamp 1676037725
transform 1 0 482172 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5235
timestamp 1676037725
transform 1 0 482724 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5237
timestamp 1676037725
transform 1 0 482908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5249
timestamp 1676037725
transform 1 0 484012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5261
timestamp 1676037725
transform 1 0 485116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5273
timestamp 1676037725
transform 1 0 486220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5285
timestamp 1676037725
transform 1 0 487324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5291
timestamp 1676037725
transform 1 0 487876 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5293
timestamp 1676037725
transform 1 0 488060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5305
timestamp 1676037725
transform 1 0 489164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5317
timestamp 1676037725
transform 1 0 490268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5329
timestamp 1676037725
transform 1 0 491372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5341
timestamp 1676037725
transform 1 0 492476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5347
timestamp 1676037725
transform 1 0 493028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5349
timestamp 1676037725
transform 1 0 493212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5361
timestamp 1676037725
transform 1 0 494316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5373
timestamp 1676037725
transform 1 0 495420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5385
timestamp 1676037725
transform 1 0 496524 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5397
timestamp 1676037725
transform 1 0 497628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5403
timestamp 1676037725
transform 1 0 498180 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5405
timestamp 1676037725
transform 1 0 498364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5417
timestamp 1676037725
transform 1 0 499468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5429
timestamp 1676037725
transform 1 0 500572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5441
timestamp 1676037725
transform 1 0 501676 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5453
timestamp 1676037725
transform 1 0 502780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5459
timestamp 1676037725
transform 1 0 503332 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5461
timestamp 1676037725
transform 1 0 503516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5473
timestamp 1676037725
transform 1 0 504620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5485
timestamp 1676037725
transform 1 0 505724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5497
timestamp 1676037725
transform 1 0 506828 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5509
timestamp 1676037725
transform 1 0 507932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5515
timestamp 1676037725
transform 1 0 508484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5517
timestamp 1676037725
transform 1 0 508668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5529
timestamp 1676037725
transform 1 0 509772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5541
timestamp 1676037725
transform 1 0 510876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5553
timestamp 1676037725
transform 1 0 511980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5565
timestamp 1676037725
transform 1 0 513084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5571
timestamp 1676037725
transform 1 0 513636 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5573
timestamp 1676037725
transform 1 0 513820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5585
timestamp 1676037725
transform 1 0 514924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5597
timestamp 1676037725
transform 1 0 516028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5609
timestamp 1676037725
transform 1 0 517132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5621
timestamp 1676037725
transform 1 0 518236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5627
timestamp 1676037725
transform 1 0 518788 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5629
timestamp 1676037725
transform 1 0 518972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5641
timestamp 1676037725
transform 1 0 520076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5653
timestamp 1676037725
transform 1 0 521180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5665
timestamp 1676037725
transform 1 0 522284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5677
timestamp 1676037725
transform 1 0 523388 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5683
timestamp 1676037725
transform 1 0 523940 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5685
timestamp 1676037725
transform 1 0 524124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5697
timestamp 1676037725
transform 1 0 525228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5709
timestamp 1676037725
transform 1 0 526332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5721
timestamp 1676037725
transform 1 0 527436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5733
timestamp 1676037725
transform 1 0 528540 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5739
timestamp 1676037725
transform 1 0 529092 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5741
timestamp 1676037725
transform 1 0 529276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5753
timestamp 1676037725
transform 1 0 530380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5765
timestamp 1676037725
transform 1 0 531484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5777
timestamp 1676037725
transform 1 0 532588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5789
timestamp 1676037725
transform 1 0 533692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5795
timestamp 1676037725
transform 1 0 534244 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5797
timestamp 1676037725
transform 1 0 534428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5809
timestamp 1676037725
transform 1 0 535532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5821
timestamp 1676037725
transform 1 0 536636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5833
timestamp 1676037725
transform 1 0 537740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5845
timestamp 1676037725
transform 1 0 538844 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5851
timestamp 1676037725
transform 1 0 539396 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5853
timestamp 1676037725
transform 1 0 539580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5865
timestamp 1676037725
transform 1 0 540684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5877
timestamp 1676037725
transform 1 0 541788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5889
timestamp 1676037725
transform 1 0 542892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5901
timestamp 1676037725
transform 1 0 543996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5907
timestamp 1676037725
transform 1 0 544548 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5909
timestamp 1676037725
transform 1 0 544732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5921
timestamp 1676037725
transform 1 0 545836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5933
timestamp 1676037725
transform 1 0 546940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5945
timestamp 1676037725
transform 1 0 548044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5957
timestamp 1676037725
transform 1 0 549148 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5963
timestamp 1676037725
transform 1 0 549700 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5965
timestamp 1676037725
transform 1 0 549884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5977
timestamp 1676037725
transform 1 0 550988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5989
timestamp 1676037725
transform 1 0 552092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6001
timestamp 1676037725
transform 1 0 553196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6013
timestamp 1676037725
transform 1 0 554300 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6019
timestamp 1676037725
transform 1 0 554852 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6021
timestamp 1676037725
transform 1 0 555036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6033
timestamp 1676037725
transform 1 0 556140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6045
timestamp 1676037725
transform 1 0 557244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6057
timestamp 1676037725
transform 1 0 558348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6069
timestamp 1676037725
transform 1 0 559452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6075
timestamp 1676037725
transform 1 0 560004 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6077
timestamp 1676037725
transform 1 0 560188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6089
timestamp 1676037725
transform 1 0 561292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6101
timestamp 1676037725
transform 1 0 562396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6113
timestamp 1676037725
transform 1 0 563500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6125
timestamp 1676037725
transform 1 0 564604 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6131
timestamp 1676037725
transform 1 0 565156 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6133
timestamp 1676037725
transform 1 0 565340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6145
timestamp 1676037725
transform 1 0 566444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6157
timestamp 1676037725
transform 1 0 567548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6169
timestamp 1676037725
transform 1 0 568652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6181
timestamp 1676037725
transform 1 0 569756 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6187
timestamp 1676037725
transform 1 0 570308 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6189
timestamp 1676037725
transform 1 0 570492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6201
timestamp 1676037725
transform 1 0 571596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6213
timestamp 1676037725
transform 1 0 572700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6225
timestamp 1676037725
transform 1 0 573804 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6237
timestamp 1676037725
transform 1 0 574908 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6243
timestamp 1676037725
transform 1 0 575460 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6245
timestamp 1676037725
transform 1 0 575644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6257
timestamp 1676037725
transform 1 0 576748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6269
timestamp 1676037725
transform 1 0 577852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6281
timestamp 1676037725
transform 1 0 578956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6293
timestamp 1676037725
transform 1 0 580060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6299
timestamp 1676037725
transform 1 0 580612 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6301
timestamp 1676037725
transform 1 0 580796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6313
timestamp 1676037725
transform 1 0 581900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6325
timestamp 1676037725
transform 1 0 583004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6337
timestamp 1676037725
transform 1 0 584108 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6349
timestamp 1676037725
transform 1 0 585212 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6355
timestamp 1676037725
transform 1 0 585764 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6357
timestamp 1676037725
transform 1 0 585948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6369
timestamp 1676037725
transform 1 0 587052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6381
timestamp 1676037725
transform 1 0 588156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6393
timestamp 1676037725
transform 1 0 589260 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6405
timestamp 1676037725
transform 1 0 590364 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6411
timestamp 1676037725
transform 1 0 590916 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6413
timestamp 1676037725
transform 1 0 591100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6425
timestamp 1676037725
transform 1 0 592204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6437
timestamp 1676037725
transform 1 0 593308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6449
timestamp 1676037725
transform 1 0 594412 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6461
timestamp 1676037725
transform 1 0 595516 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6467
timestamp 1676037725
transform 1 0 596068 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6469
timestamp 1676037725
transform 1 0 596252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6481
timestamp 1676037725
transform 1 0 597356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6493
timestamp 1676037725
transform 1 0 598460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6505
timestamp 1676037725
transform 1 0 599564 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6517
timestamp 1676037725
transform 1 0 600668 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6523
timestamp 1676037725
transform 1 0 601220 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6525
timestamp 1676037725
transform 1 0 601404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6537
timestamp 1676037725
transform 1 0 602508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6549
timestamp 1676037725
transform 1 0 603612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6561
timestamp 1676037725
transform 1 0 604716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6573
timestamp 1676037725
transform 1 0 605820 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6579
timestamp 1676037725
transform 1 0 606372 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6581
timestamp 1676037725
transform 1 0 606556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6593
timestamp 1676037725
transform 1 0 607660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6605
timestamp 1676037725
transform 1 0 608764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6617
timestamp 1676037725
transform 1 0 609868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6629
timestamp 1676037725
transform 1 0 610972 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6635
timestamp 1676037725
transform 1 0 611524 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6637
timestamp 1676037725
transform 1 0 611708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6649
timestamp 1676037725
transform 1 0 612812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6661
timestamp 1676037725
transform 1 0 613916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6673
timestamp 1676037725
transform 1 0 615020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6685
timestamp 1676037725
transform 1 0 616124 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6691
timestamp 1676037725
transform 1 0 616676 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6693
timestamp 1676037725
transform 1 0 616860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6705
timestamp 1676037725
transform 1 0 617964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6717
timestamp 1676037725
transform 1 0 619068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6729
timestamp 1676037725
transform 1 0 620172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6741
timestamp 1676037725
transform 1 0 621276 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6747
timestamp 1676037725
transform 1 0 621828 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6749
timestamp 1676037725
transform 1 0 622012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6761
timestamp 1676037725
transform 1 0 623116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6773
timestamp 1676037725
transform 1 0 624220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6785
timestamp 1676037725
transform 1 0 625324 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6797
timestamp 1676037725
transform 1 0 626428 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6803
timestamp 1676037725
transform 1 0 626980 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6805
timestamp 1676037725
transform 1 0 627164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6817
timestamp 1676037725
transform 1 0 628268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6829
timestamp 1676037725
transform 1 0 629372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6841
timestamp 1676037725
transform 1 0 630476 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6853
timestamp 1676037725
transform 1 0 631580 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6859
timestamp 1676037725
transform 1 0 632132 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6861
timestamp 1676037725
transform 1 0 632316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6873
timestamp 1676037725
transform 1 0 633420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6885
timestamp 1676037725
transform 1 0 634524 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6897
timestamp 1676037725
transform 1 0 635628 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6909
timestamp 1676037725
transform 1 0 636732 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6915
timestamp 1676037725
transform 1 0 637284 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6917
timestamp 1676037725
transform 1 0 637468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6929
timestamp 1676037725
transform 1 0 638572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6941
timestamp 1676037725
transform 1 0 639676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6953
timestamp 1676037725
transform 1 0 640780 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6965
timestamp 1676037725
transform 1 0 641884 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6971
timestamp 1676037725
transform 1 0 642436 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6973
timestamp 1676037725
transform 1 0 642620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6985
timestamp 1676037725
transform 1 0 643724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6997
timestamp 1676037725
transform 1 0 644828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7009
timestamp 1676037725
transform 1 0 645932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7021
timestamp 1676037725
transform 1 0 647036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7027
timestamp 1676037725
transform 1 0 647588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7029
timestamp 1676037725
transform 1 0 647772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7041
timestamp 1676037725
transform 1 0 648876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7053
timestamp 1676037725
transform 1 0 649980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7065
timestamp 1676037725
transform 1 0 651084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7077
timestamp 1676037725
transform 1 0 652188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7083
timestamp 1676037725
transform 1 0 652740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7085
timestamp 1676037725
transform 1 0 652924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7097
timestamp 1676037725
transform 1 0 654028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7109
timestamp 1676037725
transform 1 0 655132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7121
timestamp 1676037725
transform 1 0 656236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7133
timestamp 1676037725
transform 1 0 657340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7139
timestamp 1676037725
transform 1 0 657892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7141
timestamp 1676037725
transform 1 0 658076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7153
timestamp 1676037725
transform 1 0 659180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7165
timestamp 1676037725
transform 1 0 660284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7177
timestamp 1676037725
transform 1 0 661388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7189
timestamp 1676037725
transform 1 0 662492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7195
timestamp 1676037725
transform 1 0 663044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7197
timestamp 1676037725
transform 1 0 663228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7209
timestamp 1676037725
transform 1 0 664332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7221
timestamp 1676037725
transform 1 0 665436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7233
timestamp 1676037725
transform 1 0 666540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7245
timestamp 1676037725
transform 1 0 667644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7251
timestamp 1676037725
transform 1 0 668196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7253
timestamp 1676037725
transform 1 0 668380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7265
timestamp 1676037725
transform 1 0 669484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7277
timestamp 1676037725
transform 1 0 670588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7289
timestamp 1676037725
transform 1 0 671692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7301
timestamp 1676037725
transform 1 0 672796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7307
timestamp 1676037725
transform 1 0 673348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7309
timestamp 1676037725
transform 1 0 673532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7321
timestamp 1676037725
transform 1 0 674636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7333
timestamp 1676037725
transform 1 0 675740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7345
timestamp 1676037725
transform 1 0 676844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7357
timestamp 1676037725
transform 1 0 677948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7363
timestamp 1676037725
transform 1 0 678500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7365
timestamp 1676037725
transform 1 0 678684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7377
timestamp 1676037725
transform 1 0 679788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7389
timestamp 1676037725
transform 1 0 680892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7401
timestamp 1676037725
transform 1 0 681996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1676037725
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1676037725
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1676037725
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1676037725
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1676037725
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1676037725
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1676037725
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1676037725
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1676037725
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1676037725
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1676037725
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1676037725
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1676037725
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1676037725
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1676037725
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1676037725
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1676037725
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1676037725
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1676037725
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1676037725
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1676037725
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1676037725
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1676037725
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1676037725
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1676037725
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1676037725
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1676037725
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1676037725
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1676037725
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1676037725
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1676037725
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1676037725
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1676037725
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1676037725
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1676037725
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1676037725
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1676037725
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1676037725
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1676037725
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1676037725
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1676037725
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1676037725
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1676037725
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1676037725
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1676037725
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1676037725
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1676037725
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1676037725
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1676037725
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1676037725
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1676037725
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1676037725
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1676037725
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1676037725
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1676037725
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1676037725
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1676037725
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1676037725
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1676037725
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1676037725
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1676037725
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1676037725
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1676037725
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1189
timestamp 1676037725
transform 1 0 110492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1201
timestamp 1676037725
transform 1 0 111596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1213
timestamp 1676037725
transform 1 0 112700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1676037725
transform 1 0 113804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1676037725
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1233
timestamp 1676037725
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1245
timestamp 1676037725
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1257
timestamp 1676037725
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1269
timestamp 1676037725
transform 1 0 117852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1281
timestamp 1676037725
transform 1 0 118956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1287
timestamp 1676037725
transform 1 0 119508 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1289
timestamp 1676037725
transform 1 0 119692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1301
timestamp 1676037725
transform 1 0 120796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1313
timestamp 1676037725
transform 1 0 121900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1325
timestamp 1676037725
transform 1 0 123004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1337
timestamp 1676037725
transform 1 0 124108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1343
timestamp 1676037725
transform 1 0 124660 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1345
timestamp 1676037725
transform 1 0 124844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1357
timestamp 1676037725
transform 1 0 125948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1369
timestamp 1676037725
transform 1 0 127052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1381
timestamp 1676037725
transform 1 0 128156 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1393
timestamp 1676037725
transform 1 0 129260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1399
timestamp 1676037725
transform 1 0 129812 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1401
timestamp 1676037725
transform 1 0 129996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1413
timestamp 1676037725
transform 1 0 131100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1425
timestamp 1676037725
transform 1 0 132204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1437
timestamp 1676037725
transform 1 0 133308 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1449
timestamp 1676037725
transform 1 0 134412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1455
timestamp 1676037725
transform 1 0 134964 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1457
timestamp 1676037725
transform 1 0 135148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1469
timestamp 1676037725
transform 1 0 136252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1481
timestamp 1676037725
transform 1 0 137356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1493
timestamp 1676037725
transform 1 0 138460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1505
timestamp 1676037725
transform 1 0 139564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1511
timestamp 1676037725
transform 1 0 140116 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1513
timestamp 1676037725
transform 1 0 140300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1525
timestamp 1676037725
transform 1 0 141404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1537
timestamp 1676037725
transform 1 0 142508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1549
timestamp 1676037725
transform 1 0 143612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1561
timestamp 1676037725
transform 1 0 144716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1567
timestamp 1676037725
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1569
timestamp 1676037725
transform 1 0 145452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1581
timestamp 1676037725
transform 1 0 146556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1593
timestamp 1676037725
transform 1 0 147660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1605
timestamp 1676037725
transform 1 0 148764 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1617
timestamp 1676037725
transform 1 0 149868 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1623
timestamp 1676037725
transform 1 0 150420 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1625
timestamp 1676037725
transform 1 0 150604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1637
timestamp 1676037725
transform 1 0 151708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1649
timestamp 1676037725
transform 1 0 152812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1661
timestamp 1676037725
transform 1 0 153916 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1673
timestamp 1676037725
transform 1 0 155020 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1679
timestamp 1676037725
transform 1 0 155572 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1681
timestamp 1676037725
transform 1 0 155756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1693
timestamp 1676037725
transform 1 0 156860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1705
timestamp 1676037725
transform 1 0 157964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1717
timestamp 1676037725
transform 1 0 159068 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1729
timestamp 1676037725
transform 1 0 160172 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1735
timestamp 1676037725
transform 1 0 160724 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1737
timestamp 1676037725
transform 1 0 160908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1749
timestamp 1676037725
transform 1 0 162012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1761
timestamp 1676037725
transform 1 0 163116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1773
timestamp 1676037725
transform 1 0 164220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1785
timestamp 1676037725
transform 1 0 165324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1791
timestamp 1676037725
transform 1 0 165876 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1793
timestamp 1676037725
transform 1 0 166060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1805
timestamp 1676037725
transform 1 0 167164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1817
timestamp 1676037725
transform 1 0 168268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1829
timestamp 1676037725
transform 1 0 169372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1841
timestamp 1676037725
transform 1 0 170476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1847
timestamp 1676037725
transform 1 0 171028 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1849
timestamp 1676037725
transform 1 0 171212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1861
timestamp 1676037725
transform 1 0 172316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1873
timestamp 1676037725
transform 1 0 173420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1885
timestamp 1676037725
transform 1 0 174524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1897
timestamp 1676037725
transform 1 0 175628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1903
timestamp 1676037725
transform 1 0 176180 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1905
timestamp 1676037725
transform 1 0 176364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1917
timestamp 1676037725
transform 1 0 177468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1929
timestamp 1676037725
transform 1 0 178572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1941
timestamp 1676037725
transform 1 0 179676 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1953
timestamp 1676037725
transform 1 0 180780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1959
timestamp 1676037725
transform 1 0 181332 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1961
timestamp 1676037725
transform 1 0 181516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1973
timestamp 1676037725
transform 1 0 182620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1985
timestamp 1676037725
transform 1 0 183724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1997
timestamp 1676037725
transform 1 0 184828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2009
timestamp 1676037725
transform 1 0 185932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2015
timestamp 1676037725
transform 1 0 186484 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2017
timestamp 1676037725
transform 1 0 186668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2029
timestamp 1676037725
transform 1 0 187772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2041
timestamp 1676037725
transform 1 0 188876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2053
timestamp 1676037725
transform 1 0 189980 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2065
timestamp 1676037725
transform 1 0 191084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2071
timestamp 1676037725
transform 1 0 191636 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2073
timestamp 1676037725
transform 1 0 191820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2085
timestamp 1676037725
transform 1 0 192924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2097
timestamp 1676037725
transform 1 0 194028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2109
timestamp 1676037725
transform 1 0 195132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2121
timestamp 1676037725
transform 1 0 196236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2127
timestamp 1676037725
transform 1 0 196788 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2129
timestamp 1676037725
transform 1 0 196972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2141
timestamp 1676037725
transform 1 0 198076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2153
timestamp 1676037725
transform 1 0 199180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2165
timestamp 1676037725
transform 1 0 200284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2177
timestamp 1676037725
transform 1 0 201388 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2183
timestamp 1676037725
transform 1 0 201940 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2185
timestamp 1676037725
transform 1 0 202124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2197
timestamp 1676037725
transform 1 0 203228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2209
timestamp 1676037725
transform 1 0 204332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2221
timestamp 1676037725
transform 1 0 205436 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2233
timestamp 1676037725
transform 1 0 206540 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2239
timestamp 1676037725
transform 1 0 207092 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2241
timestamp 1676037725
transform 1 0 207276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2253
timestamp 1676037725
transform 1 0 208380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2265
timestamp 1676037725
transform 1 0 209484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2277
timestamp 1676037725
transform 1 0 210588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2289
timestamp 1676037725
transform 1 0 211692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2295
timestamp 1676037725
transform 1 0 212244 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2297
timestamp 1676037725
transform 1 0 212428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2309
timestamp 1676037725
transform 1 0 213532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2321
timestamp 1676037725
transform 1 0 214636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2333
timestamp 1676037725
transform 1 0 215740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2345
timestamp 1676037725
transform 1 0 216844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2351
timestamp 1676037725
transform 1 0 217396 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2353
timestamp 1676037725
transform 1 0 217580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2365
timestamp 1676037725
transform 1 0 218684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2377
timestamp 1676037725
transform 1 0 219788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2389
timestamp 1676037725
transform 1 0 220892 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2401
timestamp 1676037725
transform 1 0 221996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2407
timestamp 1676037725
transform 1 0 222548 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2409
timestamp 1676037725
transform 1 0 222732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2421
timestamp 1676037725
transform 1 0 223836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2433
timestamp 1676037725
transform 1 0 224940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2445
timestamp 1676037725
transform 1 0 226044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2457
timestamp 1676037725
transform 1 0 227148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2463
timestamp 1676037725
transform 1 0 227700 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2465
timestamp 1676037725
transform 1 0 227884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2477
timestamp 1676037725
transform 1 0 228988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2489
timestamp 1676037725
transform 1 0 230092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2501
timestamp 1676037725
transform 1 0 231196 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2513
timestamp 1676037725
transform 1 0 232300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2519
timestamp 1676037725
transform 1 0 232852 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2521
timestamp 1676037725
transform 1 0 233036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2533
timestamp 1676037725
transform 1 0 234140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2545
timestamp 1676037725
transform 1 0 235244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2557
timestamp 1676037725
transform 1 0 236348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2569
timestamp 1676037725
transform 1 0 237452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2575
timestamp 1676037725
transform 1 0 238004 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2577
timestamp 1676037725
transform 1 0 238188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2589
timestamp 1676037725
transform 1 0 239292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2601
timestamp 1676037725
transform 1 0 240396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2613
timestamp 1676037725
transform 1 0 241500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2625
timestamp 1676037725
transform 1 0 242604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2631
timestamp 1676037725
transform 1 0 243156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2633
timestamp 1676037725
transform 1 0 243340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2645
timestamp 1676037725
transform 1 0 244444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2657
timestamp 1676037725
transform 1 0 245548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2669
timestamp 1676037725
transform 1 0 246652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2681
timestamp 1676037725
transform 1 0 247756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2687
timestamp 1676037725
transform 1 0 248308 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2689
timestamp 1676037725
transform 1 0 248492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2701
timestamp 1676037725
transform 1 0 249596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2713
timestamp 1676037725
transform 1 0 250700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2725
timestamp 1676037725
transform 1 0 251804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2737
timestamp 1676037725
transform 1 0 252908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2743
timestamp 1676037725
transform 1 0 253460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2745
timestamp 1676037725
transform 1 0 253644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2757
timestamp 1676037725
transform 1 0 254748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2769
timestamp 1676037725
transform 1 0 255852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2781
timestamp 1676037725
transform 1 0 256956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2793
timestamp 1676037725
transform 1 0 258060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2799
timestamp 1676037725
transform 1 0 258612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2801
timestamp 1676037725
transform 1 0 258796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2813
timestamp 1676037725
transform 1 0 259900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2825
timestamp 1676037725
transform 1 0 261004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2837
timestamp 1676037725
transform 1 0 262108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2849
timestamp 1676037725
transform 1 0 263212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2855
timestamp 1676037725
transform 1 0 263764 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2857
timestamp 1676037725
transform 1 0 263948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2869
timestamp 1676037725
transform 1 0 265052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2881
timestamp 1676037725
transform 1 0 266156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2893
timestamp 1676037725
transform 1 0 267260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2905
timestamp 1676037725
transform 1 0 268364 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2911
timestamp 1676037725
transform 1 0 268916 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2913
timestamp 1676037725
transform 1 0 269100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2925
timestamp 1676037725
transform 1 0 270204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2937
timestamp 1676037725
transform 1 0 271308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2949
timestamp 1676037725
transform 1 0 272412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2961
timestamp 1676037725
transform 1 0 273516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2967
timestamp 1676037725
transform 1 0 274068 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2969
timestamp 1676037725
transform 1 0 274252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2981
timestamp 1676037725
transform 1 0 275356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2993
timestamp 1676037725
transform 1 0 276460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3005
timestamp 1676037725
transform 1 0 277564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3017
timestamp 1676037725
transform 1 0 278668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3023
timestamp 1676037725
transform 1 0 279220 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3025
timestamp 1676037725
transform 1 0 279404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3037
timestamp 1676037725
transform 1 0 280508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3049
timestamp 1676037725
transform 1 0 281612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3061
timestamp 1676037725
transform 1 0 282716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3073
timestamp 1676037725
transform 1 0 283820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3079
timestamp 1676037725
transform 1 0 284372 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3081
timestamp 1676037725
transform 1 0 284556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3093
timestamp 1676037725
transform 1 0 285660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3105
timestamp 1676037725
transform 1 0 286764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3117
timestamp 1676037725
transform 1 0 287868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3129
timestamp 1676037725
transform 1 0 288972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3135
timestamp 1676037725
transform 1 0 289524 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3137
timestamp 1676037725
transform 1 0 289708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3149
timestamp 1676037725
transform 1 0 290812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3161
timestamp 1676037725
transform 1 0 291916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3173
timestamp 1676037725
transform 1 0 293020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3185
timestamp 1676037725
transform 1 0 294124 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3191
timestamp 1676037725
transform 1 0 294676 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3193
timestamp 1676037725
transform 1 0 294860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3205
timestamp 1676037725
transform 1 0 295964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3217
timestamp 1676037725
transform 1 0 297068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3229
timestamp 1676037725
transform 1 0 298172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3241
timestamp 1676037725
transform 1 0 299276 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3247
timestamp 1676037725
transform 1 0 299828 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3249
timestamp 1676037725
transform 1 0 300012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3261
timestamp 1676037725
transform 1 0 301116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3273
timestamp 1676037725
transform 1 0 302220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3285
timestamp 1676037725
transform 1 0 303324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3297
timestamp 1676037725
transform 1 0 304428 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3303
timestamp 1676037725
transform 1 0 304980 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3305
timestamp 1676037725
transform 1 0 305164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3317
timestamp 1676037725
transform 1 0 306268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3329
timestamp 1676037725
transform 1 0 307372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3341
timestamp 1676037725
transform 1 0 308476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3353
timestamp 1676037725
transform 1 0 309580 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3359
timestamp 1676037725
transform 1 0 310132 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3361
timestamp 1676037725
transform 1 0 310316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3373
timestamp 1676037725
transform 1 0 311420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3385
timestamp 1676037725
transform 1 0 312524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3397
timestamp 1676037725
transform 1 0 313628 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3409
timestamp 1676037725
transform 1 0 314732 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3415
timestamp 1676037725
transform 1 0 315284 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3417
timestamp 1676037725
transform 1 0 315468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3429
timestamp 1676037725
transform 1 0 316572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3441
timestamp 1676037725
transform 1 0 317676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3453
timestamp 1676037725
transform 1 0 318780 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3465
timestamp 1676037725
transform 1 0 319884 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3471
timestamp 1676037725
transform 1 0 320436 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3473
timestamp 1676037725
transform 1 0 320620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3485
timestamp 1676037725
transform 1 0 321724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3497
timestamp 1676037725
transform 1 0 322828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3509
timestamp 1676037725
transform 1 0 323932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3521
timestamp 1676037725
transform 1 0 325036 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3527
timestamp 1676037725
transform 1 0 325588 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3529
timestamp 1676037725
transform 1 0 325772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3541
timestamp 1676037725
transform 1 0 326876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3553
timestamp 1676037725
transform 1 0 327980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3565
timestamp 1676037725
transform 1 0 329084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3577
timestamp 1676037725
transform 1 0 330188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3583
timestamp 1676037725
transform 1 0 330740 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3585
timestamp 1676037725
transform 1 0 330924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3597
timestamp 1676037725
transform 1 0 332028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3609
timestamp 1676037725
transform 1 0 333132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3621
timestamp 1676037725
transform 1 0 334236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3633
timestamp 1676037725
transform 1 0 335340 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3639
timestamp 1676037725
transform 1 0 335892 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3641
timestamp 1676037725
transform 1 0 336076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3653
timestamp 1676037725
transform 1 0 337180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3665
timestamp 1676037725
transform 1 0 338284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3677
timestamp 1676037725
transform 1 0 339388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3689
timestamp 1676037725
transform 1 0 340492 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3695
timestamp 1676037725
transform 1 0 341044 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3697
timestamp 1676037725
transform 1 0 341228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3709
timestamp 1676037725
transform 1 0 342332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3721
timestamp 1676037725
transform 1 0 343436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3733
timestamp 1676037725
transform 1 0 344540 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3745
timestamp 1676037725
transform 1 0 345644 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3751
timestamp 1676037725
transform 1 0 346196 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3753
timestamp 1676037725
transform 1 0 346380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3765
timestamp 1676037725
transform 1 0 347484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3777
timestamp 1676037725
transform 1 0 348588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3789
timestamp 1676037725
transform 1 0 349692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3801
timestamp 1676037725
transform 1 0 350796 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3807
timestamp 1676037725
transform 1 0 351348 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3809
timestamp 1676037725
transform 1 0 351532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3821
timestamp 1676037725
transform 1 0 352636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3833
timestamp 1676037725
transform 1 0 353740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3845
timestamp 1676037725
transform 1 0 354844 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3857
timestamp 1676037725
transform 1 0 355948 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3863
timestamp 1676037725
transform 1 0 356500 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3865
timestamp 1676037725
transform 1 0 356684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3877
timestamp 1676037725
transform 1 0 357788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3889
timestamp 1676037725
transform 1 0 358892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3901
timestamp 1676037725
transform 1 0 359996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3913
timestamp 1676037725
transform 1 0 361100 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3919
timestamp 1676037725
transform 1 0 361652 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3921
timestamp 1676037725
transform 1 0 361836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3933
timestamp 1676037725
transform 1 0 362940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3945
timestamp 1676037725
transform 1 0 364044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3957
timestamp 1676037725
transform 1 0 365148 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3969
timestamp 1676037725
transform 1 0 366252 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3975
timestamp 1676037725
transform 1 0 366804 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3977
timestamp 1676037725
transform 1 0 366988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3989
timestamp 1676037725
transform 1 0 368092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4001
timestamp 1676037725
transform 1 0 369196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4013
timestamp 1676037725
transform 1 0 370300 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4025
timestamp 1676037725
transform 1 0 371404 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4031
timestamp 1676037725
transform 1 0 371956 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4033
timestamp 1676037725
transform 1 0 372140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4045
timestamp 1676037725
transform 1 0 373244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4057
timestamp 1676037725
transform 1 0 374348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4069
timestamp 1676037725
transform 1 0 375452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4081
timestamp 1676037725
transform 1 0 376556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4087
timestamp 1676037725
transform 1 0 377108 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4089
timestamp 1676037725
transform 1 0 377292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4101
timestamp 1676037725
transform 1 0 378396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4113
timestamp 1676037725
transform 1 0 379500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4125
timestamp 1676037725
transform 1 0 380604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4137
timestamp 1676037725
transform 1 0 381708 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4143
timestamp 1676037725
transform 1 0 382260 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4145
timestamp 1676037725
transform 1 0 382444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4157
timestamp 1676037725
transform 1 0 383548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4169
timestamp 1676037725
transform 1 0 384652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4181
timestamp 1676037725
transform 1 0 385756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4193
timestamp 1676037725
transform 1 0 386860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4199
timestamp 1676037725
transform 1 0 387412 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4201
timestamp 1676037725
transform 1 0 387596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4213
timestamp 1676037725
transform 1 0 388700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4225
timestamp 1676037725
transform 1 0 389804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4237
timestamp 1676037725
transform 1 0 390908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4249
timestamp 1676037725
transform 1 0 392012 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4255
timestamp 1676037725
transform 1 0 392564 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4257
timestamp 1676037725
transform 1 0 392748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4269
timestamp 1676037725
transform 1 0 393852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4281
timestamp 1676037725
transform 1 0 394956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4293
timestamp 1676037725
transform 1 0 396060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4305
timestamp 1676037725
transform 1 0 397164 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4311
timestamp 1676037725
transform 1 0 397716 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4313
timestamp 1676037725
transform 1 0 397900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4325
timestamp 1676037725
transform 1 0 399004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4337
timestamp 1676037725
transform 1 0 400108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4349
timestamp 1676037725
transform 1 0 401212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4361
timestamp 1676037725
transform 1 0 402316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4367
timestamp 1676037725
transform 1 0 402868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4369
timestamp 1676037725
transform 1 0 403052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4381
timestamp 1676037725
transform 1 0 404156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4393
timestamp 1676037725
transform 1 0 405260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4405
timestamp 1676037725
transform 1 0 406364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4417
timestamp 1676037725
transform 1 0 407468 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4423
timestamp 1676037725
transform 1 0 408020 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4425
timestamp 1676037725
transform 1 0 408204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4437
timestamp 1676037725
transform 1 0 409308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4449
timestamp 1676037725
transform 1 0 410412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4461
timestamp 1676037725
transform 1 0 411516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4473
timestamp 1676037725
transform 1 0 412620 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4479
timestamp 1676037725
transform 1 0 413172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4481
timestamp 1676037725
transform 1 0 413356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4493
timestamp 1676037725
transform 1 0 414460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4505
timestamp 1676037725
transform 1 0 415564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4517
timestamp 1676037725
transform 1 0 416668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4529
timestamp 1676037725
transform 1 0 417772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4535
timestamp 1676037725
transform 1 0 418324 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4537
timestamp 1676037725
transform 1 0 418508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4549
timestamp 1676037725
transform 1 0 419612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4561
timestamp 1676037725
transform 1 0 420716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4573
timestamp 1676037725
transform 1 0 421820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4585
timestamp 1676037725
transform 1 0 422924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4591
timestamp 1676037725
transform 1 0 423476 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4593
timestamp 1676037725
transform 1 0 423660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4605
timestamp 1676037725
transform 1 0 424764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4617
timestamp 1676037725
transform 1 0 425868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4629
timestamp 1676037725
transform 1 0 426972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4641
timestamp 1676037725
transform 1 0 428076 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4647
timestamp 1676037725
transform 1 0 428628 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4649
timestamp 1676037725
transform 1 0 428812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4661
timestamp 1676037725
transform 1 0 429916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4673
timestamp 1676037725
transform 1 0 431020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4685
timestamp 1676037725
transform 1 0 432124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4697
timestamp 1676037725
transform 1 0 433228 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4703
timestamp 1676037725
transform 1 0 433780 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4705
timestamp 1676037725
transform 1 0 433964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4717
timestamp 1676037725
transform 1 0 435068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4729
timestamp 1676037725
transform 1 0 436172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4741
timestamp 1676037725
transform 1 0 437276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4753
timestamp 1676037725
transform 1 0 438380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4759
timestamp 1676037725
transform 1 0 438932 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4761
timestamp 1676037725
transform 1 0 439116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4773
timestamp 1676037725
transform 1 0 440220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4785
timestamp 1676037725
transform 1 0 441324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4797
timestamp 1676037725
transform 1 0 442428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4809
timestamp 1676037725
transform 1 0 443532 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4815
timestamp 1676037725
transform 1 0 444084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4817
timestamp 1676037725
transform 1 0 444268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4829
timestamp 1676037725
transform 1 0 445372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4841
timestamp 1676037725
transform 1 0 446476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4853
timestamp 1676037725
transform 1 0 447580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4865
timestamp 1676037725
transform 1 0 448684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4871
timestamp 1676037725
transform 1 0 449236 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4873
timestamp 1676037725
transform 1 0 449420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4885
timestamp 1676037725
transform 1 0 450524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4897
timestamp 1676037725
transform 1 0 451628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4909
timestamp 1676037725
transform 1 0 452732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4921
timestamp 1676037725
transform 1 0 453836 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4927
timestamp 1676037725
transform 1 0 454388 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4929
timestamp 1676037725
transform 1 0 454572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4941
timestamp 1676037725
transform 1 0 455676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4953
timestamp 1676037725
transform 1 0 456780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4965
timestamp 1676037725
transform 1 0 457884 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4977
timestamp 1676037725
transform 1 0 458988 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4983
timestamp 1676037725
transform 1 0 459540 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4985
timestamp 1676037725
transform 1 0 459724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4997
timestamp 1676037725
transform 1 0 460828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5009
timestamp 1676037725
transform 1 0 461932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5021
timestamp 1676037725
transform 1 0 463036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5033
timestamp 1676037725
transform 1 0 464140 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5039
timestamp 1676037725
transform 1 0 464692 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5041
timestamp 1676037725
transform 1 0 464876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5053
timestamp 1676037725
transform 1 0 465980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5065
timestamp 1676037725
transform 1 0 467084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5077
timestamp 1676037725
transform 1 0 468188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5089
timestamp 1676037725
transform 1 0 469292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5095
timestamp 1676037725
transform 1 0 469844 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5097
timestamp 1676037725
transform 1 0 470028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5109
timestamp 1676037725
transform 1 0 471132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5121
timestamp 1676037725
transform 1 0 472236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5133
timestamp 1676037725
transform 1 0 473340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5145
timestamp 1676037725
transform 1 0 474444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5151
timestamp 1676037725
transform 1 0 474996 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5153
timestamp 1676037725
transform 1 0 475180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5165
timestamp 1676037725
transform 1 0 476284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5177
timestamp 1676037725
transform 1 0 477388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5189
timestamp 1676037725
transform 1 0 478492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5201
timestamp 1676037725
transform 1 0 479596 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5207
timestamp 1676037725
transform 1 0 480148 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5209
timestamp 1676037725
transform 1 0 480332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5221
timestamp 1676037725
transform 1 0 481436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5233
timestamp 1676037725
transform 1 0 482540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5245
timestamp 1676037725
transform 1 0 483644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5257
timestamp 1676037725
transform 1 0 484748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5263
timestamp 1676037725
transform 1 0 485300 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5265
timestamp 1676037725
transform 1 0 485484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5277
timestamp 1676037725
transform 1 0 486588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5289
timestamp 1676037725
transform 1 0 487692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5301
timestamp 1676037725
transform 1 0 488796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5313
timestamp 1676037725
transform 1 0 489900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5319
timestamp 1676037725
transform 1 0 490452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5321
timestamp 1676037725
transform 1 0 490636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5333
timestamp 1676037725
transform 1 0 491740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5345
timestamp 1676037725
transform 1 0 492844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5357
timestamp 1676037725
transform 1 0 493948 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5369
timestamp 1676037725
transform 1 0 495052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5375
timestamp 1676037725
transform 1 0 495604 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5377
timestamp 1676037725
transform 1 0 495788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5389
timestamp 1676037725
transform 1 0 496892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5401
timestamp 1676037725
transform 1 0 497996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5413
timestamp 1676037725
transform 1 0 499100 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5425
timestamp 1676037725
transform 1 0 500204 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5431
timestamp 1676037725
transform 1 0 500756 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5433
timestamp 1676037725
transform 1 0 500940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5445
timestamp 1676037725
transform 1 0 502044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5457
timestamp 1676037725
transform 1 0 503148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5469
timestamp 1676037725
transform 1 0 504252 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5481
timestamp 1676037725
transform 1 0 505356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5487
timestamp 1676037725
transform 1 0 505908 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5489
timestamp 1676037725
transform 1 0 506092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5501
timestamp 1676037725
transform 1 0 507196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5513
timestamp 1676037725
transform 1 0 508300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5525
timestamp 1676037725
transform 1 0 509404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5537
timestamp 1676037725
transform 1 0 510508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5543
timestamp 1676037725
transform 1 0 511060 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5545
timestamp 1676037725
transform 1 0 511244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5557
timestamp 1676037725
transform 1 0 512348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5569
timestamp 1676037725
transform 1 0 513452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5581
timestamp 1676037725
transform 1 0 514556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5593
timestamp 1676037725
transform 1 0 515660 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5599
timestamp 1676037725
transform 1 0 516212 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5601
timestamp 1676037725
transform 1 0 516396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5613
timestamp 1676037725
transform 1 0 517500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5625
timestamp 1676037725
transform 1 0 518604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5637
timestamp 1676037725
transform 1 0 519708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5649
timestamp 1676037725
transform 1 0 520812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5655
timestamp 1676037725
transform 1 0 521364 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5657
timestamp 1676037725
transform 1 0 521548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5669
timestamp 1676037725
transform 1 0 522652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5681
timestamp 1676037725
transform 1 0 523756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5693
timestamp 1676037725
transform 1 0 524860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5705
timestamp 1676037725
transform 1 0 525964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5711
timestamp 1676037725
transform 1 0 526516 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5713
timestamp 1676037725
transform 1 0 526700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5725
timestamp 1676037725
transform 1 0 527804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5737
timestamp 1676037725
transform 1 0 528908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5749
timestamp 1676037725
transform 1 0 530012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5761
timestamp 1676037725
transform 1 0 531116 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5767
timestamp 1676037725
transform 1 0 531668 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5769
timestamp 1676037725
transform 1 0 531852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5781
timestamp 1676037725
transform 1 0 532956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5793
timestamp 1676037725
transform 1 0 534060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5805
timestamp 1676037725
transform 1 0 535164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5817
timestamp 1676037725
transform 1 0 536268 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5823
timestamp 1676037725
transform 1 0 536820 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5825
timestamp 1676037725
transform 1 0 537004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5837
timestamp 1676037725
transform 1 0 538108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5849
timestamp 1676037725
transform 1 0 539212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5861
timestamp 1676037725
transform 1 0 540316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5873
timestamp 1676037725
transform 1 0 541420 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5879
timestamp 1676037725
transform 1 0 541972 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5881
timestamp 1676037725
transform 1 0 542156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5893
timestamp 1676037725
transform 1 0 543260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5905
timestamp 1676037725
transform 1 0 544364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5917
timestamp 1676037725
transform 1 0 545468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5929
timestamp 1676037725
transform 1 0 546572 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5935
timestamp 1676037725
transform 1 0 547124 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5937
timestamp 1676037725
transform 1 0 547308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5949
timestamp 1676037725
transform 1 0 548412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5961
timestamp 1676037725
transform 1 0 549516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5973
timestamp 1676037725
transform 1 0 550620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5985
timestamp 1676037725
transform 1 0 551724 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5991
timestamp 1676037725
transform 1 0 552276 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5993
timestamp 1676037725
transform 1 0 552460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6005
timestamp 1676037725
transform 1 0 553564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6017
timestamp 1676037725
transform 1 0 554668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6029
timestamp 1676037725
transform 1 0 555772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6041
timestamp 1676037725
transform 1 0 556876 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6047
timestamp 1676037725
transform 1 0 557428 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6049
timestamp 1676037725
transform 1 0 557612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6061
timestamp 1676037725
transform 1 0 558716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6073
timestamp 1676037725
transform 1 0 559820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6085
timestamp 1676037725
transform 1 0 560924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6097
timestamp 1676037725
transform 1 0 562028 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6103
timestamp 1676037725
transform 1 0 562580 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6105
timestamp 1676037725
transform 1 0 562764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6117
timestamp 1676037725
transform 1 0 563868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6129
timestamp 1676037725
transform 1 0 564972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6141
timestamp 1676037725
transform 1 0 566076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6153
timestamp 1676037725
transform 1 0 567180 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6159
timestamp 1676037725
transform 1 0 567732 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6161
timestamp 1676037725
transform 1 0 567916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6173
timestamp 1676037725
transform 1 0 569020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6185
timestamp 1676037725
transform 1 0 570124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6197
timestamp 1676037725
transform 1 0 571228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6209
timestamp 1676037725
transform 1 0 572332 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6215
timestamp 1676037725
transform 1 0 572884 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6217
timestamp 1676037725
transform 1 0 573068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6229
timestamp 1676037725
transform 1 0 574172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6241
timestamp 1676037725
transform 1 0 575276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6253
timestamp 1676037725
transform 1 0 576380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6265
timestamp 1676037725
transform 1 0 577484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6271
timestamp 1676037725
transform 1 0 578036 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6273
timestamp 1676037725
transform 1 0 578220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6285
timestamp 1676037725
transform 1 0 579324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6297
timestamp 1676037725
transform 1 0 580428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6309
timestamp 1676037725
transform 1 0 581532 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6321
timestamp 1676037725
transform 1 0 582636 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6327
timestamp 1676037725
transform 1 0 583188 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6329
timestamp 1676037725
transform 1 0 583372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6341
timestamp 1676037725
transform 1 0 584476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6353
timestamp 1676037725
transform 1 0 585580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6365
timestamp 1676037725
transform 1 0 586684 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6377
timestamp 1676037725
transform 1 0 587788 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6383
timestamp 1676037725
transform 1 0 588340 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6385
timestamp 1676037725
transform 1 0 588524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6397
timestamp 1676037725
transform 1 0 589628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6409
timestamp 1676037725
transform 1 0 590732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6421
timestamp 1676037725
transform 1 0 591836 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6433
timestamp 1676037725
transform 1 0 592940 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6439
timestamp 1676037725
transform 1 0 593492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6441
timestamp 1676037725
transform 1 0 593676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6453
timestamp 1676037725
transform 1 0 594780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6465
timestamp 1676037725
transform 1 0 595884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6477
timestamp 1676037725
transform 1 0 596988 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6489
timestamp 1676037725
transform 1 0 598092 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6495
timestamp 1676037725
transform 1 0 598644 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6497
timestamp 1676037725
transform 1 0 598828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6509
timestamp 1676037725
transform 1 0 599932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6521
timestamp 1676037725
transform 1 0 601036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6533
timestamp 1676037725
transform 1 0 602140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6545
timestamp 1676037725
transform 1 0 603244 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6551
timestamp 1676037725
transform 1 0 603796 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6553
timestamp 1676037725
transform 1 0 603980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6565
timestamp 1676037725
transform 1 0 605084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6577
timestamp 1676037725
transform 1 0 606188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6589
timestamp 1676037725
transform 1 0 607292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6601
timestamp 1676037725
transform 1 0 608396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6607
timestamp 1676037725
transform 1 0 608948 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6609
timestamp 1676037725
transform 1 0 609132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6621
timestamp 1676037725
transform 1 0 610236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6633
timestamp 1676037725
transform 1 0 611340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6645
timestamp 1676037725
transform 1 0 612444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6657
timestamp 1676037725
transform 1 0 613548 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6663
timestamp 1676037725
transform 1 0 614100 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6665
timestamp 1676037725
transform 1 0 614284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6677
timestamp 1676037725
transform 1 0 615388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6689
timestamp 1676037725
transform 1 0 616492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6701
timestamp 1676037725
transform 1 0 617596 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6713
timestamp 1676037725
transform 1 0 618700 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6719
timestamp 1676037725
transform 1 0 619252 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6721
timestamp 1676037725
transform 1 0 619436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6733
timestamp 1676037725
transform 1 0 620540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6745
timestamp 1676037725
transform 1 0 621644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6757
timestamp 1676037725
transform 1 0 622748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6769
timestamp 1676037725
transform 1 0 623852 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6775
timestamp 1676037725
transform 1 0 624404 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6777
timestamp 1676037725
transform 1 0 624588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6789
timestamp 1676037725
transform 1 0 625692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6801
timestamp 1676037725
transform 1 0 626796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6813
timestamp 1676037725
transform 1 0 627900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6825
timestamp 1676037725
transform 1 0 629004 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6831
timestamp 1676037725
transform 1 0 629556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6833
timestamp 1676037725
transform 1 0 629740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6845
timestamp 1676037725
transform 1 0 630844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6857
timestamp 1676037725
transform 1 0 631948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6869
timestamp 1676037725
transform 1 0 633052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6881
timestamp 1676037725
transform 1 0 634156 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6887
timestamp 1676037725
transform 1 0 634708 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6889
timestamp 1676037725
transform 1 0 634892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6901
timestamp 1676037725
transform 1 0 635996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6913
timestamp 1676037725
transform 1 0 637100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6925
timestamp 1676037725
transform 1 0 638204 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6937
timestamp 1676037725
transform 1 0 639308 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6943
timestamp 1676037725
transform 1 0 639860 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6945
timestamp 1676037725
transform 1 0 640044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6957
timestamp 1676037725
transform 1 0 641148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6969
timestamp 1676037725
transform 1 0 642252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6981
timestamp 1676037725
transform 1 0 643356 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6993
timestamp 1676037725
transform 1 0 644460 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6999
timestamp 1676037725
transform 1 0 645012 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7001
timestamp 1676037725
transform 1 0 645196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7013
timestamp 1676037725
transform 1 0 646300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7025
timestamp 1676037725
transform 1 0 647404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7037
timestamp 1676037725
transform 1 0 648508 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_7049
timestamp 1676037725
transform 1 0 649612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7055
timestamp 1676037725
transform 1 0 650164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7057
timestamp 1676037725
transform 1 0 650348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7069
timestamp 1676037725
transform 1 0 651452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7081
timestamp 1676037725
transform 1 0 652556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7093
timestamp 1676037725
transform 1 0 653660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_7105
timestamp 1676037725
transform 1 0 654764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7111
timestamp 1676037725
transform 1 0 655316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7113
timestamp 1676037725
transform 1 0 655500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7125
timestamp 1676037725
transform 1 0 656604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7137
timestamp 1676037725
transform 1 0 657708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7149
timestamp 1676037725
transform 1 0 658812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_7161
timestamp 1676037725
transform 1 0 659916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7167
timestamp 1676037725
transform 1 0 660468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7169
timestamp 1676037725
transform 1 0 660652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7181
timestamp 1676037725
transform 1 0 661756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7193
timestamp 1676037725
transform 1 0 662860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7205
timestamp 1676037725
transform 1 0 663964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_7217
timestamp 1676037725
transform 1 0 665068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7223
timestamp 1676037725
transform 1 0 665620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7225
timestamp 1676037725
transform 1 0 665804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7237
timestamp 1676037725
transform 1 0 666908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7249
timestamp 1676037725
transform 1 0 668012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7261
timestamp 1676037725
transform 1 0 669116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_7273
timestamp 1676037725
transform 1 0 670220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7279
timestamp 1676037725
transform 1 0 670772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7281
timestamp 1676037725
transform 1 0 670956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7293
timestamp 1676037725
transform 1 0 672060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7305
timestamp 1676037725
transform 1 0 673164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7317
timestamp 1676037725
transform 1 0 674268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_7329
timestamp 1676037725
transform 1 0 675372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7335
timestamp 1676037725
transform 1 0 675924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7337
timestamp 1676037725
transform 1 0 676108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7349
timestamp 1676037725
transform 1 0 677212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7361
timestamp 1676037725
transform 1 0 678316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7373
timestamp 1676037725
transform 1 0 679420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_7385
timestamp 1676037725
transform 1 0 680524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7391
timestamp 1676037725
transform 1 0 681076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7393
timestamp 1676037725
transform 1 0 681260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7405
timestamp 1676037725
transform 1 0 682364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1676037725
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1676037725
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1676037725
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1676037725
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1676037725
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1676037725
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1676037725
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1676037725
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1676037725
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1676037725
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1676037725
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1676037725
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1676037725
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1676037725
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1676037725
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1676037725
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1676037725
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1676037725
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1676037725
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1676037725
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1676037725
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1676037725
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1676037725
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1676037725
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1676037725
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1676037725
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1676037725
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1676037725
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1676037725
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1676037725
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1676037725
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1676037725
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1676037725
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1676037725
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1676037725
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1676037725
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1676037725
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1676037725
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1676037725
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1676037725
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1676037725
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1676037725
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1676037725
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1676037725
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1676037725
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1676037725
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1676037725
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1676037725
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1676037725
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1676037725
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1676037725
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1676037725
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1676037725
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1676037725
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1676037725
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1676037725
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1676037725
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1676037725
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1676037725
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1676037725
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1161
timestamp 1676037725
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1676037725
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1185
timestamp 1676037725
transform 1 0 110124 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1676037725
transform 1 0 111228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1676037725
transform 1 0 111780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1205
timestamp 1676037725
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1217
timestamp 1676037725
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1229
timestamp 1676037725
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1241
timestamp 1676037725
transform 1 0 115276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1676037725
transform 1 0 116380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1676037725
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1261
timestamp 1676037725
transform 1 0 117116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1273
timestamp 1676037725
transform 1 0 118220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1285
timestamp 1676037725
transform 1 0 119324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1297
timestamp 1676037725
transform 1 0 120428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1309
timestamp 1676037725
transform 1 0 121532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1315
timestamp 1676037725
transform 1 0 122084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1317
timestamp 1676037725
transform 1 0 122268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1329
timestamp 1676037725
transform 1 0 123372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1341
timestamp 1676037725
transform 1 0 124476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1353
timestamp 1676037725
transform 1 0 125580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1365
timestamp 1676037725
transform 1 0 126684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1371
timestamp 1676037725
transform 1 0 127236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1373
timestamp 1676037725
transform 1 0 127420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1385
timestamp 1676037725
transform 1 0 128524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1397
timestamp 1676037725
transform 1 0 129628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1409
timestamp 1676037725
transform 1 0 130732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1421
timestamp 1676037725
transform 1 0 131836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1427
timestamp 1676037725
transform 1 0 132388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1429
timestamp 1676037725
transform 1 0 132572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1441
timestamp 1676037725
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1453
timestamp 1676037725
transform 1 0 134780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1465
timestamp 1676037725
transform 1 0 135884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1477
timestamp 1676037725
transform 1 0 136988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1483
timestamp 1676037725
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1485
timestamp 1676037725
transform 1 0 137724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1497
timestamp 1676037725
transform 1 0 138828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1509
timestamp 1676037725
transform 1 0 139932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1521
timestamp 1676037725
transform 1 0 141036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1533
timestamp 1676037725
transform 1 0 142140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1539
timestamp 1676037725
transform 1 0 142692 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1541
timestamp 1676037725
transform 1 0 142876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1553
timestamp 1676037725
transform 1 0 143980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1565
timestamp 1676037725
transform 1 0 145084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1577
timestamp 1676037725
transform 1 0 146188 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1589
timestamp 1676037725
transform 1 0 147292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1595
timestamp 1676037725
transform 1 0 147844 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1597
timestamp 1676037725
transform 1 0 148028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1609
timestamp 1676037725
transform 1 0 149132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1621
timestamp 1676037725
transform 1 0 150236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1633
timestamp 1676037725
transform 1 0 151340 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1645
timestamp 1676037725
transform 1 0 152444 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1651
timestamp 1676037725
transform 1 0 152996 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1653
timestamp 1676037725
transform 1 0 153180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1665
timestamp 1676037725
transform 1 0 154284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1677
timestamp 1676037725
transform 1 0 155388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1689
timestamp 1676037725
transform 1 0 156492 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1701
timestamp 1676037725
transform 1 0 157596 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1707
timestamp 1676037725
transform 1 0 158148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1709
timestamp 1676037725
transform 1 0 158332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1721
timestamp 1676037725
transform 1 0 159436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1733
timestamp 1676037725
transform 1 0 160540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1745
timestamp 1676037725
transform 1 0 161644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1757
timestamp 1676037725
transform 1 0 162748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1763
timestamp 1676037725
transform 1 0 163300 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1765
timestamp 1676037725
transform 1 0 163484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1777
timestamp 1676037725
transform 1 0 164588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1789
timestamp 1676037725
transform 1 0 165692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1801
timestamp 1676037725
transform 1 0 166796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1813
timestamp 1676037725
transform 1 0 167900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1819
timestamp 1676037725
transform 1 0 168452 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1821
timestamp 1676037725
transform 1 0 168636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1833
timestamp 1676037725
transform 1 0 169740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1845
timestamp 1676037725
transform 1 0 170844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1857
timestamp 1676037725
transform 1 0 171948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1869
timestamp 1676037725
transform 1 0 173052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1875
timestamp 1676037725
transform 1 0 173604 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1877
timestamp 1676037725
transform 1 0 173788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1889
timestamp 1676037725
transform 1 0 174892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1901
timestamp 1676037725
transform 1 0 175996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1913
timestamp 1676037725
transform 1 0 177100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1925
timestamp 1676037725
transform 1 0 178204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1931
timestamp 1676037725
transform 1 0 178756 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1933
timestamp 1676037725
transform 1 0 178940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1945
timestamp 1676037725
transform 1 0 180044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1957
timestamp 1676037725
transform 1 0 181148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1969
timestamp 1676037725
transform 1 0 182252 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1981
timestamp 1676037725
transform 1 0 183356 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1987
timestamp 1676037725
transform 1 0 183908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1989
timestamp 1676037725
transform 1 0 184092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2001
timestamp 1676037725
transform 1 0 185196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2013
timestamp 1676037725
transform 1 0 186300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2025
timestamp 1676037725
transform 1 0 187404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2037
timestamp 1676037725
transform 1 0 188508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2043
timestamp 1676037725
transform 1 0 189060 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2045
timestamp 1676037725
transform 1 0 189244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2057
timestamp 1676037725
transform 1 0 190348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2069
timestamp 1676037725
transform 1 0 191452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2081
timestamp 1676037725
transform 1 0 192556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2093
timestamp 1676037725
transform 1 0 193660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2099
timestamp 1676037725
transform 1 0 194212 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2101
timestamp 1676037725
transform 1 0 194396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2113
timestamp 1676037725
transform 1 0 195500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2125
timestamp 1676037725
transform 1 0 196604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2137
timestamp 1676037725
transform 1 0 197708 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2149
timestamp 1676037725
transform 1 0 198812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2155
timestamp 1676037725
transform 1 0 199364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2157
timestamp 1676037725
transform 1 0 199548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2169
timestamp 1676037725
transform 1 0 200652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2181
timestamp 1676037725
transform 1 0 201756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2193
timestamp 1676037725
transform 1 0 202860 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2205
timestamp 1676037725
transform 1 0 203964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2211
timestamp 1676037725
transform 1 0 204516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2213
timestamp 1676037725
transform 1 0 204700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2225
timestamp 1676037725
transform 1 0 205804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2237
timestamp 1676037725
transform 1 0 206908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2249
timestamp 1676037725
transform 1 0 208012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2261
timestamp 1676037725
transform 1 0 209116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2267
timestamp 1676037725
transform 1 0 209668 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2269
timestamp 1676037725
transform 1 0 209852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2281
timestamp 1676037725
transform 1 0 210956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2293
timestamp 1676037725
transform 1 0 212060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2305
timestamp 1676037725
transform 1 0 213164 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2317
timestamp 1676037725
transform 1 0 214268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2323
timestamp 1676037725
transform 1 0 214820 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2325
timestamp 1676037725
transform 1 0 215004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2337
timestamp 1676037725
transform 1 0 216108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2349
timestamp 1676037725
transform 1 0 217212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2361
timestamp 1676037725
transform 1 0 218316 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2373
timestamp 1676037725
transform 1 0 219420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2379
timestamp 1676037725
transform 1 0 219972 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2381
timestamp 1676037725
transform 1 0 220156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2393
timestamp 1676037725
transform 1 0 221260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2405
timestamp 1676037725
transform 1 0 222364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2417
timestamp 1676037725
transform 1 0 223468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2429
timestamp 1676037725
transform 1 0 224572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2435
timestamp 1676037725
transform 1 0 225124 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2437
timestamp 1676037725
transform 1 0 225308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2449
timestamp 1676037725
transform 1 0 226412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2461
timestamp 1676037725
transform 1 0 227516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2473
timestamp 1676037725
transform 1 0 228620 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2485
timestamp 1676037725
transform 1 0 229724 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2491
timestamp 1676037725
transform 1 0 230276 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2493
timestamp 1676037725
transform 1 0 230460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2505
timestamp 1676037725
transform 1 0 231564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2517
timestamp 1676037725
transform 1 0 232668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2529
timestamp 1676037725
transform 1 0 233772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2541
timestamp 1676037725
transform 1 0 234876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2547
timestamp 1676037725
transform 1 0 235428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2549
timestamp 1676037725
transform 1 0 235612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2561
timestamp 1676037725
transform 1 0 236716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2573
timestamp 1676037725
transform 1 0 237820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2585
timestamp 1676037725
transform 1 0 238924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2597
timestamp 1676037725
transform 1 0 240028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2603
timestamp 1676037725
transform 1 0 240580 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2605
timestamp 1676037725
transform 1 0 240764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2617
timestamp 1676037725
transform 1 0 241868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2629
timestamp 1676037725
transform 1 0 242972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2641
timestamp 1676037725
transform 1 0 244076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2653
timestamp 1676037725
transform 1 0 245180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2659
timestamp 1676037725
transform 1 0 245732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2661
timestamp 1676037725
transform 1 0 245916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2673
timestamp 1676037725
transform 1 0 247020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2685
timestamp 1676037725
transform 1 0 248124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2697
timestamp 1676037725
transform 1 0 249228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2709
timestamp 1676037725
transform 1 0 250332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2715
timestamp 1676037725
transform 1 0 250884 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2717
timestamp 1676037725
transform 1 0 251068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2729
timestamp 1676037725
transform 1 0 252172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2741
timestamp 1676037725
transform 1 0 253276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2753
timestamp 1676037725
transform 1 0 254380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2765
timestamp 1676037725
transform 1 0 255484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2771
timestamp 1676037725
transform 1 0 256036 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2773
timestamp 1676037725
transform 1 0 256220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2785
timestamp 1676037725
transform 1 0 257324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2797
timestamp 1676037725
transform 1 0 258428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2809
timestamp 1676037725
transform 1 0 259532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2821
timestamp 1676037725
transform 1 0 260636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2827
timestamp 1676037725
transform 1 0 261188 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2829
timestamp 1676037725
transform 1 0 261372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2841
timestamp 1676037725
transform 1 0 262476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2853
timestamp 1676037725
transform 1 0 263580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2865
timestamp 1676037725
transform 1 0 264684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2877
timestamp 1676037725
transform 1 0 265788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2883
timestamp 1676037725
transform 1 0 266340 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2885
timestamp 1676037725
transform 1 0 266524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2897
timestamp 1676037725
transform 1 0 267628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2909
timestamp 1676037725
transform 1 0 268732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2921
timestamp 1676037725
transform 1 0 269836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2933
timestamp 1676037725
transform 1 0 270940 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2939
timestamp 1676037725
transform 1 0 271492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2941
timestamp 1676037725
transform 1 0 271676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2953
timestamp 1676037725
transform 1 0 272780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2965
timestamp 1676037725
transform 1 0 273884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2977
timestamp 1676037725
transform 1 0 274988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2989
timestamp 1676037725
transform 1 0 276092 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2995
timestamp 1676037725
transform 1 0 276644 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2997
timestamp 1676037725
transform 1 0 276828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3009
timestamp 1676037725
transform 1 0 277932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3021
timestamp 1676037725
transform 1 0 279036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3033
timestamp 1676037725
transform 1 0 280140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3045
timestamp 1676037725
transform 1 0 281244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3051
timestamp 1676037725
transform 1 0 281796 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3053
timestamp 1676037725
transform 1 0 281980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3065
timestamp 1676037725
transform 1 0 283084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3077
timestamp 1676037725
transform 1 0 284188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3089
timestamp 1676037725
transform 1 0 285292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3101
timestamp 1676037725
transform 1 0 286396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3107
timestamp 1676037725
transform 1 0 286948 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3109
timestamp 1676037725
transform 1 0 287132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3121
timestamp 1676037725
transform 1 0 288236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3133
timestamp 1676037725
transform 1 0 289340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3145
timestamp 1676037725
transform 1 0 290444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3157
timestamp 1676037725
transform 1 0 291548 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3163
timestamp 1676037725
transform 1 0 292100 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3165
timestamp 1676037725
transform 1 0 292284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3177
timestamp 1676037725
transform 1 0 293388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3189
timestamp 1676037725
transform 1 0 294492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3201
timestamp 1676037725
transform 1 0 295596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3213
timestamp 1676037725
transform 1 0 296700 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3219
timestamp 1676037725
transform 1 0 297252 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3221
timestamp 1676037725
transform 1 0 297436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3233
timestamp 1676037725
transform 1 0 298540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3245
timestamp 1676037725
transform 1 0 299644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3257
timestamp 1676037725
transform 1 0 300748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3269
timestamp 1676037725
transform 1 0 301852 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3275
timestamp 1676037725
transform 1 0 302404 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3277
timestamp 1676037725
transform 1 0 302588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3289
timestamp 1676037725
transform 1 0 303692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3301
timestamp 1676037725
transform 1 0 304796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3313
timestamp 1676037725
transform 1 0 305900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3325
timestamp 1676037725
transform 1 0 307004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3331
timestamp 1676037725
transform 1 0 307556 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3333
timestamp 1676037725
transform 1 0 307740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3345
timestamp 1676037725
transform 1 0 308844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3357
timestamp 1676037725
transform 1 0 309948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3369
timestamp 1676037725
transform 1 0 311052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3381
timestamp 1676037725
transform 1 0 312156 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3387
timestamp 1676037725
transform 1 0 312708 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3389
timestamp 1676037725
transform 1 0 312892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3401
timestamp 1676037725
transform 1 0 313996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3413
timestamp 1676037725
transform 1 0 315100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3425
timestamp 1676037725
transform 1 0 316204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3437
timestamp 1676037725
transform 1 0 317308 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3443
timestamp 1676037725
transform 1 0 317860 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3445
timestamp 1676037725
transform 1 0 318044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3457
timestamp 1676037725
transform 1 0 319148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3469
timestamp 1676037725
transform 1 0 320252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3481
timestamp 1676037725
transform 1 0 321356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3493
timestamp 1676037725
transform 1 0 322460 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3499
timestamp 1676037725
transform 1 0 323012 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3501
timestamp 1676037725
transform 1 0 323196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3513
timestamp 1676037725
transform 1 0 324300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3525
timestamp 1676037725
transform 1 0 325404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3537
timestamp 1676037725
transform 1 0 326508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3549
timestamp 1676037725
transform 1 0 327612 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3555
timestamp 1676037725
transform 1 0 328164 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3557
timestamp 1676037725
transform 1 0 328348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3569
timestamp 1676037725
transform 1 0 329452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3581
timestamp 1676037725
transform 1 0 330556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3593
timestamp 1676037725
transform 1 0 331660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3605
timestamp 1676037725
transform 1 0 332764 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3611
timestamp 1676037725
transform 1 0 333316 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3613
timestamp 1676037725
transform 1 0 333500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3625
timestamp 1676037725
transform 1 0 334604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3637
timestamp 1676037725
transform 1 0 335708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3649
timestamp 1676037725
transform 1 0 336812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3661
timestamp 1676037725
transform 1 0 337916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3667
timestamp 1676037725
transform 1 0 338468 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3669
timestamp 1676037725
transform 1 0 338652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3681
timestamp 1676037725
transform 1 0 339756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3693
timestamp 1676037725
transform 1 0 340860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3705
timestamp 1676037725
transform 1 0 341964 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3717
timestamp 1676037725
transform 1 0 343068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3723
timestamp 1676037725
transform 1 0 343620 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3725
timestamp 1676037725
transform 1 0 343804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3737
timestamp 1676037725
transform 1 0 344908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3749
timestamp 1676037725
transform 1 0 346012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3761
timestamp 1676037725
transform 1 0 347116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3773
timestamp 1676037725
transform 1 0 348220 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3779
timestamp 1676037725
transform 1 0 348772 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3781
timestamp 1676037725
transform 1 0 348956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3793
timestamp 1676037725
transform 1 0 350060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3805
timestamp 1676037725
transform 1 0 351164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3817
timestamp 1676037725
transform 1 0 352268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3829
timestamp 1676037725
transform 1 0 353372 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3835
timestamp 1676037725
transform 1 0 353924 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3837
timestamp 1676037725
transform 1 0 354108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3849
timestamp 1676037725
transform 1 0 355212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3861
timestamp 1676037725
transform 1 0 356316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3873
timestamp 1676037725
transform 1 0 357420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3885
timestamp 1676037725
transform 1 0 358524 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3891
timestamp 1676037725
transform 1 0 359076 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3893
timestamp 1676037725
transform 1 0 359260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3905
timestamp 1676037725
transform 1 0 360364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3917
timestamp 1676037725
transform 1 0 361468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3929
timestamp 1676037725
transform 1 0 362572 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3941
timestamp 1676037725
transform 1 0 363676 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3947
timestamp 1676037725
transform 1 0 364228 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3949
timestamp 1676037725
transform 1 0 364412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3961
timestamp 1676037725
transform 1 0 365516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3973
timestamp 1676037725
transform 1 0 366620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3985
timestamp 1676037725
transform 1 0 367724 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3997
timestamp 1676037725
transform 1 0 368828 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4003
timestamp 1676037725
transform 1 0 369380 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4005
timestamp 1676037725
transform 1 0 369564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4017
timestamp 1676037725
transform 1 0 370668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4029
timestamp 1676037725
transform 1 0 371772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4041
timestamp 1676037725
transform 1 0 372876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4053
timestamp 1676037725
transform 1 0 373980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4059
timestamp 1676037725
transform 1 0 374532 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4061
timestamp 1676037725
transform 1 0 374716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4073
timestamp 1676037725
transform 1 0 375820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4085
timestamp 1676037725
transform 1 0 376924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4097
timestamp 1676037725
transform 1 0 378028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4109
timestamp 1676037725
transform 1 0 379132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4115
timestamp 1676037725
transform 1 0 379684 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4117
timestamp 1676037725
transform 1 0 379868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4129
timestamp 1676037725
transform 1 0 380972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4141
timestamp 1676037725
transform 1 0 382076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4153
timestamp 1676037725
transform 1 0 383180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4165
timestamp 1676037725
transform 1 0 384284 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4171
timestamp 1676037725
transform 1 0 384836 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4173
timestamp 1676037725
transform 1 0 385020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4185
timestamp 1676037725
transform 1 0 386124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4197
timestamp 1676037725
transform 1 0 387228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4209
timestamp 1676037725
transform 1 0 388332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4221
timestamp 1676037725
transform 1 0 389436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4227
timestamp 1676037725
transform 1 0 389988 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4229
timestamp 1676037725
transform 1 0 390172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4241
timestamp 1676037725
transform 1 0 391276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4253
timestamp 1676037725
transform 1 0 392380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4265
timestamp 1676037725
transform 1 0 393484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4277
timestamp 1676037725
transform 1 0 394588 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4283
timestamp 1676037725
transform 1 0 395140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4285
timestamp 1676037725
transform 1 0 395324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4297
timestamp 1676037725
transform 1 0 396428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4309
timestamp 1676037725
transform 1 0 397532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4321
timestamp 1676037725
transform 1 0 398636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4333
timestamp 1676037725
transform 1 0 399740 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4339
timestamp 1676037725
transform 1 0 400292 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4341
timestamp 1676037725
transform 1 0 400476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4353
timestamp 1676037725
transform 1 0 401580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4365
timestamp 1676037725
transform 1 0 402684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4377
timestamp 1676037725
transform 1 0 403788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4389
timestamp 1676037725
transform 1 0 404892 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4395
timestamp 1676037725
transform 1 0 405444 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4397
timestamp 1676037725
transform 1 0 405628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4409
timestamp 1676037725
transform 1 0 406732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4421
timestamp 1676037725
transform 1 0 407836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4433
timestamp 1676037725
transform 1 0 408940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4445
timestamp 1676037725
transform 1 0 410044 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4451
timestamp 1676037725
transform 1 0 410596 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4453
timestamp 1676037725
transform 1 0 410780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4465
timestamp 1676037725
transform 1 0 411884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4477
timestamp 1676037725
transform 1 0 412988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4489
timestamp 1676037725
transform 1 0 414092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4501
timestamp 1676037725
transform 1 0 415196 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4507
timestamp 1676037725
transform 1 0 415748 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4509
timestamp 1676037725
transform 1 0 415932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4521
timestamp 1676037725
transform 1 0 417036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4533
timestamp 1676037725
transform 1 0 418140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4545
timestamp 1676037725
transform 1 0 419244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4557
timestamp 1676037725
transform 1 0 420348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4563
timestamp 1676037725
transform 1 0 420900 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4565
timestamp 1676037725
transform 1 0 421084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4577
timestamp 1676037725
transform 1 0 422188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4589
timestamp 1676037725
transform 1 0 423292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4601
timestamp 1676037725
transform 1 0 424396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4613
timestamp 1676037725
transform 1 0 425500 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4619
timestamp 1676037725
transform 1 0 426052 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4621
timestamp 1676037725
transform 1 0 426236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4633
timestamp 1676037725
transform 1 0 427340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4645
timestamp 1676037725
transform 1 0 428444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4657
timestamp 1676037725
transform 1 0 429548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4669
timestamp 1676037725
transform 1 0 430652 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4675
timestamp 1676037725
transform 1 0 431204 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4677
timestamp 1676037725
transform 1 0 431388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4689
timestamp 1676037725
transform 1 0 432492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4701
timestamp 1676037725
transform 1 0 433596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4713
timestamp 1676037725
transform 1 0 434700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4725
timestamp 1676037725
transform 1 0 435804 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4731
timestamp 1676037725
transform 1 0 436356 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4733
timestamp 1676037725
transform 1 0 436540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4745
timestamp 1676037725
transform 1 0 437644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4757
timestamp 1676037725
transform 1 0 438748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4769
timestamp 1676037725
transform 1 0 439852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4781
timestamp 1676037725
transform 1 0 440956 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4787
timestamp 1676037725
transform 1 0 441508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4789
timestamp 1676037725
transform 1 0 441692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4801
timestamp 1676037725
transform 1 0 442796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4813
timestamp 1676037725
transform 1 0 443900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4825
timestamp 1676037725
transform 1 0 445004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4837
timestamp 1676037725
transform 1 0 446108 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4843
timestamp 1676037725
transform 1 0 446660 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4845
timestamp 1676037725
transform 1 0 446844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4857
timestamp 1676037725
transform 1 0 447948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4869
timestamp 1676037725
transform 1 0 449052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4881
timestamp 1676037725
transform 1 0 450156 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4893
timestamp 1676037725
transform 1 0 451260 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4899
timestamp 1676037725
transform 1 0 451812 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4901
timestamp 1676037725
transform 1 0 451996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4913
timestamp 1676037725
transform 1 0 453100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4925
timestamp 1676037725
transform 1 0 454204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4937
timestamp 1676037725
transform 1 0 455308 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4949
timestamp 1676037725
transform 1 0 456412 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4955
timestamp 1676037725
transform 1 0 456964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4957
timestamp 1676037725
transform 1 0 457148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4969
timestamp 1676037725
transform 1 0 458252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4981
timestamp 1676037725
transform 1 0 459356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4993
timestamp 1676037725
transform 1 0 460460 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5005
timestamp 1676037725
transform 1 0 461564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5011
timestamp 1676037725
transform 1 0 462116 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5013
timestamp 1676037725
transform 1 0 462300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5025
timestamp 1676037725
transform 1 0 463404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5037
timestamp 1676037725
transform 1 0 464508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5049
timestamp 1676037725
transform 1 0 465612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5061
timestamp 1676037725
transform 1 0 466716 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5067
timestamp 1676037725
transform 1 0 467268 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5069
timestamp 1676037725
transform 1 0 467452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5081
timestamp 1676037725
transform 1 0 468556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5093
timestamp 1676037725
transform 1 0 469660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5105
timestamp 1676037725
transform 1 0 470764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5117
timestamp 1676037725
transform 1 0 471868 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5123
timestamp 1676037725
transform 1 0 472420 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5125
timestamp 1676037725
transform 1 0 472604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5137
timestamp 1676037725
transform 1 0 473708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5149
timestamp 1676037725
transform 1 0 474812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5161
timestamp 1676037725
transform 1 0 475916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5173
timestamp 1676037725
transform 1 0 477020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5179
timestamp 1676037725
transform 1 0 477572 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5181
timestamp 1676037725
transform 1 0 477756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5193
timestamp 1676037725
transform 1 0 478860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5205
timestamp 1676037725
transform 1 0 479964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5217
timestamp 1676037725
transform 1 0 481068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5229
timestamp 1676037725
transform 1 0 482172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5235
timestamp 1676037725
transform 1 0 482724 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5237
timestamp 1676037725
transform 1 0 482908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5249
timestamp 1676037725
transform 1 0 484012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5261
timestamp 1676037725
transform 1 0 485116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5273
timestamp 1676037725
transform 1 0 486220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5285
timestamp 1676037725
transform 1 0 487324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5291
timestamp 1676037725
transform 1 0 487876 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5293
timestamp 1676037725
transform 1 0 488060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5305
timestamp 1676037725
transform 1 0 489164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5317
timestamp 1676037725
transform 1 0 490268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5329
timestamp 1676037725
transform 1 0 491372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5341
timestamp 1676037725
transform 1 0 492476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5347
timestamp 1676037725
transform 1 0 493028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5349
timestamp 1676037725
transform 1 0 493212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5361
timestamp 1676037725
transform 1 0 494316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5373
timestamp 1676037725
transform 1 0 495420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5385
timestamp 1676037725
transform 1 0 496524 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5397
timestamp 1676037725
transform 1 0 497628 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5403
timestamp 1676037725
transform 1 0 498180 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5405
timestamp 1676037725
transform 1 0 498364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5417
timestamp 1676037725
transform 1 0 499468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5429
timestamp 1676037725
transform 1 0 500572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5441
timestamp 1676037725
transform 1 0 501676 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5453
timestamp 1676037725
transform 1 0 502780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5459
timestamp 1676037725
transform 1 0 503332 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5461
timestamp 1676037725
transform 1 0 503516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5473
timestamp 1676037725
transform 1 0 504620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5485
timestamp 1676037725
transform 1 0 505724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5497
timestamp 1676037725
transform 1 0 506828 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5509
timestamp 1676037725
transform 1 0 507932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5515
timestamp 1676037725
transform 1 0 508484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5517
timestamp 1676037725
transform 1 0 508668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5529
timestamp 1676037725
transform 1 0 509772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5541
timestamp 1676037725
transform 1 0 510876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5553
timestamp 1676037725
transform 1 0 511980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5565
timestamp 1676037725
transform 1 0 513084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5571
timestamp 1676037725
transform 1 0 513636 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5573
timestamp 1676037725
transform 1 0 513820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5585
timestamp 1676037725
transform 1 0 514924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5597
timestamp 1676037725
transform 1 0 516028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5609
timestamp 1676037725
transform 1 0 517132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5621
timestamp 1676037725
transform 1 0 518236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5627
timestamp 1676037725
transform 1 0 518788 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5629
timestamp 1676037725
transform 1 0 518972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5641
timestamp 1676037725
transform 1 0 520076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5653
timestamp 1676037725
transform 1 0 521180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5665
timestamp 1676037725
transform 1 0 522284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5677
timestamp 1676037725
transform 1 0 523388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5683
timestamp 1676037725
transform 1 0 523940 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5685
timestamp 1676037725
transform 1 0 524124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5697
timestamp 1676037725
transform 1 0 525228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5709
timestamp 1676037725
transform 1 0 526332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5721
timestamp 1676037725
transform 1 0 527436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5733
timestamp 1676037725
transform 1 0 528540 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5739
timestamp 1676037725
transform 1 0 529092 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5741
timestamp 1676037725
transform 1 0 529276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5753
timestamp 1676037725
transform 1 0 530380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5765
timestamp 1676037725
transform 1 0 531484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5777
timestamp 1676037725
transform 1 0 532588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5789
timestamp 1676037725
transform 1 0 533692 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5795
timestamp 1676037725
transform 1 0 534244 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5797
timestamp 1676037725
transform 1 0 534428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5809
timestamp 1676037725
transform 1 0 535532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5821
timestamp 1676037725
transform 1 0 536636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5833
timestamp 1676037725
transform 1 0 537740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5845
timestamp 1676037725
transform 1 0 538844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5851
timestamp 1676037725
transform 1 0 539396 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5853
timestamp 1676037725
transform 1 0 539580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5865
timestamp 1676037725
transform 1 0 540684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5877
timestamp 1676037725
transform 1 0 541788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5889
timestamp 1676037725
transform 1 0 542892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5901
timestamp 1676037725
transform 1 0 543996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5907
timestamp 1676037725
transform 1 0 544548 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5909
timestamp 1676037725
transform 1 0 544732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5921
timestamp 1676037725
transform 1 0 545836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5933
timestamp 1676037725
transform 1 0 546940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5945
timestamp 1676037725
transform 1 0 548044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5957
timestamp 1676037725
transform 1 0 549148 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5963
timestamp 1676037725
transform 1 0 549700 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5965
timestamp 1676037725
transform 1 0 549884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5977
timestamp 1676037725
transform 1 0 550988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5989
timestamp 1676037725
transform 1 0 552092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6001
timestamp 1676037725
transform 1 0 553196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6013
timestamp 1676037725
transform 1 0 554300 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6019
timestamp 1676037725
transform 1 0 554852 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6021
timestamp 1676037725
transform 1 0 555036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6033
timestamp 1676037725
transform 1 0 556140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6045
timestamp 1676037725
transform 1 0 557244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6057
timestamp 1676037725
transform 1 0 558348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6069
timestamp 1676037725
transform 1 0 559452 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6075
timestamp 1676037725
transform 1 0 560004 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6077
timestamp 1676037725
transform 1 0 560188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6089
timestamp 1676037725
transform 1 0 561292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6101
timestamp 1676037725
transform 1 0 562396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6113
timestamp 1676037725
transform 1 0 563500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6125
timestamp 1676037725
transform 1 0 564604 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6131
timestamp 1676037725
transform 1 0 565156 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6133
timestamp 1676037725
transform 1 0 565340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6145
timestamp 1676037725
transform 1 0 566444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6157
timestamp 1676037725
transform 1 0 567548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6169
timestamp 1676037725
transform 1 0 568652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6181
timestamp 1676037725
transform 1 0 569756 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6187
timestamp 1676037725
transform 1 0 570308 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6189
timestamp 1676037725
transform 1 0 570492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6201
timestamp 1676037725
transform 1 0 571596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6213
timestamp 1676037725
transform 1 0 572700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6225
timestamp 1676037725
transform 1 0 573804 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6237
timestamp 1676037725
transform 1 0 574908 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6243
timestamp 1676037725
transform 1 0 575460 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6245
timestamp 1676037725
transform 1 0 575644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6257
timestamp 1676037725
transform 1 0 576748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6269
timestamp 1676037725
transform 1 0 577852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6281
timestamp 1676037725
transform 1 0 578956 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6293
timestamp 1676037725
transform 1 0 580060 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6299
timestamp 1676037725
transform 1 0 580612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6301
timestamp 1676037725
transform 1 0 580796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6313
timestamp 1676037725
transform 1 0 581900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6325
timestamp 1676037725
transform 1 0 583004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6337
timestamp 1676037725
transform 1 0 584108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6349
timestamp 1676037725
transform 1 0 585212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6355
timestamp 1676037725
transform 1 0 585764 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6357
timestamp 1676037725
transform 1 0 585948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6369
timestamp 1676037725
transform 1 0 587052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6381
timestamp 1676037725
transform 1 0 588156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6393
timestamp 1676037725
transform 1 0 589260 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6405
timestamp 1676037725
transform 1 0 590364 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6411
timestamp 1676037725
transform 1 0 590916 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6413
timestamp 1676037725
transform 1 0 591100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6425
timestamp 1676037725
transform 1 0 592204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6437
timestamp 1676037725
transform 1 0 593308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6449
timestamp 1676037725
transform 1 0 594412 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6461
timestamp 1676037725
transform 1 0 595516 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6467
timestamp 1676037725
transform 1 0 596068 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6469
timestamp 1676037725
transform 1 0 596252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6481
timestamp 1676037725
transform 1 0 597356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6493
timestamp 1676037725
transform 1 0 598460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6505
timestamp 1676037725
transform 1 0 599564 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6517
timestamp 1676037725
transform 1 0 600668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6523
timestamp 1676037725
transform 1 0 601220 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6525
timestamp 1676037725
transform 1 0 601404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6537
timestamp 1676037725
transform 1 0 602508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6549
timestamp 1676037725
transform 1 0 603612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6561
timestamp 1676037725
transform 1 0 604716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6573
timestamp 1676037725
transform 1 0 605820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6579
timestamp 1676037725
transform 1 0 606372 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6581
timestamp 1676037725
transform 1 0 606556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6593
timestamp 1676037725
transform 1 0 607660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6605
timestamp 1676037725
transform 1 0 608764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6617
timestamp 1676037725
transform 1 0 609868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6629
timestamp 1676037725
transform 1 0 610972 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6635
timestamp 1676037725
transform 1 0 611524 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6637
timestamp 1676037725
transform 1 0 611708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6649
timestamp 1676037725
transform 1 0 612812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6661
timestamp 1676037725
transform 1 0 613916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6673
timestamp 1676037725
transform 1 0 615020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6685
timestamp 1676037725
transform 1 0 616124 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6691
timestamp 1676037725
transform 1 0 616676 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6693
timestamp 1676037725
transform 1 0 616860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6705
timestamp 1676037725
transform 1 0 617964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6717
timestamp 1676037725
transform 1 0 619068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6729
timestamp 1676037725
transform 1 0 620172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6741
timestamp 1676037725
transform 1 0 621276 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6747
timestamp 1676037725
transform 1 0 621828 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6749
timestamp 1676037725
transform 1 0 622012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6761
timestamp 1676037725
transform 1 0 623116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6773
timestamp 1676037725
transform 1 0 624220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6785
timestamp 1676037725
transform 1 0 625324 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6797
timestamp 1676037725
transform 1 0 626428 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6803
timestamp 1676037725
transform 1 0 626980 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6805
timestamp 1676037725
transform 1 0 627164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6817
timestamp 1676037725
transform 1 0 628268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6829
timestamp 1676037725
transform 1 0 629372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6841
timestamp 1676037725
transform 1 0 630476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6853
timestamp 1676037725
transform 1 0 631580 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6859
timestamp 1676037725
transform 1 0 632132 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6861
timestamp 1676037725
transform 1 0 632316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6873
timestamp 1676037725
transform 1 0 633420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6885
timestamp 1676037725
transform 1 0 634524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6897
timestamp 1676037725
transform 1 0 635628 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6909
timestamp 1676037725
transform 1 0 636732 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6915
timestamp 1676037725
transform 1 0 637284 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6917
timestamp 1676037725
transform 1 0 637468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6929
timestamp 1676037725
transform 1 0 638572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6941
timestamp 1676037725
transform 1 0 639676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6953
timestamp 1676037725
transform 1 0 640780 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_6965
timestamp 1676037725
transform 1 0 641884 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6971
timestamp 1676037725
transform 1 0 642436 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6973
timestamp 1676037725
transform 1 0 642620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6985
timestamp 1676037725
transform 1 0 643724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6997
timestamp 1676037725
transform 1 0 644828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7009
timestamp 1676037725
transform 1 0 645932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7021
timestamp 1676037725
transform 1 0 647036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7027
timestamp 1676037725
transform 1 0 647588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7029
timestamp 1676037725
transform 1 0 647772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7041
timestamp 1676037725
transform 1 0 648876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7053
timestamp 1676037725
transform 1 0 649980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7065
timestamp 1676037725
transform 1 0 651084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7077
timestamp 1676037725
transform 1 0 652188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7083
timestamp 1676037725
transform 1 0 652740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7085
timestamp 1676037725
transform 1 0 652924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7097
timestamp 1676037725
transform 1 0 654028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7109
timestamp 1676037725
transform 1 0 655132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7121
timestamp 1676037725
transform 1 0 656236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7133
timestamp 1676037725
transform 1 0 657340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7139
timestamp 1676037725
transform 1 0 657892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7141
timestamp 1676037725
transform 1 0 658076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7153
timestamp 1676037725
transform 1 0 659180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7165
timestamp 1676037725
transform 1 0 660284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7177
timestamp 1676037725
transform 1 0 661388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7189
timestamp 1676037725
transform 1 0 662492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7195
timestamp 1676037725
transform 1 0 663044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7197
timestamp 1676037725
transform 1 0 663228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7209
timestamp 1676037725
transform 1 0 664332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7221
timestamp 1676037725
transform 1 0 665436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7233
timestamp 1676037725
transform 1 0 666540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7245
timestamp 1676037725
transform 1 0 667644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7251
timestamp 1676037725
transform 1 0 668196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7253
timestamp 1676037725
transform 1 0 668380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7265
timestamp 1676037725
transform 1 0 669484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7277
timestamp 1676037725
transform 1 0 670588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7289
timestamp 1676037725
transform 1 0 671692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7301
timestamp 1676037725
transform 1 0 672796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7307
timestamp 1676037725
transform 1 0 673348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7309
timestamp 1676037725
transform 1 0 673532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7321
timestamp 1676037725
transform 1 0 674636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7333
timestamp 1676037725
transform 1 0 675740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7345
timestamp 1676037725
transform 1 0 676844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7357
timestamp 1676037725
transform 1 0 677948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7363
timestamp 1676037725
transform 1 0 678500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7365
timestamp 1676037725
transform 1 0 678684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7377
timestamp 1676037725
transform 1 0 679788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7389
timestamp 1676037725
transform 1 0 680892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7401
timestamp 1676037725
transform 1 0 681996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1676037725
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1676037725
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_85
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1676037725
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1676037725
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_141
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_153
timestamp 1676037725
transform 1 0 15180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1676037725
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1676037725
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1676037725
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1676037725
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1676037725
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1676037725
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_309
timestamp 1676037725
transform 1 0 29532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1676037725
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1676037725
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_365
timestamp 1676037725
transform 1 0 34684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_377
timestamp 1676037725
transform 1 0 35788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1676037725
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_421
timestamp 1676037725
transform 1 0 39836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_433
timestamp 1676037725
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1676037725
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_477
timestamp 1676037725
transform 1 0 44988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_489
timestamp 1676037725
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1676037725
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_533
timestamp 1676037725
transform 1 0 50140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_545
timestamp 1676037725
transform 1 0 51244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_557
timestamp 1676037725
transform 1 0 52348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_589
timestamp 1676037725
transform 1 0 55292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_601
timestamp 1676037725
transform 1 0 56396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_613
timestamp 1676037725
transform 1 0 57500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1676037725
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_641
timestamp 1676037725
transform 1 0 60076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_645
timestamp 1676037725
transform 1 0 60444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_657
timestamp 1676037725
transform 1 0 61548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_669
timestamp 1676037725
transform 1 0 62652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1676037725
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1676037725
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_697
timestamp 1676037725
transform 1 0 65228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_701
timestamp 1676037725
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_713
timestamp 1676037725
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_725
timestamp 1676037725
transform 1 0 67804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1676037725
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1676037725
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_753
timestamp 1676037725
transform 1 0 70380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_757
timestamp 1676037725
transform 1 0 70748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_769
timestamp 1676037725
transform 1 0 71852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_781
timestamp 1676037725
transform 1 0 72956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1676037725
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1676037725
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_809
timestamp 1676037725
transform 1 0 75532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_813
timestamp 1676037725
transform 1 0 75900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_825
timestamp 1676037725
transform 1 0 77004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_837
timestamp 1676037725
transform 1 0 78108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1676037725
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1676037725
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_865
timestamp 1676037725
transform 1 0 80684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_869
timestamp 1676037725
transform 1 0 81052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_881
timestamp 1676037725
transform 1 0 82156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_893
timestamp 1676037725
transform 1 0 83260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1676037725
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1676037725
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_921
timestamp 1676037725
transform 1 0 85836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_925
timestamp 1676037725
transform 1 0 86204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_937
timestamp 1676037725
transform 1 0 87308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_949
timestamp 1676037725
transform 1 0 88412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1676037725
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1676037725
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_977
timestamp 1676037725
transform 1 0 90988 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_981
timestamp 1676037725
transform 1 0 91356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_993
timestamp 1676037725
transform 1 0 92460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1005
timestamp 1676037725
transform 1 0 93564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1676037725
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1676037725
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1033
timestamp 1676037725
transform 1 0 96140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1037
timestamp 1676037725
transform 1 0 96508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1049
timestamp 1676037725
transform 1 0 97612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1061
timestamp 1676037725
transform 1 0 98716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1676037725
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1676037725
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1089
timestamp 1676037725
transform 1 0 101292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1093
timestamp 1676037725
transform 1 0 101660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1105
timestamp 1676037725
transform 1 0 102764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1117
timestamp 1676037725
transform 1 0 103868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1676037725
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1676037725
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1145
timestamp 1676037725
transform 1 0 106444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1149
timestamp 1676037725
transform 1 0 106812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1161
timestamp 1676037725
transform 1 0 107916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1173
timestamp 1676037725
transform 1 0 109020 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1676037725
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1189
timestamp 1676037725
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1201
timestamp 1676037725
transform 1 0 111596 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1205
timestamp 1676037725
transform 1 0 111964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1217
timestamp 1676037725
transform 1 0 113068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1229
timestamp 1676037725
transform 1 0 114172 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1676037725
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1676037725
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1257
timestamp 1676037725
transform 1 0 116748 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1261
timestamp 1676037725
transform 1 0 117116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1273
timestamp 1676037725
transform 1 0 118220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1285
timestamp 1676037725
transform 1 0 119324 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1289
timestamp 1676037725
transform 1 0 119692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1301
timestamp 1676037725
transform 1 0 120796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1313
timestamp 1676037725
transform 1 0 121900 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1317
timestamp 1676037725
transform 1 0 122268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1329
timestamp 1676037725
transform 1 0 123372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1341
timestamp 1676037725
transform 1 0 124476 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1345
timestamp 1676037725
transform 1 0 124844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1357
timestamp 1676037725
transform 1 0 125948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1369
timestamp 1676037725
transform 1 0 127052 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1373
timestamp 1676037725
transform 1 0 127420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1385
timestamp 1676037725
transform 1 0 128524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1397
timestamp 1676037725
transform 1 0 129628 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1401
timestamp 1676037725
transform 1 0 129996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1413
timestamp 1676037725
transform 1 0 131100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1425
timestamp 1676037725
transform 1 0 132204 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1429
timestamp 1676037725
transform 1 0 132572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1441
timestamp 1676037725
transform 1 0 133676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1453
timestamp 1676037725
transform 1 0 134780 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1457
timestamp 1676037725
transform 1 0 135148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1469
timestamp 1676037725
transform 1 0 136252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1481
timestamp 1676037725
transform 1 0 137356 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1485
timestamp 1676037725
transform 1 0 137724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1497
timestamp 1676037725
transform 1 0 138828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1509
timestamp 1676037725
transform 1 0 139932 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1513
timestamp 1676037725
transform 1 0 140300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1525
timestamp 1676037725
transform 1 0 141404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1537
timestamp 1676037725
transform 1 0 142508 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1541
timestamp 1676037725
transform 1 0 142876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1553
timestamp 1676037725
transform 1 0 143980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1565
timestamp 1676037725
transform 1 0 145084 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1569
timestamp 1676037725
transform 1 0 145452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1581
timestamp 1676037725
transform 1 0 146556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1593
timestamp 1676037725
transform 1 0 147660 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1597
timestamp 1676037725
transform 1 0 148028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1609
timestamp 1676037725
transform 1 0 149132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1621
timestamp 1676037725
transform 1 0 150236 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1625
timestamp 1676037725
transform 1 0 150604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1637
timestamp 1676037725
transform 1 0 151708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1649
timestamp 1676037725
transform 1 0 152812 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1653
timestamp 1676037725
transform 1 0 153180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1665
timestamp 1676037725
transform 1 0 154284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1677
timestamp 1676037725
transform 1 0 155388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1681
timestamp 1676037725
transform 1 0 155756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1693
timestamp 1676037725
transform 1 0 156860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1705
timestamp 1676037725
transform 1 0 157964 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1709
timestamp 1676037725
transform 1 0 158332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1721
timestamp 1676037725
transform 1 0 159436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1733
timestamp 1676037725
transform 1 0 160540 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1737
timestamp 1676037725
transform 1 0 160908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1749
timestamp 1676037725
transform 1 0 162012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1761
timestamp 1676037725
transform 1 0 163116 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1765
timestamp 1676037725
transform 1 0 163484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1777
timestamp 1676037725
transform 1 0 164588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1789
timestamp 1676037725
transform 1 0 165692 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1793
timestamp 1676037725
transform 1 0 166060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1805
timestamp 1676037725
transform 1 0 167164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1817
timestamp 1676037725
transform 1 0 168268 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1821
timestamp 1676037725
transform 1 0 168636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1833
timestamp 1676037725
transform 1 0 169740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1845
timestamp 1676037725
transform 1 0 170844 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1849
timestamp 1676037725
transform 1 0 171212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1861
timestamp 1676037725
transform 1 0 172316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1873
timestamp 1676037725
transform 1 0 173420 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1877
timestamp 1676037725
transform 1 0 173788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1889
timestamp 1676037725
transform 1 0 174892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1901
timestamp 1676037725
transform 1 0 175996 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1905
timestamp 1676037725
transform 1 0 176364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1917
timestamp 1676037725
transform 1 0 177468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1929
timestamp 1676037725
transform 1 0 178572 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1933
timestamp 1676037725
transform 1 0 178940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1945
timestamp 1676037725
transform 1 0 180044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1957
timestamp 1676037725
transform 1 0 181148 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1961
timestamp 1676037725
transform 1 0 181516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1973
timestamp 1676037725
transform 1 0 182620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1985
timestamp 1676037725
transform 1 0 183724 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1989
timestamp 1676037725
transform 1 0 184092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2001
timestamp 1676037725
transform 1 0 185196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2013
timestamp 1676037725
transform 1 0 186300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2017
timestamp 1676037725
transform 1 0 186668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2029
timestamp 1676037725
transform 1 0 187772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2041
timestamp 1676037725
transform 1 0 188876 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2045
timestamp 1676037725
transform 1 0 189244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2057
timestamp 1676037725
transform 1 0 190348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2069
timestamp 1676037725
transform 1 0 191452 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2073
timestamp 1676037725
transform 1 0 191820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2085
timestamp 1676037725
transform 1 0 192924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2097
timestamp 1676037725
transform 1 0 194028 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2101
timestamp 1676037725
transform 1 0 194396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2113
timestamp 1676037725
transform 1 0 195500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2125
timestamp 1676037725
transform 1 0 196604 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2129
timestamp 1676037725
transform 1 0 196972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2141
timestamp 1676037725
transform 1 0 198076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2153
timestamp 1676037725
transform 1 0 199180 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2157
timestamp 1676037725
transform 1 0 199548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2169
timestamp 1676037725
transform 1 0 200652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2181
timestamp 1676037725
transform 1 0 201756 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2185
timestamp 1676037725
transform 1 0 202124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2197
timestamp 1676037725
transform 1 0 203228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2209
timestamp 1676037725
transform 1 0 204332 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2213
timestamp 1676037725
transform 1 0 204700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2225
timestamp 1676037725
transform 1 0 205804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2237
timestamp 1676037725
transform 1 0 206908 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2241
timestamp 1676037725
transform 1 0 207276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2253
timestamp 1676037725
transform 1 0 208380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2265
timestamp 1676037725
transform 1 0 209484 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2269
timestamp 1676037725
transform 1 0 209852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2281
timestamp 1676037725
transform 1 0 210956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2293
timestamp 1676037725
transform 1 0 212060 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2297
timestamp 1676037725
transform 1 0 212428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2309
timestamp 1676037725
transform 1 0 213532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2321
timestamp 1676037725
transform 1 0 214636 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2325
timestamp 1676037725
transform 1 0 215004 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2337
timestamp 1676037725
transform 1 0 216108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2349
timestamp 1676037725
transform 1 0 217212 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2353
timestamp 1676037725
transform 1 0 217580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2365
timestamp 1676037725
transform 1 0 218684 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2377
timestamp 1676037725
transform 1 0 219788 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2381
timestamp 1676037725
transform 1 0 220156 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2393
timestamp 1676037725
transform 1 0 221260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2405
timestamp 1676037725
transform 1 0 222364 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2409
timestamp 1676037725
transform 1 0 222732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2421
timestamp 1676037725
transform 1 0 223836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2433
timestamp 1676037725
transform 1 0 224940 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2437
timestamp 1676037725
transform 1 0 225308 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2449
timestamp 1676037725
transform 1 0 226412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2461
timestamp 1676037725
transform 1 0 227516 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2465
timestamp 1676037725
transform 1 0 227884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2477
timestamp 1676037725
transform 1 0 228988 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2489
timestamp 1676037725
transform 1 0 230092 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2493
timestamp 1676037725
transform 1 0 230460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2505
timestamp 1676037725
transform 1 0 231564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2517
timestamp 1676037725
transform 1 0 232668 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2521
timestamp 1676037725
transform 1 0 233036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2533
timestamp 1676037725
transform 1 0 234140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2545
timestamp 1676037725
transform 1 0 235244 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2549
timestamp 1676037725
transform 1 0 235612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2561
timestamp 1676037725
transform 1 0 236716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2573
timestamp 1676037725
transform 1 0 237820 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2577
timestamp 1676037725
transform 1 0 238188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2589
timestamp 1676037725
transform 1 0 239292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2601
timestamp 1676037725
transform 1 0 240396 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2605
timestamp 1676037725
transform 1 0 240764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2617
timestamp 1676037725
transform 1 0 241868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2629
timestamp 1676037725
transform 1 0 242972 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2633
timestamp 1676037725
transform 1 0 243340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2645
timestamp 1676037725
transform 1 0 244444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2657
timestamp 1676037725
transform 1 0 245548 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2661
timestamp 1676037725
transform 1 0 245916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2673
timestamp 1676037725
transform 1 0 247020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2685
timestamp 1676037725
transform 1 0 248124 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2689
timestamp 1676037725
transform 1 0 248492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2701
timestamp 1676037725
transform 1 0 249596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2713
timestamp 1676037725
transform 1 0 250700 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2717
timestamp 1676037725
transform 1 0 251068 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2729
timestamp 1676037725
transform 1 0 252172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2741
timestamp 1676037725
transform 1 0 253276 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2745
timestamp 1676037725
transform 1 0 253644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2757
timestamp 1676037725
transform 1 0 254748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2769
timestamp 1676037725
transform 1 0 255852 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2773
timestamp 1676037725
transform 1 0 256220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2785
timestamp 1676037725
transform 1 0 257324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2797
timestamp 1676037725
transform 1 0 258428 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2801
timestamp 1676037725
transform 1 0 258796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2813
timestamp 1676037725
transform 1 0 259900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2825
timestamp 1676037725
transform 1 0 261004 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2829
timestamp 1676037725
transform 1 0 261372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2841
timestamp 1676037725
transform 1 0 262476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2853
timestamp 1676037725
transform 1 0 263580 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2857
timestamp 1676037725
transform 1 0 263948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2869
timestamp 1676037725
transform 1 0 265052 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2881
timestamp 1676037725
transform 1 0 266156 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2885
timestamp 1676037725
transform 1 0 266524 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2897
timestamp 1676037725
transform 1 0 267628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2909
timestamp 1676037725
transform 1 0 268732 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2913
timestamp 1676037725
transform 1 0 269100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2925
timestamp 1676037725
transform 1 0 270204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2937
timestamp 1676037725
transform 1 0 271308 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2941
timestamp 1676037725
transform 1 0 271676 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2953
timestamp 1676037725
transform 1 0 272780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2965
timestamp 1676037725
transform 1 0 273884 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2969
timestamp 1676037725
transform 1 0 274252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2981
timestamp 1676037725
transform 1 0 275356 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_2993
timestamp 1676037725
transform 1 0 276460 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2997
timestamp 1676037725
transform 1 0 276828 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3009
timestamp 1676037725
transform 1 0 277932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3021
timestamp 1676037725
transform 1 0 279036 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3025
timestamp 1676037725
transform 1 0 279404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3037
timestamp 1676037725
transform 1 0 280508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3049
timestamp 1676037725
transform 1 0 281612 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3053
timestamp 1676037725
transform 1 0 281980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3065
timestamp 1676037725
transform 1 0 283084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3077
timestamp 1676037725
transform 1 0 284188 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3081
timestamp 1676037725
transform 1 0 284556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3093
timestamp 1676037725
transform 1 0 285660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3105
timestamp 1676037725
transform 1 0 286764 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3109
timestamp 1676037725
transform 1 0 287132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3121
timestamp 1676037725
transform 1 0 288236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3133
timestamp 1676037725
transform 1 0 289340 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3137
timestamp 1676037725
transform 1 0 289708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3149
timestamp 1676037725
transform 1 0 290812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3161
timestamp 1676037725
transform 1 0 291916 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3165
timestamp 1676037725
transform 1 0 292284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3177
timestamp 1676037725
transform 1 0 293388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3189
timestamp 1676037725
transform 1 0 294492 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3193
timestamp 1676037725
transform 1 0 294860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3205
timestamp 1676037725
transform 1 0 295964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3217
timestamp 1676037725
transform 1 0 297068 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3221
timestamp 1676037725
transform 1 0 297436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3233
timestamp 1676037725
transform 1 0 298540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3245
timestamp 1676037725
transform 1 0 299644 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3249
timestamp 1676037725
transform 1 0 300012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3261
timestamp 1676037725
transform 1 0 301116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3273
timestamp 1676037725
transform 1 0 302220 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3277
timestamp 1676037725
transform 1 0 302588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3289
timestamp 1676037725
transform 1 0 303692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3301
timestamp 1676037725
transform 1 0 304796 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3305
timestamp 1676037725
transform 1 0 305164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3317
timestamp 1676037725
transform 1 0 306268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3329
timestamp 1676037725
transform 1 0 307372 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3333
timestamp 1676037725
transform 1 0 307740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3345
timestamp 1676037725
transform 1 0 308844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3357
timestamp 1676037725
transform 1 0 309948 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3361
timestamp 1676037725
transform 1 0 310316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3373
timestamp 1676037725
transform 1 0 311420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3385
timestamp 1676037725
transform 1 0 312524 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3389
timestamp 1676037725
transform 1 0 312892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3401
timestamp 1676037725
transform 1 0 313996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3413
timestamp 1676037725
transform 1 0 315100 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3417
timestamp 1676037725
transform 1 0 315468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3429
timestamp 1676037725
transform 1 0 316572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3441
timestamp 1676037725
transform 1 0 317676 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3445
timestamp 1676037725
transform 1 0 318044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3457
timestamp 1676037725
transform 1 0 319148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3469
timestamp 1676037725
transform 1 0 320252 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3473
timestamp 1676037725
transform 1 0 320620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3485
timestamp 1676037725
transform 1 0 321724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3497
timestamp 1676037725
transform 1 0 322828 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3501
timestamp 1676037725
transform 1 0 323196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3513
timestamp 1676037725
transform 1 0 324300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3525
timestamp 1676037725
transform 1 0 325404 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3529
timestamp 1676037725
transform 1 0 325772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3541
timestamp 1676037725
transform 1 0 326876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3553
timestamp 1676037725
transform 1 0 327980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3557
timestamp 1676037725
transform 1 0 328348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3569
timestamp 1676037725
transform 1 0 329452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3581
timestamp 1676037725
transform 1 0 330556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3585
timestamp 1676037725
transform 1 0 330924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3597
timestamp 1676037725
transform 1 0 332028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3609
timestamp 1676037725
transform 1 0 333132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3613
timestamp 1676037725
transform 1 0 333500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3625
timestamp 1676037725
transform 1 0 334604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3637
timestamp 1676037725
transform 1 0 335708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3641
timestamp 1676037725
transform 1 0 336076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3653
timestamp 1676037725
transform 1 0 337180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3665
timestamp 1676037725
transform 1 0 338284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3669
timestamp 1676037725
transform 1 0 338652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3681
timestamp 1676037725
transform 1 0 339756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3693
timestamp 1676037725
transform 1 0 340860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3697
timestamp 1676037725
transform 1 0 341228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3709
timestamp 1676037725
transform 1 0 342332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3721
timestamp 1676037725
transform 1 0 343436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3725
timestamp 1676037725
transform 1 0 343804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3737
timestamp 1676037725
transform 1 0 344908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3749
timestamp 1676037725
transform 1 0 346012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3753
timestamp 1676037725
transform 1 0 346380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3765
timestamp 1676037725
transform 1 0 347484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3777
timestamp 1676037725
transform 1 0 348588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3781
timestamp 1676037725
transform 1 0 348956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3793
timestamp 1676037725
transform 1 0 350060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3805
timestamp 1676037725
transform 1 0 351164 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3809
timestamp 1676037725
transform 1 0 351532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3821
timestamp 1676037725
transform 1 0 352636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3833
timestamp 1676037725
transform 1 0 353740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3837
timestamp 1676037725
transform 1 0 354108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3849
timestamp 1676037725
transform 1 0 355212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3861
timestamp 1676037725
transform 1 0 356316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3865
timestamp 1676037725
transform 1 0 356684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3877
timestamp 1676037725
transform 1 0 357788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3889
timestamp 1676037725
transform 1 0 358892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3893
timestamp 1676037725
transform 1 0 359260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3905
timestamp 1676037725
transform 1 0 360364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3917
timestamp 1676037725
transform 1 0 361468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3921
timestamp 1676037725
transform 1 0 361836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3933
timestamp 1676037725
transform 1 0 362940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3945
timestamp 1676037725
transform 1 0 364044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3949
timestamp 1676037725
transform 1 0 364412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3961
timestamp 1676037725
transform 1 0 365516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3973
timestamp 1676037725
transform 1 0 366620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3977
timestamp 1676037725
transform 1 0 366988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3989
timestamp 1676037725
transform 1 0 368092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4001
timestamp 1676037725
transform 1 0 369196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4005
timestamp 1676037725
transform 1 0 369564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4017
timestamp 1676037725
transform 1 0 370668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4029
timestamp 1676037725
transform 1 0 371772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4033
timestamp 1676037725
transform 1 0 372140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4045
timestamp 1676037725
transform 1 0 373244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4057
timestamp 1676037725
transform 1 0 374348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4061
timestamp 1676037725
transform 1 0 374716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4073
timestamp 1676037725
transform 1 0 375820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4085
timestamp 1676037725
transform 1 0 376924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4089
timestamp 1676037725
transform 1 0 377292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4101
timestamp 1676037725
transform 1 0 378396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4113
timestamp 1676037725
transform 1 0 379500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4117
timestamp 1676037725
transform 1 0 379868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4129
timestamp 1676037725
transform 1 0 380972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4141
timestamp 1676037725
transform 1 0 382076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4145
timestamp 1676037725
transform 1 0 382444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4157
timestamp 1676037725
transform 1 0 383548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4169
timestamp 1676037725
transform 1 0 384652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4173
timestamp 1676037725
transform 1 0 385020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4185
timestamp 1676037725
transform 1 0 386124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4197
timestamp 1676037725
transform 1 0 387228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4201
timestamp 1676037725
transform 1 0 387596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4213
timestamp 1676037725
transform 1 0 388700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4225
timestamp 1676037725
transform 1 0 389804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4229
timestamp 1676037725
transform 1 0 390172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4241
timestamp 1676037725
transform 1 0 391276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4253
timestamp 1676037725
transform 1 0 392380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4257
timestamp 1676037725
transform 1 0 392748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4269
timestamp 1676037725
transform 1 0 393852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4281
timestamp 1676037725
transform 1 0 394956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4285
timestamp 1676037725
transform 1 0 395324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4297
timestamp 1676037725
transform 1 0 396428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4309
timestamp 1676037725
transform 1 0 397532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4313
timestamp 1676037725
transform 1 0 397900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4325
timestamp 1676037725
transform 1 0 399004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4337
timestamp 1676037725
transform 1 0 400108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4341
timestamp 1676037725
transform 1 0 400476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4353
timestamp 1676037725
transform 1 0 401580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4365
timestamp 1676037725
transform 1 0 402684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4369
timestamp 1676037725
transform 1 0 403052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4381
timestamp 1676037725
transform 1 0 404156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4393
timestamp 1676037725
transform 1 0 405260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4397
timestamp 1676037725
transform 1 0 405628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4409
timestamp 1676037725
transform 1 0 406732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4421
timestamp 1676037725
transform 1 0 407836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4425
timestamp 1676037725
transform 1 0 408204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4437
timestamp 1676037725
transform 1 0 409308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4449
timestamp 1676037725
transform 1 0 410412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4453
timestamp 1676037725
transform 1 0 410780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4465
timestamp 1676037725
transform 1 0 411884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4477
timestamp 1676037725
transform 1 0 412988 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4481
timestamp 1676037725
transform 1 0 413356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4493
timestamp 1676037725
transform 1 0 414460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4505
timestamp 1676037725
transform 1 0 415564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4509
timestamp 1676037725
transform 1 0 415932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4521
timestamp 1676037725
transform 1 0 417036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4533
timestamp 1676037725
transform 1 0 418140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4537
timestamp 1676037725
transform 1 0 418508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4549
timestamp 1676037725
transform 1 0 419612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4561
timestamp 1676037725
transform 1 0 420716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4565
timestamp 1676037725
transform 1 0 421084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4577
timestamp 1676037725
transform 1 0 422188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4589
timestamp 1676037725
transform 1 0 423292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4593
timestamp 1676037725
transform 1 0 423660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4605
timestamp 1676037725
transform 1 0 424764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4617
timestamp 1676037725
transform 1 0 425868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4621
timestamp 1676037725
transform 1 0 426236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4633
timestamp 1676037725
transform 1 0 427340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4645
timestamp 1676037725
transform 1 0 428444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4649
timestamp 1676037725
transform 1 0 428812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4661
timestamp 1676037725
transform 1 0 429916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4673
timestamp 1676037725
transform 1 0 431020 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4677
timestamp 1676037725
transform 1 0 431388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4689
timestamp 1676037725
transform 1 0 432492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4701
timestamp 1676037725
transform 1 0 433596 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4705
timestamp 1676037725
transform 1 0 433964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4717
timestamp 1676037725
transform 1 0 435068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4729
timestamp 1676037725
transform 1 0 436172 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4733
timestamp 1676037725
transform 1 0 436540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4745
timestamp 1676037725
transform 1 0 437644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4757
timestamp 1676037725
transform 1 0 438748 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4761
timestamp 1676037725
transform 1 0 439116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4773
timestamp 1676037725
transform 1 0 440220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4785
timestamp 1676037725
transform 1 0 441324 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4789
timestamp 1676037725
transform 1 0 441692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4801
timestamp 1676037725
transform 1 0 442796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4813
timestamp 1676037725
transform 1 0 443900 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4817
timestamp 1676037725
transform 1 0 444268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4829
timestamp 1676037725
transform 1 0 445372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4841
timestamp 1676037725
transform 1 0 446476 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4845
timestamp 1676037725
transform 1 0 446844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4857
timestamp 1676037725
transform 1 0 447948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4869
timestamp 1676037725
transform 1 0 449052 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4873
timestamp 1676037725
transform 1 0 449420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4885
timestamp 1676037725
transform 1 0 450524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4897
timestamp 1676037725
transform 1 0 451628 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4901
timestamp 1676037725
transform 1 0 451996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4913
timestamp 1676037725
transform 1 0 453100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4925
timestamp 1676037725
transform 1 0 454204 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4929
timestamp 1676037725
transform 1 0 454572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4941
timestamp 1676037725
transform 1 0 455676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4953
timestamp 1676037725
transform 1 0 456780 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4957
timestamp 1676037725
transform 1 0 457148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4969
timestamp 1676037725
transform 1 0 458252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_4981
timestamp 1676037725
transform 1 0 459356 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4985
timestamp 1676037725
transform 1 0 459724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4997
timestamp 1676037725
transform 1 0 460828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5009
timestamp 1676037725
transform 1 0 461932 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5013
timestamp 1676037725
transform 1 0 462300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5025
timestamp 1676037725
transform 1 0 463404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5037
timestamp 1676037725
transform 1 0 464508 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5041
timestamp 1676037725
transform 1 0 464876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5053
timestamp 1676037725
transform 1 0 465980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5065
timestamp 1676037725
transform 1 0 467084 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5069
timestamp 1676037725
transform 1 0 467452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5081
timestamp 1676037725
transform 1 0 468556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5093
timestamp 1676037725
transform 1 0 469660 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5097
timestamp 1676037725
transform 1 0 470028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5109
timestamp 1676037725
transform 1 0 471132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5121
timestamp 1676037725
transform 1 0 472236 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5125
timestamp 1676037725
transform 1 0 472604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5137
timestamp 1676037725
transform 1 0 473708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5149
timestamp 1676037725
transform 1 0 474812 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5153
timestamp 1676037725
transform 1 0 475180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5165
timestamp 1676037725
transform 1 0 476284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5177
timestamp 1676037725
transform 1 0 477388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5181
timestamp 1676037725
transform 1 0 477756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5193
timestamp 1676037725
transform 1 0 478860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5205
timestamp 1676037725
transform 1 0 479964 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5209
timestamp 1676037725
transform 1 0 480332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5221
timestamp 1676037725
transform 1 0 481436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5233
timestamp 1676037725
transform 1 0 482540 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5237
timestamp 1676037725
transform 1 0 482908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5249
timestamp 1676037725
transform 1 0 484012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5261
timestamp 1676037725
transform 1 0 485116 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5265
timestamp 1676037725
transform 1 0 485484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5277
timestamp 1676037725
transform 1 0 486588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5289
timestamp 1676037725
transform 1 0 487692 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5293
timestamp 1676037725
transform 1 0 488060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5305
timestamp 1676037725
transform 1 0 489164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5317
timestamp 1676037725
transform 1 0 490268 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5321
timestamp 1676037725
transform 1 0 490636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5333
timestamp 1676037725
transform 1 0 491740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5345
timestamp 1676037725
transform 1 0 492844 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5349
timestamp 1676037725
transform 1 0 493212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5361
timestamp 1676037725
transform 1 0 494316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5373
timestamp 1676037725
transform 1 0 495420 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5377
timestamp 1676037725
transform 1 0 495788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5389
timestamp 1676037725
transform 1 0 496892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5401
timestamp 1676037725
transform 1 0 497996 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5405
timestamp 1676037725
transform 1 0 498364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5417
timestamp 1676037725
transform 1 0 499468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5429
timestamp 1676037725
transform 1 0 500572 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5433
timestamp 1676037725
transform 1 0 500940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5445
timestamp 1676037725
transform 1 0 502044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5457
timestamp 1676037725
transform 1 0 503148 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5461
timestamp 1676037725
transform 1 0 503516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5473
timestamp 1676037725
transform 1 0 504620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5485
timestamp 1676037725
transform 1 0 505724 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5489
timestamp 1676037725
transform 1 0 506092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5501
timestamp 1676037725
transform 1 0 507196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5513
timestamp 1676037725
transform 1 0 508300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5517
timestamp 1676037725
transform 1 0 508668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5529
timestamp 1676037725
transform 1 0 509772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5541
timestamp 1676037725
transform 1 0 510876 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5545
timestamp 1676037725
transform 1 0 511244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5557
timestamp 1676037725
transform 1 0 512348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5569
timestamp 1676037725
transform 1 0 513452 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5573
timestamp 1676037725
transform 1 0 513820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5585
timestamp 1676037725
transform 1 0 514924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5597
timestamp 1676037725
transform 1 0 516028 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5601
timestamp 1676037725
transform 1 0 516396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5613
timestamp 1676037725
transform 1 0 517500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5625
timestamp 1676037725
transform 1 0 518604 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5629
timestamp 1676037725
transform 1 0 518972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5641
timestamp 1676037725
transform 1 0 520076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5653
timestamp 1676037725
transform 1 0 521180 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5657
timestamp 1676037725
transform 1 0 521548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5669
timestamp 1676037725
transform 1 0 522652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5681
timestamp 1676037725
transform 1 0 523756 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5685
timestamp 1676037725
transform 1 0 524124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5697
timestamp 1676037725
transform 1 0 525228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5709
timestamp 1676037725
transform 1 0 526332 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5713
timestamp 1676037725
transform 1 0 526700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5725
timestamp 1676037725
transform 1 0 527804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5737
timestamp 1676037725
transform 1 0 528908 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5741
timestamp 1676037725
transform 1 0 529276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5753
timestamp 1676037725
transform 1 0 530380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5765
timestamp 1676037725
transform 1 0 531484 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5769
timestamp 1676037725
transform 1 0 531852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5781
timestamp 1676037725
transform 1 0 532956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5793
timestamp 1676037725
transform 1 0 534060 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5797
timestamp 1676037725
transform 1 0 534428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5809
timestamp 1676037725
transform 1 0 535532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5821
timestamp 1676037725
transform 1 0 536636 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5825
timestamp 1676037725
transform 1 0 537004 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5837
timestamp 1676037725
transform 1 0 538108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5849
timestamp 1676037725
transform 1 0 539212 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5853
timestamp 1676037725
transform 1 0 539580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5865
timestamp 1676037725
transform 1 0 540684 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5877
timestamp 1676037725
transform 1 0 541788 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5881
timestamp 1676037725
transform 1 0 542156 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5893
timestamp 1676037725
transform 1 0 543260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5905
timestamp 1676037725
transform 1 0 544364 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5909
timestamp 1676037725
transform 1 0 544732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5921
timestamp 1676037725
transform 1 0 545836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5933
timestamp 1676037725
transform 1 0 546940 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5937
timestamp 1676037725
transform 1 0 547308 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5949
timestamp 1676037725
transform 1 0 548412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5961
timestamp 1676037725
transform 1 0 549516 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5965
timestamp 1676037725
transform 1 0 549884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5977
timestamp 1676037725
transform 1 0 550988 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_5989
timestamp 1676037725
transform 1 0 552092 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5993
timestamp 1676037725
transform 1 0 552460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6005
timestamp 1676037725
transform 1 0 553564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6017
timestamp 1676037725
transform 1 0 554668 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6021
timestamp 1676037725
transform 1 0 555036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6033
timestamp 1676037725
transform 1 0 556140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6045
timestamp 1676037725
transform 1 0 557244 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6049
timestamp 1676037725
transform 1 0 557612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6061
timestamp 1676037725
transform 1 0 558716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6073
timestamp 1676037725
transform 1 0 559820 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6077
timestamp 1676037725
transform 1 0 560188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6089
timestamp 1676037725
transform 1 0 561292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6101
timestamp 1676037725
transform 1 0 562396 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6105
timestamp 1676037725
transform 1 0 562764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6117
timestamp 1676037725
transform 1 0 563868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6129
timestamp 1676037725
transform 1 0 564972 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6133
timestamp 1676037725
transform 1 0 565340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6145
timestamp 1676037725
transform 1 0 566444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6157
timestamp 1676037725
transform 1 0 567548 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6161
timestamp 1676037725
transform 1 0 567916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6173
timestamp 1676037725
transform 1 0 569020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6185
timestamp 1676037725
transform 1 0 570124 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6189
timestamp 1676037725
transform 1 0 570492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6201
timestamp 1676037725
transform 1 0 571596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6213
timestamp 1676037725
transform 1 0 572700 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6217
timestamp 1676037725
transform 1 0 573068 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6229
timestamp 1676037725
transform 1 0 574172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6241
timestamp 1676037725
transform 1 0 575276 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6245
timestamp 1676037725
transform 1 0 575644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6257
timestamp 1676037725
transform 1 0 576748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6269
timestamp 1676037725
transform 1 0 577852 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6273
timestamp 1676037725
transform 1 0 578220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6285
timestamp 1676037725
transform 1 0 579324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6297
timestamp 1676037725
transform 1 0 580428 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6301
timestamp 1676037725
transform 1 0 580796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6313
timestamp 1676037725
transform 1 0 581900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6325
timestamp 1676037725
transform 1 0 583004 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6329
timestamp 1676037725
transform 1 0 583372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6341
timestamp 1676037725
transform 1 0 584476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6353
timestamp 1676037725
transform 1 0 585580 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6357
timestamp 1676037725
transform 1 0 585948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6369
timestamp 1676037725
transform 1 0 587052 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6381
timestamp 1676037725
transform 1 0 588156 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6385
timestamp 1676037725
transform 1 0 588524 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6397
timestamp 1676037725
transform 1 0 589628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6409
timestamp 1676037725
transform 1 0 590732 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6413
timestamp 1676037725
transform 1 0 591100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6425
timestamp 1676037725
transform 1 0 592204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6437
timestamp 1676037725
transform 1 0 593308 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6441
timestamp 1676037725
transform 1 0 593676 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6453
timestamp 1676037725
transform 1 0 594780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6465
timestamp 1676037725
transform 1 0 595884 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6469
timestamp 1676037725
transform 1 0 596252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6481
timestamp 1676037725
transform 1 0 597356 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6493
timestamp 1676037725
transform 1 0 598460 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6497
timestamp 1676037725
transform 1 0 598828 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6509
timestamp 1676037725
transform 1 0 599932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6521
timestamp 1676037725
transform 1 0 601036 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6525
timestamp 1676037725
transform 1 0 601404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6537
timestamp 1676037725
transform 1 0 602508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6549
timestamp 1676037725
transform 1 0 603612 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6553
timestamp 1676037725
transform 1 0 603980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6565
timestamp 1676037725
transform 1 0 605084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6577
timestamp 1676037725
transform 1 0 606188 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6581
timestamp 1676037725
transform 1 0 606556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6593
timestamp 1676037725
transform 1 0 607660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6605
timestamp 1676037725
transform 1 0 608764 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6609
timestamp 1676037725
transform 1 0 609132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6621
timestamp 1676037725
transform 1 0 610236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6633
timestamp 1676037725
transform 1 0 611340 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6637
timestamp 1676037725
transform 1 0 611708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6649
timestamp 1676037725
transform 1 0 612812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6661
timestamp 1676037725
transform 1 0 613916 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6665
timestamp 1676037725
transform 1 0 614284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6677
timestamp 1676037725
transform 1 0 615388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6689
timestamp 1676037725
transform 1 0 616492 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6693
timestamp 1676037725
transform 1 0 616860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6705
timestamp 1676037725
transform 1 0 617964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6717
timestamp 1676037725
transform 1 0 619068 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6721
timestamp 1676037725
transform 1 0 619436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6733
timestamp 1676037725
transform 1 0 620540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6745
timestamp 1676037725
transform 1 0 621644 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6749
timestamp 1676037725
transform 1 0 622012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6761
timestamp 1676037725
transform 1 0 623116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6773
timestamp 1676037725
transform 1 0 624220 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6777
timestamp 1676037725
transform 1 0 624588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6789
timestamp 1676037725
transform 1 0 625692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6801
timestamp 1676037725
transform 1 0 626796 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6805
timestamp 1676037725
transform 1 0 627164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6817
timestamp 1676037725
transform 1 0 628268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6829
timestamp 1676037725
transform 1 0 629372 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6833
timestamp 1676037725
transform 1 0 629740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6845
timestamp 1676037725
transform 1 0 630844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6857
timestamp 1676037725
transform 1 0 631948 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6861
timestamp 1676037725
transform 1 0 632316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6873
timestamp 1676037725
transform 1 0 633420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6885
timestamp 1676037725
transform 1 0 634524 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6889
timestamp 1676037725
transform 1 0 634892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6901
timestamp 1676037725
transform 1 0 635996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6913
timestamp 1676037725
transform 1 0 637100 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6917
timestamp 1676037725
transform 1 0 637468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6929
timestamp 1676037725
transform 1 0 638572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6941
timestamp 1676037725
transform 1 0 639676 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6945
timestamp 1676037725
transform 1 0 640044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6957
timestamp 1676037725
transform 1 0 641148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6969
timestamp 1676037725
transform 1 0 642252 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6973
timestamp 1676037725
transform 1 0 642620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_6985
timestamp 1676037725
transform 1 0 643724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6997
timestamp 1676037725
transform 1 0 644828 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7001
timestamp 1676037725
transform 1 0 645196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7013
timestamp 1676037725
transform 1 0 646300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7025
timestamp 1676037725
transform 1 0 647404 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7029
timestamp 1676037725
transform 1 0 647772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7041
timestamp 1676037725
transform 1 0 648876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7053
timestamp 1676037725
transform 1 0 649980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7057
timestamp 1676037725
transform 1 0 650348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7069
timestamp 1676037725
transform 1 0 651452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7081
timestamp 1676037725
transform 1 0 652556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7085
timestamp 1676037725
transform 1 0 652924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7097
timestamp 1676037725
transform 1 0 654028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7109
timestamp 1676037725
transform 1 0 655132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7113
timestamp 1676037725
transform 1 0 655500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7125
timestamp 1676037725
transform 1 0 656604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7137
timestamp 1676037725
transform 1 0 657708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7141
timestamp 1676037725
transform 1 0 658076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7153
timestamp 1676037725
transform 1 0 659180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7165
timestamp 1676037725
transform 1 0 660284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7169
timestamp 1676037725
transform 1 0 660652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7181
timestamp 1676037725
transform 1 0 661756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7193
timestamp 1676037725
transform 1 0 662860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7197
timestamp 1676037725
transform 1 0 663228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7209
timestamp 1676037725
transform 1 0 664332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7221
timestamp 1676037725
transform 1 0 665436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7225
timestamp 1676037725
transform 1 0 665804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7237
timestamp 1676037725
transform 1 0 666908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7249
timestamp 1676037725
transform 1 0 668012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7253
timestamp 1676037725
transform 1 0 668380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7265
timestamp 1676037725
transform 1 0 669484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7277
timestamp 1676037725
transform 1 0 670588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7281
timestamp 1676037725
transform 1 0 670956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7293
timestamp 1676037725
transform 1 0 672060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7305
timestamp 1676037725
transform 1 0 673164 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7309
timestamp 1676037725
transform 1 0 673532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7321
timestamp 1676037725
transform 1 0 674636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7333
timestamp 1676037725
transform 1 0 675740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7337
timestamp 1676037725
transform 1 0 676108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7349
timestamp 1676037725
transform 1 0 677212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7361
timestamp 1676037725
transform 1 0 678316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7365
timestamp 1676037725
transform 1 0 678684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7377
timestamp 1676037725
transform 1 0 679788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7389
timestamp 1676037725
transform 1 0 680892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7393
timestamp 1676037725
transform 1 0 681260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7405
timestamp 1676037725
transform 1 0 682364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 682824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 682824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 682824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 682824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 682824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 682824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 682824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 682824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 682824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 682824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1676037725
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1676037725
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1676037725
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1676037725
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1676037725
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1676037725
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1676037725
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1676037725
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1676037725
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1676037725
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1676037725
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1676037725
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1676037725
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1676037725
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1676037725
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1676037725
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 119600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 124752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 129904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 135056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 140208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 145360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 150512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 153088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 155664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 160816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 163392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 165968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 168544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 171120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 173696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 176272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 178848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 181424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 184000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 186576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 189152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 191728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 194304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 196880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 199456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 202032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 204608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 207184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 209760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 212336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 214912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 217488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 220064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 222640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 225216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 227792 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 230368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 232944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 235520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 238096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 240672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 243248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 245824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 248400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 250976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 253552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 256128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 258704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 261280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 263856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 266432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 269008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 271584 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 274160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 276736 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 279312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 281888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 284464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 287040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 289616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 292192 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 294768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 297344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 299920 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 302496 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 305072 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 307648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 310224 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 312800 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 315376 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 317952 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 320528 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 323104 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 325680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 328256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 330832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 333408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 335984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 338560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 341136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 343712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 346288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 348864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 351440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 354016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 356592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 359168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 361744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 364320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 366896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 369472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 372048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 374624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 377200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 379776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 382352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 384928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 387504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 390080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 392656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 395232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 397808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 400384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 402960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 405536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 408112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 410688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 413264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 415840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 418416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 420992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 423568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 426144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 428720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 431296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 433872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 436448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 439024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 441600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 444176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 446752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 449328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 451904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 454480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 457056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 459632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 462208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 464784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 467360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 469936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 472512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 475088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 477664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 480240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 482816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 485392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 487968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 490544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 493120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 495696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 498272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 500848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 503424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 506000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 508576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 511152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 513728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 516304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 518880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 521456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 524032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 526608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 529184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 531760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 534336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 536912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 539488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 542064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 544640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 547216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 549792 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 552368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 554944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 557520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 560096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 562672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 565248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 567824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 570400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 572976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 575552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 578128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 580704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 583280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 585856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 588432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 591008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 593584 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 596160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 598736 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 601312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 603888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 606464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 609040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 611616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 614192 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 616768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 619344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 621920 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 624496 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 627072 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 629648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 632224 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 634800 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 637376 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 639952 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 642528 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 645104 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 647680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 650256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 652832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 655408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 657984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 660560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 663136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 665712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 668288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 670864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 673440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 676016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 678592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 681168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 150512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 155664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 160816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 165968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 171120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 176272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 181424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 186576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 191728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 196880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 202032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 207184 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 212336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 217488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 222640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 227792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 232944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 238096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 243248 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 248400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 253552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 258704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 263856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 269008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 274160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 279312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 284464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 289616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 294768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 299920 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 305072 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 310224 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 315376 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 320528 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 325680 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 330832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 335984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 341136 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 346288 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 351440 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 356592 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 361744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 366896 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 372048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 377200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 382352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 387504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 392656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 397808 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 402960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 408112 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 413264 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 418416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 423568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 428720 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 433872 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 439024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 444176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 449328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 454480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 459632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 464784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 469936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 475088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 480240 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 485392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 490544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 495696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 500848 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 506000 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 511152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 516304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 521456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 526608 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 531760 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 536912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 542064 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 547216 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 552368 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 557520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 562672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 567824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 572976 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 578128 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 583280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 588432 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 593584 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 598736 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 603888 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 609040 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 614192 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 619344 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 624496 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 629648 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 634800 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 639952 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 645104 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 650256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 655408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 660560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 665712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 670864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 676016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 681168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 153088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 158240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 163392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 168544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 173696 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 178848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 184000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 189152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 194304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 199456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 204608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 209760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 214912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 220064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 225216 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 230368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 235520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 240672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 245824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 250976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 256128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 261280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 266432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 271584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 276736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 281888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 287040 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 292192 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 297344 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 302496 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 307648 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 312800 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 317952 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 323104 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 328256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 333408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 338560 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 343712 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 348864 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 354016 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 359168 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 364320 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 369472 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 374624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 379776 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 384928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 390080 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 395232 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 400384 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 405536 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 410688 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 415840 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 420992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 426144 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 431296 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 436448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 441600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 446752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 451904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 457056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 462208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 467360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 472512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 477664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 482816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 487968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 493120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 498272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 503424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 508576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 513728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 518880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 524032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 529184 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 534336 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 539488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 544640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 549792 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 554944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 560096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 565248 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 570400 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 575552 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 580704 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 585856 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 591008 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 596160 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 601312 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 606464 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 611616 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 616768 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 621920 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 627072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 632224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 637376 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 642528 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 647680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 652832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 657984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 663136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 668288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 673440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 678592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 150512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 155664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 160816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 165968 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 171120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 176272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 181424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 186576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 191728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 196880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 202032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 207184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 212336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 217488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 222640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 227792 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 232944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 238096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 243248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 248400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 253552 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 258704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 263856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 269008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 274160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 279312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 284464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 289616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 294768 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 299920 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 305072 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 310224 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 315376 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 320528 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 325680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 330832 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 335984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 341136 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 346288 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 351440 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 356592 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 361744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 366896 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 372048 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 377200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 382352 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 387504 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 392656 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 397808 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 402960 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 408112 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 413264 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 418416 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 423568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 428720 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 433872 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 439024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 444176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 449328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 454480 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 459632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 464784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 469936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 475088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 480240 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 485392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 490544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 495696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 500848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 506000 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 511152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 516304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 521456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 526608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 531760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 536912 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 542064 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 547216 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 552368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 557520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 562672 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 567824 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 572976 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 578128 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 583280 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 588432 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 593584 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 598736 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 603888 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 609040 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 614192 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 619344 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 624496 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 629648 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 634800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 639952 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 645104 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 650256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 655408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 660560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 665712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 670864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 676016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 681168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 153088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 158240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 163392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 168544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 173696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 178848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 184000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 189152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 194304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 199456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 204608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 209760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 214912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 220064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 225216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 230368 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 235520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 240672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 245824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 250976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 256128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 261280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 266432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 271584 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 276736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 281888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 287040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 292192 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 297344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 302496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 307648 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 312800 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 317952 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 323104 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 328256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 333408 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 338560 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 343712 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 348864 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 354016 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 359168 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 364320 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 369472 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 374624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 379776 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 384928 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 390080 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 395232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 400384 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 405536 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 410688 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 415840 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 420992 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 426144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 431296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 436448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 441600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 446752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 451904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 457056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 462208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 467360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 472512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 477664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 482816 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 487968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 493120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 498272 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 503424 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 508576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 513728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 518880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 524032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 529184 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 534336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 539488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 544640 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 549792 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 554944 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 560096 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 565248 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 570400 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 575552 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 580704 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 585856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 591008 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 596160 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 601312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 606464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 611616 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 616768 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 621920 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 627072 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 632224 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 637376 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 642528 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 647680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 652832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 657984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 663136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 668288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 673440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 678592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 150512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 155664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 160816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 165968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 171120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 176272 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 181424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 186576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 191728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 196880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 202032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 207184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 212336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 217488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 222640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 227792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 232944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 238096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 243248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 248400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 253552 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 258704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 263856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 269008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 274160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 279312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 284464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 289616 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 294768 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 299920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 305072 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 310224 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 315376 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 320528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 325680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 330832 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 335984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 341136 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 346288 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 351440 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 356592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 361744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 366896 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 372048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 377200 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 382352 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 387504 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 392656 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 397808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 402960 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 408112 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 413264 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 418416 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 423568 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 428720 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 433872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 439024 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 444176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 449328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 454480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 459632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 464784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 469936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 475088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 480240 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 485392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 490544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 495696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 500848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 506000 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 511152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 516304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 521456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 526608 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 531760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 536912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 542064 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 547216 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 552368 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 557520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 562672 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 567824 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 572976 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 578128 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 583280 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 588432 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 593584 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 598736 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 603888 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 609040 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 614192 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 619344 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 624496 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 629648 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 634800 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 639952 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 645104 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 650256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 655408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 660560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 665712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 670864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 676016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 681168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 153088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 158240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 163392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 168544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 173696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 178848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 184000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 189152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 194304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 199456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 204608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 209760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 214912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 220064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 225216 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 230368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 235520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 240672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 245824 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 250976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 256128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 261280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 266432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 271584 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 276736 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 281888 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 287040 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 292192 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 297344 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 302496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 307648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 312800 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 317952 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 323104 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 328256 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 333408 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 338560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 343712 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 348864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 354016 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 359168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 364320 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 369472 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 374624 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 379776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 384928 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 390080 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 395232 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 400384 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 405536 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 410688 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 415840 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 420992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 426144 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 431296 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 436448 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 441600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 446752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 451904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 457056 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 462208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 467360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 472512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 477664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 482816 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 487968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 493120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 498272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 503424 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 508576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 513728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 518880 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 524032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 529184 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 534336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 539488 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 544640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 549792 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 554944 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 560096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 565248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 570400 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 575552 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 580704 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 585856 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 591008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 596160 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 601312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 606464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 611616 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 616768 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 621920 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 627072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 632224 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 637376 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 642528 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 647680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 652832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 657984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 663136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 668288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1676037725
transform 1 0 673440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1676037725
transform 1 0 678592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1676037725
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1676037725
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1676037725
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1676037725
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1676037725
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1676037725
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1676037725
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1676037725
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1676037725
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1676037725
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1676037725
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1676037725
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1676037725
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1676037725
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1676037725
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1676037725
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1676037725
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1676037725
transform 1 0 150512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1676037725
transform 1 0 155664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1676037725
transform 1 0 160816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1676037725
transform 1 0 165968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1676037725
transform 1 0 171120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1676037725
transform 1 0 176272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1676037725
transform 1 0 181424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1676037725
transform 1 0 186576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1676037725
transform 1 0 191728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1676037725
transform 1 0 196880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1676037725
transform 1 0 202032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1676037725
transform 1 0 207184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1676037725
transform 1 0 212336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1676037725
transform 1 0 217488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1676037725
transform 1 0 222640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1676037725
transform 1 0 227792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1676037725
transform 1 0 232944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1676037725
transform 1 0 238096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1676037725
transform 1 0 243248 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1676037725
transform 1 0 248400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1676037725
transform 1 0 253552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1676037725
transform 1 0 258704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1676037725
transform 1 0 263856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1676037725
transform 1 0 269008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1676037725
transform 1 0 274160 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1676037725
transform 1 0 279312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1676037725
transform 1 0 284464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1676037725
transform 1 0 289616 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1676037725
transform 1 0 294768 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1676037725
transform 1 0 299920 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1676037725
transform 1 0 305072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1676037725
transform 1 0 310224 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1676037725
transform 1 0 315376 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1676037725
transform 1 0 320528 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1676037725
transform 1 0 325680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1676037725
transform 1 0 330832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1676037725
transform 1 0 335984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1676037725
transform 1 0 341136 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1676037725
transform 1 0 346288 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1676037725
transform 1 0 351440 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1676037725
transform 1 0 356592 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1676037725
transform 1 0 361744 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1676037725
transform 1 0 366896 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1676037725
transform 1 0 372048 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1676037725
transform 1 0 377200 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1676037725
transform 1 0 382352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1676037725
transform 1 0 387504 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1676037725
transform 1 0 392656 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1676037725
transform 1 0 397808 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1676037725
transform 1 0 402960 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1676037725
transform 1 0 408112 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1676037725
transform 1 0 413264 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1676037725
transform 1 0 418416 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1676037725
transform 1 0 423568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1676037725
transform 1 0 428720 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1676037725
transform 1 0 433872 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1676037725
transform 1 0 439024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1676037725
transform 1 0 444176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1676037725
transform 1 0 449328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1676037725
transform 1 0 454480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1676037725
transform 1 0 459632 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1676037725
transform 1 0 464784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1676037725
transform 1 0 469936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1676037725
transform 1 0 475088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1676037725
transform 1 0 480240 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1676037725
transform 1 0 485392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1676037725
transform 1 0 490544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1676037725
transform 1 0 495696 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1676037725
transform 1 0 500848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1676037725
transform 1 0 506000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1676037725
transform 1 0 511152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1676037725
transform 1 0 516304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1676037725
transform 1 0 521456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1676037725
transform 1 0 526608 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1676037725
transform 1 0 531760 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1676037725
transform 1 0 536912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1676037725
transform 1 0 542064 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1676037725
transform 1 0 547216 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1676037725
transform 1 0 552368 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1676037725
transform 1 0 557520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1676037725
transform 1 0 562672 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1676037725
transform 1 0 567824 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1676037725
transform 1 0 572976 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1676037725
transform 1 0 578128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1676037725
transform 1 0 583280 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1676037725
transform 1 0 588432 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1676037725
transform 1 0 593584 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1676037725
transform 1 0 598736 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1676037725
transform 1 0 603888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1676037725
transform 1 0 609040 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1676037725
transform 1 0 614192 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1676037725
transform 1 0 619344 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1676037725
transform 1 0 624496 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1676037725
transform 1 0 629648 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1676037725
transform 1 0 634800 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1676037725
transform 1 0 639952 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1676037725
transform 1 0 645104 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1676037725
transform 1 0 650256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1676037725
transform 1 0 655408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1676037725
transform 1 0 660560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1676037725
transform 1 0 665712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1676037725
transform 1 0 670864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1676037725
transform 1 0 676016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1676037725
transform 1 0 681168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1676037725
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1676037725
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1676037725
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1676037725
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1676037725
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1676037725
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1676037725
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1676037725
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1676037725
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1676037725
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1676037725
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1676037725
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1676037725
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1676037725
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1676037725
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1676037725
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1676037725
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1676037725
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1676037725
transform 1 0 153088 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1676037725
transform 1 0 158240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1676037725
transform 1 0 163392 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1676037725
transform 1 0 168544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1676037725
transform 1 0 173696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1676037725
transform 1 0 178848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1676037725
transform 1 0 184000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1676037725
transform 1 0 189152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1676037725
transform 1 0 194304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1676037725
transform 1 0 199456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1676037725
transform 1 0 204608 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1676037725
transform 1 0 209760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1676037725
transform 1 0 214912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1676037725
transform 1 0 220064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1676037725
transform 1 0 225216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1676037725
transform 1 0 230368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1676037725
transform 1 0 235520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1676037725
transform 1 0 240672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1676037725
transform 1 0 245824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1676037725
transform 1 0 250976 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1676037725
transform 1 0 256128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1676037725
transform 1 0 261280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1676037725
transform 1 0 266432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1676037725
transform 1 0 271584 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1676037725
transform 1 0 276736 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1676037725
transform 1 0 281888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1676037725
transform 1 0 287040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1676037725
transform 1 0 292192 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1676037725
transform 1 0 297344 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1676037725
transform 1 0 302496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1676037725
transform 1 0 307648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1676037725
transform 1 0 312800 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1676037725
transform 1 0 317952 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1676037725
transform 1 0 323104 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1676037725
transform 1 0 328256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1676037725
transform 1 0 333408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1676037725
transform 1 0 338560 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1676037725
transform 1 0 343712 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1676037725
transform 1 0 348864 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1676037725
transform 1 0 354016 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1676037725
transform 1 0 359168 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1676037725
transform 1 0 364320 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1676037725
transform 1 0 369472 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1676037725
transform 1 0 374624 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1676037725
transform 1 0 379776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1676037725
transform 1 0 384928 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1676037725
transform 1 0 390080 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1676037725
transform 1 0 395232 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1676037725
transform 1 0 400384 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1676037725
transform 1 0 405536 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1676037725
transform 1 0 410688 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1676037725
transform 1 0 415840 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1676037725
transform 1 0 420992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1676037725
transform 1 0 426144 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1676037725
transform 1 0 431296 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1676037725
transform 1 0 436448 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1676037725
transform 1 0 441600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1676037725
transform 1 0 446752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1676037725
transform 1 0 451904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1676037725
transform 1 0 457056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1676037725
transform 1 0 462208 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1676037725
transform 1 0 467360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1676037725
transform 1 0 472512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1676037725
transform 1 0 477664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1676037725
transform 1 0 482816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1676037725
transform 1 0 487968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1676037725
transform 1 0 493120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1676037725
transform 1 0 498272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1676037725
transform 1 0 503424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1676037725
transform 1 0 508576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1676037725
transform 1 0 513728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1676037725
transform 1 0 518880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1676037725
transform 1 0 524032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1676037725
transform 1 0 529184 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1676037725
transform 1 0 534336 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1676037725
transform 1 0 539488 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1676037725
transform 1 0 544640 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1676037725
transform 1 0 549792 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1676037725
transform 1 0 554944 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1676037725
transform 1 0 560096 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1676037725
transform 1 0 565248 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1676037725
transform 1 0 570400 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1676037725
transform 1 0 575552 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1676037725
transform 1 0 580704 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1676037725
transform 1 0 585856 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1676037725
transform 1 0 591008 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1676037725
transform 1 0 596160 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1676037725
transform 1 0 601312 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1676037725
transform 1 0 606464 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1676037725
transform 1 0 611616 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1676037725
transform 1 0 616768 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1676037725
transform 1 0 621920 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1676037725
transform 1 0 627072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1676037725
transform 1 0 632224 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1676037725
transform 1 0 637376 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1676037725
transform 1 0 642528 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1676037725
transform 1 0 647680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1676037725
transform 1 0 652832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1676037725
transform 1 0 657984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1676037725
transform 1 0 663136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1676037725
transform 1 0 668288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1676037725
transform 1 0 673440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1676037725
transform 1 0 678592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1676037725
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1676037725
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1676037725
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1676037725
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1676037725
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1676037725
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1676037725
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1676037725
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1676037725
transform 1 0 44896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1676037725
transform 1 0 50048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1676037725
transform 1 0 55200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1676037725
transform 1 0 60352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1676037725
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1676037725
transform 1 0 65504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1676037725
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1676037725
transform 1 0 70656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1676037725
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1676037725
transform 1 0 75808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1676037725
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1676037725
transform 1 0 80960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1676037725
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1676037725
transform 1 0 86112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1676037725
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1676037725
transform 1 0 91264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1676037725
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1676037725
transform 1 0 96416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1676037725
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1676037725
transform 1 0 101568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1676037725
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1676037725
transform 1 0 106720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1676037725
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1676037725
transform 1 0 111872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1676037725
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1676037725
transform 1 0 117024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1676037725
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1676037725
transform 1 0 122176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1676037725
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1676037725
transform 1 0 127328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1676037725
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1676037725
transform 1 0 132480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1676037725
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1676037725
transform 1 0 137632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1676037725
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1676037725
transform 1 0 142784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1676037725
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1676037725
transform 1 0 147936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1676037725
transform 1 0 150512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1676037725
transform 1 0 153088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1676037725
transform 1 0 155664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1676037725
transform 1 0 158240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1676037725
transform 1 0 160816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1676037725
transform 1 0 163392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1676037725
transform 1 0 165968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1676037725
transform 1 0 168544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1676037725
transform 1 0 171120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1676037725
transform 1 0 173696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1676037725
transform 1 0 176272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1676037725
transform 1 0 178848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1676037725
transform 1 0 181424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1676037725
transform 1 0 184000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1676037725
transform 1 0 186576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1676037725
transform 1 0 189152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1676037725
transform 1 0 191728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1676037725
transform 1 0 194304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1676037725
transform 1 0 196880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1676037725
transform 1 0 199456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1676037725
transform 1 0 202032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1676037725
transform 1 0 204608 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1676037725
transform 1 0 207184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1676037725
transform 1 0 209760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1676037725
transform 1 0 212336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1676037725
transform 1 0 214912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1676037725
transform 1 0 217488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1676037725
transform 1 0 220064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1676037725
transform 1 0 222640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1676037725
transform 1 0 225216 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1676037725
transform 1 0 227792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1676037725
transform 1 0 230368 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1676037725
transform 1 0 232944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1676037725
transform 1 0 235520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1676037725
transform 1 0 238096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1676037725
transform 1 0 240672 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1676037725
transform 1 0 243248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1676037725
transform 1 0 245824 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1676037725
transform 1 0 248400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1676037725
transform 1 0 250976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1676037725
transform 1 0 253552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1676037725
transform 1 0 256128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1676037725
transform 1 0 258704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1676037725
transform 1 0 261280 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1676037725
transform 1 0 263856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1676037725
transform 1 0 266432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1676037725
transform 1 0 269008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1676037725
transform 1 0 271584 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1676037725
transform 1 0 274160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1676037725
transform 1 0 276736 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1676037725
transform 1 0 279312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1676037725
transform 1 0 281888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1676037725
transform 1 0 284464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1676037725
transform 1 0 287040 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1676037725
transform 1 0 289616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1676037725
transform 1 0 292192 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1676037725
transform 1 0 294768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1676037725
transform 1 0 297344 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1676037725
transform 1 0 299920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1676037725
transform 1 0 302496 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1676037725
transform 1 0 305072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1676037725
transform 1 0 307648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1676037725
transform 1 0 310224 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1676037725
transform 1 0 312800 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1676037725
transform 1 0 315376 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1676037725
transform 1 0 317952 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1676037725
transform 1 0 320528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1676037725
transform 1 0 323104 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1676037725
transform 1 0 325680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1676037725
transform 1 0 328256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1676037725
transform 1 0 330832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1676037725
transform 1 0 333408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1676037725
transform 1 0 335984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1676037725
transform 1 0 338560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1676037725
transform 1 0 341136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1676037725
transform 1 0 343712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1676037725
transform 1 0 346288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1676037725
transform 1 0 348864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1676037725
transform 1 0 351440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1676037725
transform 1 0 354016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1676037725
transform 1 0 356592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1676037725
transform 1 0 359168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1676037725
transform 1 0 361744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1676037725
transform 1 0 364320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1676037725
transform 1 0 366896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1676037725
transform 1 0 369472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1676037725
transform 1 0 372048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1676037725
transform 1 0 374624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1676037725
transform 1 0 377200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1676037725
transform 1 0 379776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1676037725
transform 1 0 382352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1676037725
transform 1 0 384928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1676037725
transform 1 0 387504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1676037725
transform 1 0 390080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1676037725
transform 1 0 392656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1676037725
transform 1 0 395232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1676037725
transform 1 0 397808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1676037725
transform 1 0 400384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1676037725
transform 1 0 402960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1676037725
transform 1 0 405536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1676037725
transform 1 0 408112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1676037725
transform 1 0 410688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1676037725
transform 1 0 413264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1676037725
transform 1 0 415840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1676037725
transform 1 0 418416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1676037725
transform 1 0 420992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1676037725
transform 1 0 423568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1676037725
transform 1 0 426144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1676037725
transform 1 0 428720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1676037725
transform 1 0 431296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1676037725
transform 1 0 433872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1676037725
transform 1 0 436448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1676037725
transform 1 0 439024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1676037725
transform 1 0 441600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1676037725
transform 1 0 444176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1676037725
transform 1 0 446752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1676037725
transform 1 0 449328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1676037725
transform 1 0 451904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1676037725
transform 1 0 454480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1676037725
transform 1 0 457056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1676037725
transform 1 0 459632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1676037725
transform 1 0 462208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1676037725
transform 1 0 464784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1676037725
transform 1 0 467360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1676037725
transform 1 0 469936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1676037725
transform 1 0 472512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1676037725
transform 1 0 475088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1676037725
transform 1 0 477664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1676037725
transform 1 0 480240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1676037725
transform 1 0 482816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1676037725
transform 1 0 485392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1676037725
transform 1 0 487968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1676037725
transform 1 0 490544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1676037725
transform 1 0 493120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1676037725
transform 1 0 495696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1676037725
transform 1 0 498272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1676037725
transform 1 0 500848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1676037725
transform 1 0 503424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1676037725
transform 1 0 506000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1676037725
transform 1 0 508576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1676037725
transform 1 0 511152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1676037725
transform 1 0 513728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1676037725
transform 1 0 516304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1676037725
transform 1 0 518880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1676037725
transform 1 0 521456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1676037725
transform 1 0 524032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1676037725
transform 1 0 526608 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1676037725
transform 1 0 529184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1676037725
transform 1 0 531760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1676037725
transform 1 0 534336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1676037725
transform 1 0 536912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1676037725
transform 1 0 539488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1676037725
transform 1 0 542064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1676037725
transform 1 0 544640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1676037725
transform 1 0 547216 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1676037725
transform 1 0 549792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1676037725
transform 1 0 552368 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1676037725
transform 1 0 554944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1676037725
transform 1 0 557520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1676037725
transform 1 0 560096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1676037725
transform 1 0 562672 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1676037725
transform 1 0 565248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1676037725
transform 1 0 567824 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1676037725
transform 1 0 570400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1676037725
transform 1 0 572976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1676037725
transform 1 0 575552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1676037725
transform 1 0 578128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1676037725
transform 1 0 580704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1676037725
transform 1 0 583280 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1676037725
transform 1 0 585856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1676037725
transform 1 0 588432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1676037725
transform 1 0 591008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1676037725
transform 1 0 593584 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1676037725
transform 1 0 596160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1676037725
transform 1 0 598736 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1676037725
transform 1 0 601312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1676037725
transform 1 0 603888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1676037725
transform 1 0 606464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1676037725
transform 1 0 609040 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1676037725
transform 1 0 611616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1676037725
transform 1 0 614192 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1676037725
transform 1 0 616768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1676037725
transform 1 0 619344 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1676037725
transform 1 0 621920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1676037725
transform 1 0 624496 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1676037725
transform 1 0 627072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1676037725
transform 1 0 629648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1676037725
transform 1 0 632224 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1676037725
transform 1 0 634800 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1676037725
transform 1 0 637376 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1676037725
transform 1 0 639952 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1676037725
transform 1 0 642528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1676037725
transform 1 0 645104 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1676037725
transform 1 0 647680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1676037725
transform 1 0 650256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1676037725
transform 1 0 652832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1676037725
transform 1 0 655408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1676037725
transform 1 0 657984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1676037725
transform 1 0 660560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1676037725
transform 1 0 663136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1676037725
transform 1 0 665712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1676037725
transform 1 0 668288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1676037725
transform 1 0 670864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1676037725
transform 1 0 673440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1676037725
transform 1 0 676016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1676037725
transform 1 0 678592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1676037725
transform 1 0 681168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  u_rp\[0\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[1\].u_buf
timestamp 1676037725
transform -1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[2\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[3\].u_buf
timestamp 1676037725
transform -1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[4\].u_buf
timestamp 1676037725
transform -1 0 63940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[5\].u_buf
timestamp 1676037725
transform -1 0 79396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[6\].u_buf
timestamp 1676037725
transform -1 0 94852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[7\].u_buf
timestamp 1676037725
transform -1 0 110308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[8\].u_buf
timestamp 1676037725
transform -1 0 125764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[9\].u_buf
timestamp 1676037725
transform -1 0 141220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[10\].u_buf
timestamp 1676037725
transform -1 0 156676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[11\].u_buf
timestamp 1676037725
transform -1 0 172132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[12\].u_buf
timestamp 1676037725
transform -1 0 187588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[13\].u_buf
timestamp 1676037725
transform -1 0 203044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[14\].u_buf
timestamp 1676037725
transform -1 0 218500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[15\].u_buf
timestamp 1676037725
transform -1 0 233956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[16\].u_buf
timestamp 1676037725
transform -1 0 249412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[17\].u_buf
timestamp 1676037725
transform -1 0 264868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[18\].u_buf
timestamp 1676037725
transform -1 0 280324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[19\].u_buf
timestamp 1676037725
transform -1 0 295780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[20\].u_buf
timestamp 1676037725
transform -1 0 311236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[21\].u_buf
timestamp 1676037725
transform -1 0 326692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[22\].u_buf
timestamp 1676037725
transform -1 0 342148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[23\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 357604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[24\].u_buf
timestamp 1676037725
transform -1 0 373060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[25\].u_buf
timestamp 1676037725
transform -1 0 388516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[26\].u_buf
timestamp 1676037725
transform -1 0 403972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[27\].u_buf
timestamp 1676037725
transform -1 0 419428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[28\].u_buf
timestamp 1676037725
transform -1 0 434884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[29\].u_buf
timestamp 1676037725
transform -1 0 450340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[30\].u_buf
timestamp 1676037725
transform -1 0 465796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[31\].u_buf
timestamp 1676037725
transform -1 0 481252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[32\].u_buf
timestamp 1676037725
transform -1 0 496708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[33\].u_buf
timestamp 1676037725
transform -1 0 512164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[34\].u_buf
timestamp 1676037725
transform -1 0 527620 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[35\].u_buf
timestamp 1676037725
transform -1 0 543076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[36\].u_buf
timestamp 1676037725
transform -1 0 558532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[37\].u_buf
timestamp 1676037725
transform -1 0 573988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[38\].u_buf
timestamp 1676037725
transform -1 0 589444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[39\].u_buf
timestamp 1676037725
transform -1 0 604900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[40\].u_buf
timestamp 1676037725
transform -1 0 620356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[41\].u_buf
timestamp 1676037725
transform -1 0 635812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[42\].u_buf
timestamp 1676037725
transform -1 0 651268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[43\].u_buf
timestamp 1676037725
transform -1 0 666724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[44\].u_buf
timestamp 1676037725
transform -1 0 682180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  wire1
timestamp 1676037725
transform 1 0 138092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  wire2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 136528 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 342240 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire4
timestamp 1676037725
transform -1 0 436080 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire5
timestamp 1676037725
transform -1 0 530472 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire6
timestamp 1676037725
transform -1 0 625600 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire7
timestamp 1676037725
transform -1 0 339756 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire8
timestamp 1676037725
transform -1 0 434976 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire9
timestamp 1676037725
transform -1 0 529000 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire10
timestamp 1676037725
transform -1 0 623392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire11
timestamp 1676037725
transform -1 0 338376 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire12
timestamp 1676037725
transform -1 0 433596 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire13
timestamp 1676037725
transform -1 0 527712 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire14
timestamp 1676037725
transform -1 0 337548 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire15
timestamp 1676037725
transform -1 0 432400 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire16
timestamp 1676037725
transform -1 0 525964 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire17
timestamp 1676037725
transform -1 0 335800 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire18
timestamp 1676037725
transform -1 0 430468 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire19
timestamp 1676037725
transform 1 0 135332 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire20
timestamp 1676037725
transform 1 0 40756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire21
timestamp 1676037725
transform -1 0 334788 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire22
timestamp 1676037725
transform -1 0 428536 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire23
timestamp 1676037725
transform -1 0 333224 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire24
timestamp 1676037725
transform -1 0 331660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire25
timestamp 1676037725
transform -1 0 204240 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire26
timestamp 1676037725
transform -1 0 188968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire27
timestamp 1676037725
transform -1 0 159344 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  wire28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 571320 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 477940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire30
timestamp 1676037725
transform 1 0 382996 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire31
timestamp 1676037725
transform 1 0 288512 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  wire32
timestamp 1676037725
transform 1 0 555864 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  wire33
timestamp 1676037725
transform 1 0 462484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  wire34
timestamp 1676037725
transform 1 0 367632 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire35
timestamp 1676037725
transform 1 0 273056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire36
timestamp 1676037725
transform 1 0 525596 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire37
timestamp 1676037725
transform 1 0 431296 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire38
timestamp 1676037725
transform 1 0 336352 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire39
timestamp 1676037725
transform -1 0 143888 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire40
timestamp 1676037725
transform 1 0 510140 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire41
timestamp 1676037725
transform 1 0 416116 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire42
timestamp 1676037725
transform 1 0 321448 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire43
timestamp 1676037725
transform 1 0 479228 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire44
timestamp 1676037725
transform 1 0 385204 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire45
timestamp 1676037725
transform 1 0 290628 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire46
timestamp 1676037725
transform 1 0 463772 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire47
timestamp 1676037725
transform 1 0 369748 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire48
timestamp 1676037725
transform 1 0 275264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire49
timestamp 1676037725
transform 1 0 432860 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire50
timestamp 1676037725
transform 1 0 338928 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire51
timestamp 1676037725
transform 1 0 417404 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire52
timestamp 1676037725
transform 1 0 323472 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire53
timestamp 1676037725
transform 1 0 386492 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire54
timestamp 1676037725
transform 1 0 292744 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire55
timestamp 1676037725
transform 1 0 371036 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire56
timestamp 1676037725
transform 1 0 277380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire57
timestamp 1676037725
transform 1 0 340124 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire58
timestamp 1676037725
transform 1 0 246744 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire59
timestamp 1676037725
transform 1 0 324668 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire60
timestamp 1676037725
transform 1 0 295044 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire61
timestamp 1676037725
transform 1 0 279588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  wire62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 248860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire63
timestamp 1676037725
transform -1 0 112976 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire64
timestamp 1676037725
transform -1 0 206264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire65
timestamp 1676037725
transform -1 0 97520 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire66
timestamp 1676037725
transform -1 0 190900 0 1 2176
box -38 -48 590 592
<< labels >>
flabel metal1 s 228010 0 228066 800 0 FreeSans 224 90 0 0 ch_in[0]
port 0 nsew signal input
flabel metal1 s 232090 0 232146 800 0 FreeSans 224 90 0 0 ch_in[10]
port 1 nsew signal input
flabel metal1 s 168374 9200 168430 10000 0 FreeSans 224 90 0 0 ch_in[11]
port 2 nsew signal input
flabel metal1 s 232906 0 232962 800 0 FreeSans 224 90 0 0 ch_in[12]
port 3 nsew signal input
flabel metal1 s 233314 0 233370 800 0 FreeSans 224 90 0 0 ch_in[13]
port 4 nsew signal input
flabel metal1 s 214274 9200 214330 10000 0 FreeSans 224 90 0 0 ch_in[14]
port 5 nsew signal input
flabel metal1 s 234130 0 234186 800 0 FreeSans 224 90 0 0 ch_in[15]
port 6 nsew signal input
flabel metal1 s 234538 0 234594 800 0 FreeSans 224 90 0 0 ch_in[16]
port 7 nsew signal input
flabel metal1 s 260174 9200 260230 10000 0 FreeSans 224 90 0 0 ch_in[17]
port 8 nsew signal input
flabel metal1 s 235354 0 235410 800 0 FreeSans 224 90 0 0 ch_in[18]
port 9 nsew signal input
flabel metal1 s 235762 0 235818 800 0 FreeSans 224 90 0 0 ch_in[19]
port 10 nsew signal input
flabel metal1 s 228418 0 228474 800 0 FreeSans 224 90 0 0 ch_in[1]
port 11 nsew signal input
flabel metal1 s 306074 9200 306130 10000 0 FreeSans 224 90 0 0 ch_in[20]
port 12 nsew signal input
flabel metal1 s 236578 0 236634 800 0 FreeSans 224 90 0 0 ch_in[21]
port 13 nsew signal input
flabel metal1 s 236986 0 237042 800 0 FreeSans 224 90 0 0 ch_in[22]
port 14 nsew signal input
flabel metal1 s 351974 9200 352030 10000 0 FreeSans 224 90 0 0 ch_in[23]
port 15 nsew signal input
flabel metal1 s 237802 0 237858 800 0 FreeSans 224 90 0 0 ch_in[24]
port 16 nsew signal input
flabel metal1 s 238210 0 238266 800 0 FreeSans 224 90 0 0 ch_in[25]
port 17 nsew signal input
flabel metal1 s 397874 9200 397930 10000 0 FreeSans 224 90 0 0 ch_in[26]
port 18 nsew signal input
flabel metal1 s 239026 0 239082 800 0 FreeSans 224 90 0 0 ch_in[27]
port 19 nsew signal input
flabel metal1 s 239434 0 239490 800 0 FreeSans 224 90 0 0 ch_in[28]
port 20 nsew signal input
flabel metal1 s 443774 9200 443830 10000 0 FreeSans 224 90 0 0 ch_in[29]
port 21 nsew signal input
flabel metal1 s 30674 9200 30730 10000 0 FreeSans 224 90 0 0 ch_in[2]
port 22 nsew signal input
flabel metal1 s 240250 0 240306 800 0 FreeSans 224 90 0 0 ch_in[30]
port 23 nsew signal input
flabel metal1 s 240658 0 240714 800 0 FreeSans 224 90 0 0 ch_in[31]
port 24 nsew signal input
flabel metal1 s 489674 9200 489730 10000 0 FreeSans 224 90 0 0 ch_in[32]
port 25 nsew signal input
flabel metal1 s 241474 0 241530 800 0 FreeSans 224 90 0 0 ch_in[33]
port 26 nsew signal input
flabel metal1 s 241882 0 241938 800 0 FreeSans 224 90 0 0 ch_in[34]
port 27 nsew signal input
flabel metal1 s 535574 9200 535630 10000 0 FreeSans 224 90 0 0 ch_in[35]
port 28 nsew signal input
flabel metal1 s 242698 0 242754 800 0 FreeSans 224 90 0 0 ch_in[36]
port 29 nsew signal input
flabel metal1 s 243106 0 243162 800 0 FreeSans 224 90 0 0 ch_in[37]
port 30 nsew signal input
flabel metal1 s 581474 9200 581530 10000 0 FreeSans 224 90 0 0 ch_in[38]
port 31 nsew signal input
flabel metal1 s 243922 0 243978 800 0 FreeSans 224 90 0 0 ch_in[39]
port 32 nsew signal input
flabel metal1 s 229234 0 229290 800 0 FreeSans 224 90 0 0 ch_in[3]
port 33 nsew signal input
flabel metal1 s 244330 0 244386 800 0 FreeSans 224 90 0 0 ch_in[40]
port 34 nsew signal input
flabel metal1 s 627374 9200 627430 10000 0 FreeSans 224 90 0 0 ch_in[41]
port 35 nsew signal input
flabel metal1 s 245146 0 245202 800 0 FreeSans 224 90 0 0 ch_in[42]
port 36 nsew signal input
flabel metal1 s 245554 0 245610 800 0 FreeSans 224 90 0 0 ch_in[43]
port 37 nsew signal input
flabel metal1 s 673274 9200 673330 10000 0 FreeSans 224 90 0 0 ch_in[44]
port 38 nsew signal input
flabel metal1 s 229642 0 229698 800 0 FreeSans 224 90 0 0 ch_in[4]
port 39 nsew signal input
flabel metal1 s 76574 9200 76630 10000 0 FreeSans 224 90 0 0 ch_in[5]
port 40 nsew signal input
flabel metal1 s 230458 0 230514 800 0 FreeSans 224 90 0 0 ch_in[6]
port 41 nsew signal input
flabel metal1 s 230866 0 230922 800 0 FreeSans 224 90 0 0 ch_in[7]
port 42 nsew signal input
flabel metal1 s 122474 9200 122530 10000 0 FreeSans 224 90 0 0 ch_in[8]
port 43 nsew signal input
flabel metal1 s 231682 0 231738 800 0 FreeSans 224 90 0 0 ch_in[9]
port 44 nsew signal input
flabel metal1 s 74 9200 130 10000 0 FreeSans 224 90 0 0 ch_out[0]
port 45 nsew signal tristate
flabel metal1 s 153074 9200 153130 10000 0 FreeSans 224 90 0 0 ch_out[10]
port 46 nsew signal tristate
flabel metal1 s 232498 0 232554 800 0 FreeSans 224 90 0 0 ch_out[11]
port 47 nsew signal tristate
flabel metal1 s 183674 9200 183730 10000 0 FreeSans 224 90 0 0 ch_out[12]
port 48 nsew signal tristate
flabel metal1 s 198974 9200 199030 10000 0 FreeSans 224 90 0 0 ch_out[13]
port 49 nsew signal tristate
flabel metal1 s 233722 0 233778 800 0 FreeSans 224 90 0 0 ch_out[14]
port 50 nsew signal tristate
flabel metal1 s 229574 9200 229630 10000 0 FreeSans 224 90 0 0 ch_out[15]
port 51 nsew signal tristate
flabel metal1 s 244874 9200 244930 10000 0 FreeSans 224 90 0 0 ch_out[16]
port 52 nsew signal tristate
flabel metal1 s 234946 0 235002 800 0 FreeSans 224 90 0 0 ch_out[17]
port 53 nsew signal tristate
flabel metal1 s 275474 9200 275530 10000 0 FreeSans 224 90 0 0 ch_out[18]
port 54 nsew signal tristate
flabel metal1 s 290774 9200 290830 10000 0 FreeSans 224 90 0 0 ch_out[19]
port 55 nsew signal tristate
flabel metal1 s 15374 9200 15430 10000 0 FreeSans 224 90 0 0 ch_out[1]
port 56 nsew signal tristate
flabel metal1 s 236170 0 236226 800 0 FreeSans 224 90 0 0 ch_out[20]
port 57 nsew signal tristate
flabel metal1 s 321374 9200 321430 10000 0 FreeSans 224 90 0 0 ch_out[21]
port 58 nsew signal tristate
flabel metal1 s 336674 9200 336730 10000 0 FreeSans 224 90 0 0 ch_out[22]
port 59 nsew signal tristate
flabel metal1 s 237394 0 237450 800 0 FreeSans 224 90 0 0 ch_out[23]
port 60 nsew signal tristate
flabel metal1 s 367274 9200 367330 10000 0 FreeSans 224 90 0 0 ch_out[24]
port 61 nsew signal tristate
flabel metal1 s 382574 9200 382630 10000 0 FreeSans 224 90 0 0 ch_out[25]
port 62 nsew signal tristate
flabel metal1 s 238618 0 238674 800 0 FreeSans 224 90 0 0 ch_out[26]
port 63 nsew signal tristate
flabel metal1 s 413174 9200 413230 10000 0 FreeSans 224 90 0 0 ch_out[27]
port 64 nsew signal tristate
flabel metal1 s 428474 9200 428530 10000 0 FreeSans 224 90 0 0 ch_out[28]
port 65 nsew signal tristate
flabel metal1 s 239842 0 239898 800 0 FreeSans 224 90 0 0 ch_out[29]
port 66 nsew signal tristate
flabel metal1 s 228826 0 228882 800 0 FreeSans 224 90 0 0 ch_out[2]
port 67 nsew signal tristate
flabel metal1 s 459074 9200 459130 10000 0 FreeSans 224 90 0 0 ch_out[30]
port 68 nsew signal tristate
flabel metal1 s 474374 9200 474430 10000 0 FreeSans 224 90 0 0 ch_out[31]
port 69 nsew signal tristate
flabel metal1 s 241066 0 241122 800 0 FreeSans 224 90 0 0 ch_out[32]
port 70 nsew signal tristate
flabel metal1 s 504974 9200 505030 10000 0 FreeSans 224 90 0 0 ch_out[33]
port 71 nsew signal tristate
flabel metal1 s 520274 9200 520330 10000 0 FreeSans 224 90 0 0 ch_out[34]
port 72 nsew signal tristate
flabel metal1 s 242290 0 242346 800 0 FreeSans 224 90 0 0 ch_out[35]
port 73 nsew signal tristate
flabel metal1 s 550874 9200 550930 10000 0 FreeSans 224 90 0 0 ch_out[36]
port 74 nsew signal tristate
flabel metal1 s 566174 9200 566230 10000 0 FreeSans 224 90 0 0 ch_out[37]
port 75 nsew signal tristate
flabel metal1 s 243514 0 243570 800 0 FreeSans 224 90 0 0 ch_out[38]
port 76 nsew signal tristate
flabel metal1 s 596774 9200 596830 10000 0 FreeSans 224 90 0 0 ch_out[39]
port 77 nsew signal tristate
flabel metal1 s 45974 9200 46030 10000 0 FreeSans 224 90 0 0 ch_out[3]
port 78 nsew signal tristate
flabel metal1 s 612074 9200 612130 10000 0 FreeSans 224 90 0 0 ch_out[40]
port 79 nsew signal tristate
flabel metal1 s 244738 0 244794 800 0 FreeSans 224 90 0 0 ch_out[41]
port 80 nsew signal tristate
flabel metal1 s 642674 9200 642730 10000 0 FreeSans 224 90 0 0 ch_out[42]
port 81 nsew signal tristate
flabel metal1 s 657974 9200 658030 10000 0 FreeSans 224 90 0 0 ch_out[43]
port 82 nsew signal tristate
flabel metal1 s 245962 0 246018 800 0 FreeSans 224 90 0 0 ch_out[44]
port 83 nsew signal tristate
flabel metal1 s 61274 9200 61330 10000 0 FreeSans 224 90 0 0 ch_out[4]
port 84 nsew signal tristate
flabel metal1 s 230050 0 230106 800 0 FreeSans 224 90 0 0 ch_out[5]
port 85 nsew signal tristate
flabel metal1 s 91874 9200 91930 10000 0 FreeSans 224 90 0 0 ch_out[6]
port 86 nsew signal tristate
flabel metal1 s 107174 9200 107230 10000 0 FreeSans 224 90 0 0 ch_out[7]
port 87 nsew signal tristate
flabel metal1 s 231274 0 231330 800 0 FreeSans 224 90 0 0 ch_out[8]
port 88 nsew signal tristate
flabel metal1 s 137774 9200 137830 10000 0 FreeSans 224 90 0 0 ch_out[9]
port 89 nsew signal tristate
flabel metal2 s -416 656 -96 9136 0 FreeSans 1792 90 0 0 vccd1
port 90 nsew power bidirectional
flabel metal3 s -416 656 684344 976 0 FreeSans 1920 0 0 0 vccd1
port 90 nsew power bidirectional
flabel metal3 s -416 8816 684344 9136 0 FreeSans 1920 0 0 0 vccd1
port 90 nsew power bidirectional
flabel metal2 s 684024 656 684344 9136 0 FreeSans 1792 90 0 0 vccd1
port 90 nsew power bidirectional
flabel metal2 s 86159 -4 86479 9796 0 FreeSans 1792 90 0 0 vccd1
port 90 nsew power bidirectional
flabel metal2 s 256589 -4 256909 9796 0 FreeSans 1792 90 0 0 vccd1
port 90 nsew power bidirectional
flabel metal2 s 427019 -4 427339 9796 0 FreeSans 1792 90 0 0 vccd1
port 90 nsew power bidirectional
flabel metal2 s 597449 -4 597769 9796 0 FreeSans 1792 90 0 0 vccd1
port 90 nsew power bidirectional
flabel metal3 s -1076 2695 685004 3015 0 FreeSans 1920 0 0 0 vccd1
port 90 nsew power bidirectional
flabel metal3 s -1076 4054 685004 4374 0 FreeSans 1920 0 0 0 vccd1
port 90 nsew power bidirectional
flabel metal3 s -1076 5413 685004 5733 0 FreeSans 1920 0 0 0 vccd1
port 90 nsew power bidirectional
flabel metal3 s -1076 6772 685004 7092 0 FreeSans 1920 0 0 0 vccd1
port 90 nsew power bidirectional
flabel metal2 s -1076 -4 -756 9796 0 FreeSans 1792 90 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal3 s -1076 -4 685004 316 0 FreeSans 1920 0 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal3 s -1076 9476 685004 9796 0 FreeSans 1920 0 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal2 s 684684 -4 685004 9796 0 FreeSans 1792 90 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal2 s 86819 -4 87139 9796 0 FreeSans 1792 90 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal2 s 257249 -4 257569 9796 0 FreeSans 1792 90 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal2 s 427679 -4 427999 9796 0 FreeSans 1792 90 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal2 s 598109 -4 598429 9796 0 FreeSans 1792 90 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal3 s -1076 3355 685004 3675 0 FreeSans 1920 0 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal3 s -1076 4714 685004 5034 0 FreeSans 1920 0 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal3 s -1076 6073 685004 6393 0 FreeSans 1920 0 0 0 vssd1
port 91 nsew ground bidirectional
flabel metal3 s -1076 7432 685004 7752 0 FreeSans 1920 0 0 0 vssd1
port 91 nsew ground bidirectional
rlabel metal1 341964 7072 341964 7072 0 vccd1
rlabel metal1 341964 7616 341964 7616 0 vssd1
rlabel metal2 191406 1156 191406 1156 0 ch_in[0]
rlabel metal2 157182 1700 157182 1700 0 ch_in[10]
rlabel metal2 171626 4998 171626 4998 0 ch_in[11]
rlabel metal1 190854 2312 190854 2312 0 ch_in[12]
rlabel metal2 202998 1292 202998 1292 0 ch_in[13]
rlabel metal2 218086 4998 218086 4998 0 ch_in[14]
rlabel metal2 234370 1530 234370 1530 0 ch_in[15]
rlabel metal1 246192 2618 246192 2618 0 ch_in[16]
rlabel metal2 264362 4930 264362 4930 0 ch_in[17]
rlabel metal2 278990 2142 278990 2142 0 ch_in[18]
rlabel metal1 235918 782 235918 782 0 ch_in[19]
rlabel metal1 206494 2414 206494 2414 0 ch_in[1]
rlabel metal2 310730 4590 310730 4590 0 ch_in[20]
rlabel metal2 326186 2669 326186 2669 0 ch_in[21]
rlabel metal1 248722 3026 248722 3026 0 ch_in[22]
rlabel metal1 352613 8874 352613 8874 0 ch_in[23]
rlabel metal1 279634 3060 279634 3060 0 ch_in[24]
rlabel metal1 294814 3026 294814 3026 0 ch_in[25]
rlabel metal2 403466 4998 403466 4998 0 ch_in[26]
rlabel metal1 291134 2414 291134 2414 0 ch_in[27]
rlabel metal1 246514 2414 246514 2414 0 ch_in[28]
rlabel metal2 449926 4964 449926 4964 0 ch_in[29]
rlabel metal1 32292 2414 32292 2414 0 ch_in[2]
rlabel metal2 276046 2040 276046 2040 0 ch_in[30]
rlabel metal1 292790 2822 292790 2822 0 ch_in[31]
rlabel metal1 489785 8942 489785 8942 0 ch_in[32]
rlabel metal2 323610 1904 323610 1904 0 ch_in[33]
rlabel metal1 338744 3026 338744 3026 0 ch_in[34]
rlabel metal1 542570 2414 542570 2414 0 ch_in[35]
rlabel metal2 274758 2176 274758 2176 0 ch_in[36]
rlabel metal2 290214 2142 290214 2142 0 ch_in[37]
rlabel metal1 581915 9214 581915 9214 0 ch_in[38]
rlabel metal2 320942 2040 320942 2040 0 ch_in[39]
rlabel metal1 224066 952 224066 952 0 ch_in[3]
rlabel metal2 336490 1496 336490 1496 0 ch_in[40]
rlabel metal2 635582 4284 635582 4284 0 ch_in[41]
rlabel metal2 272550 1292 272550 1292 0 ch_in[42]
rlabel metal2 288006 1224 288006 1224 0 ch_in[43]
rlabel metal2 681766 4658 681766 4658 0 ch_in[44]
rlabel metal2 159850 1734 159850 1734 0 ch_in[4]
rlabel metal2 78890 4998 78890 4998 0 ch_in[5]
rlabel metal2 189566 1870 189566 1870 0 ch_in[6]
rlabel metal1 204608 2414 204608 2414 0 ch_in[7]
rlabel metal1 122643 9214 122643 9214 0 ch_in[8]
rlabel metal1 223974 884 223974 884 0 ch_in[9]
rlabel metal1 996 9214 996 9214 0 ch_out[0]
rlabel metal1 156170 2550 156170 2550 0 ch_out[10]
rlabel metal2 171902 1768 171902 1768 0 ch_out[11]
rlabel metal2 187358 4726 187358 4726 0 ch_out[12]
rlabel metal1 199525 8942 199525 8942 0 ch_out[13]
rlabel metal2 218270 2312 218270 2312 0 ch_out[14]
rlabel metal1 231748 6834 231748 6834 0 ch_out[15]
rlabel metal1 247388 6834 247388 6834 0 ch_out[16]
rlabel metal2 264638 1258 264638 1258 0 ch_out[17]
rlabel metal1 275731 9214 275731 9214 0 ch_out[18]
rlabel metal1 293342 6834 293342 6834 0 ch_out[19]
rlabel metal1 16974 2618 16974 2618 0 ch_out[1]
rlabel metal2 311006 1190 311006 1190 0 ch_out[20]
rlabel metal2 326462 4556 326462 4556 0 ch_out[21]
rlabel metal2 341918 4556 341918 4556 0 ch_out[22]
rlabel metal2 331338 1802 331338 1802 0 ch_out[23]
rlabel metal2 372830 4692 372830 4692 0 ch_out[24]
rlabel metal2 388286 4352 388286 4352 0 ch_out[25]
rlabel metal2 332626 1700 332626 1700 0 ch_out[26]
rlabel metal2 419198 4556 419198 4556 0 ch_out[27]
rlabel metal1 428819 9214 428819 9214 0 ch_out[28]
rlabel metal2 334098 1598 334098 1598 0 ch_out[29]
rlabel metal2 224250 969 224250 969 0 ch_out[2]
rlabel metal1 465290 2278 465290 2278 0 ch_out[30]
rlabel metal1 476790 6834 476790 6834 0 ch_out[31]
rlabel metal2 335478 1632 335478 1632 0 ch_out[32]
rlabel via1 505011 8942 505011 8942 0 ch_out[33]
rlabel metal1 527252 2278 527252 2278 0 ch_out[34]
rlabel metal2 336858 1972 336858 1972 0 ch_out[35]
rlabel metal1 554070 6834 554070 6834 0 ch_out[36]
rlabel metal1 566681 9214 566681 9214 0 ch_out[37]
rlabel metal2 337686 1734 337686 1734 0 ch_out[38]
rlabel metal2 604670 4726 604670 4726 0 ch_out[39]
rlabel metal1 47610 2618 47610 2618 0 ch_out[3]
rlabel metal2 620126 4386 620126 4386 0 ch_out[40]
rlabel metal2 339066 1394 339066 1394 0 ch_out[41]
rlabel metal1 642873 8942 642873 8942 0 ch_out[42]
rlabel metal1 658108 8942 658108 8942 0 ch_out[43]
rlabel metal2 341550 1496 341550 1496 0 ch_out[44]
rlabel metal2 63710 4726 63710 4726 0 ch_out[4]
rlabel metal2 224158 289 224158 289 0 ch_out[5]
rlabel metal2 94622 4726 94622 4726 0 ch_out[6]
rlabel metal2 110078 4556 110078 4556 0 ch_out[7]
rlabel metal1 219420 748 219420 748 0 ch_out[8]
rlabel metal1 139334 6834 139334 6834 0 ch_out[9]
rlabel metal2 125718 2108 125718 2108 0 net1
rlabel metal2 623070 2108 623070 2108 0 net10
rlabel metal2 528218 2448 528218 2448 0 net11
rlabel metal2 338238 1870 338238 1870 0 net12
rlabel metal2 527022 3230 527022 3230 0 net13
rlabel metal1 525918 3060 525918 3060 0 net14
rlabel metal2 431710 2924 431710 2924 0 net15
rlabel metal1 525642 3128 525642 3128 0 net16
rlabel metal2 430974 2006 430974 2006 0 net17
rlabel metal2 429778 1802 429778 1802 0 net18
rlabel metal1 38341 2414 38341 2414 0 net19
rlabel metal2 79166 2142 79166 2142 0 net2
rlabel metal1 43309 2482 43309 2482 0 net20
rlabel metal2 429134 2142 429134 2142 0 net21
rlabel metal2 334650 1802 334650 1802 0 net22
rlabel metal2 333086 1734 333086 1734 0 net23
rlabel metal2 331614 2074 331614 2074 0 net24
rlabel metal2 110722 2176 110722 2176 0 net25
rlabel metal2 95358 2040 95358 2040 0 net26
rlabel metal1 64170 2414 64170 2414 0 net27
rlabel metal1 623162 2414 623162 2414 0 net28
rlabel metal1 526378 2414 526378 2414 0 net29
rlabel metal2 625462 2516 625462 2516 0 net3
rlabel metal2 383686 1972 383686 1972 0 net30
rlabel metal1 288834 2312 288834 2312 0 net31
rlabel metal1 620310 2312 620310 2312 0 net32
rlabel metal2 463358 2176 463358 2176 0 net33
rlabel metal2 368322 1734 368322 1734 0 net34
rlabel metal2 273378 2516 273378 2516 0 net35
rlabel metal1 526286 2482 526286 2482 0 net36
rlabel metal2 431894 2737 431894 2737 0 net37
rlabel metal2 430790 2601 430790 2601 0 net38
rlabel metal1 48438 2482 48438 2482 0 net39
rlabel metal2 342746 2312 342746 2312 0 net4
rlabel metal2 604486 2720 604486 2720 0 net40
rlabel metal2 416806 2210 416806 2210 0 net41
rlabel metal2 322138 2176 322138 2176 0 net42
rlabel metal1 526010 2992 526010 2992 0 net43
rlabel metal1 389597 2482 389597 2482 0 net44
rlabel metal2 290950 2210 290950 2210 0 net45
rlabel metal2 558118 2618 558118 2618 0 net46
rlabel metal2 370438 2108 370438 2108 0 net47
rlabel metal2 275586 1972 275586 1972 0 net48
rlabel metal2 527574 2924 527574 2924 0 net49
rlabel metal2 436862 2040 436862 2040 0 net5
rlabel metal2 339618 3264 339618 3264 0 net50
rlabel metal1 463266 2380 463266 2380 0 net51
rlabel metal2 324162 2006 324162 2006 0 net52
rlabel metal2 387182 1904 387182 1904 0 net53
rlabel metal2 386630 2176 386630 2176 0 net54
rlabel metal1 371726 2516 371726 2516 0 net55
rlabel metal1 370760 2414 370760 2414 0 net56
rlabel metal2 340814 1870 340814 1870 0 net57
rlabel metal2 340262 1938 340262 1938 0 net58
rlabel metal2 325358 1938 325358 1938 0 net59
rlabel metal2 624910 2142 624910 2142 0 net6
rlabel metal2 388470 2754 388470 2754 0 net60
rlabel metal2 373014 2652 373014 2652 0 net61
rlabel metal1 342102 2482 342102 2482 0 net62
rlabel metal2 18078 2108 18078 2108 0 net63
rlabel metal2 113482 2006 113482 2006 0 net64
rlabel metal2 2622 2176 2622 2176 0 net65
rlabel metal2 97382 2516 97382 2516 0 net66
rlabel metal1 623254 2482 623254 2482 0 net7
rlabel metal2 426926 3264 426926 3264 0 net8
rlabel metal2 528310 2006 528310 2006 0 net9
<< properties >>
string FIXED_BBOX 0 0 684000 10000
<< end >>
