magic
tech sky130A
magscale 1 2
timestamp 1698826257
<< viali >>
rect 2421 17221 2455 17255
rect 2605 17221 2639 17255
rect 4169 17221 4203 17255
rect 3065 17153 3099 17187
rect 3341 17153 3375 17187
rect 4353 17153 4387 17187
rect 4905 17153 4939 17187
rect 5089 17153 5123 17187
rect 3433 17085 3467 17119
rect 2237 17017 2271 17051
rect 3985 17017 4019 17051
rect 5089 17017 5123 17051
rect 2421 16949 2455 16983
rect 6377 16677 6411 16711
rect 1593 16541 1627 16575
rect 1869 16541 1903 16575
rect 2697 16541 2731 16575
rect 4169 16541 4203 16575
rect 5365 16541 5399 16575
rect 5457 16541 5491 16575
rect 6285 16541 6319 16575
rect 6469 16541 6503 16575
rect 1961 16473 1995 16507
rect 2421 16473 2455 16507
rect 2881 16473 2915 16507
rect 3985 16473 4019 16507
rect 4353 16473 4387 16507
rect 2513 16405 2547 16439
rect 5549 16405 5583 16439
rect 2237 16133 2271 16167
rect 4445 16133 4479 16167
rect 4629 16133 4663 16167
rect 5641 16133 5675 16167
rect 6745 16133 6779 16167
rect 2145 16065 2179 16099
rect 2421 16065 2455 16099
rect 3433 16065 3467 16099
rect 3525 16065 3559 16099
rect 3709 16065 3743 16099
rect 5825 16065 5859 16099
rect 6929 16065 6963 16099
rect 7481 16065 7515 16099
rect 7665 16065 7699 16099
rect 3893 15929 3927 15963
rect 7665 15929 7699 15963
rect 2605 15861 2639 15895
rect 4629 15861 4663 15895
rect 4813 15861 4847 15895
rect 5549 15861 5583 15895
rect 6653 15861 6687 15895
rect 5365 15657 5399 15691
rect 6193 15657 6227 15691
rect 3065 15589 3099 15623
rect 4445 15521 4479 15555
rect 9137 15521 9171 15555
rect 1961 15453 1995 15487
rect 2697 15453 2731 15487
rect 3065 15453 3099 15487
rect 3249 15453 3283 15487
rect 3985 15453 4019 15487
rect 4077 15453 4111 15487
rect 4261 15453 4295 15487
rect 5641 15453 5675 15487
rect 9321 15453 9355 15487
rect 9413 15453 9447 15487
rect 1685 15385 1719 15419
rect 2145 15385 2179 15419
rect 5181 15385 5215 15419
rect 6285 15385 6319 15419
rect 6469 15385 6503 15419
rect 6929 15385 6963 15419
rect 7113 15385 7147 15419
rect 7297 15385 7331 15419
rect 8125 15385 8159 15419
rect 8309 15385 8343 15419
rect 8493 15385 8527 15419
rect 1777 15317 1811 15351
rect 5365 15317 5399 15351
rect 1869 15113 1903 15147
rect 3617 15113 3651 15147
rect 6929 15113 6963 15147
rect 1777 15045 1811 15079
rect 6561 15045 6595 15079
rect 6745 15045 6779 15079
rect 2053 14977 2087 15011
rect 3617 14977 3651 15011
rect 3985 14977 4019 15011
rect 4445 14977 4479 15011
rect 4537 14977 4571 15011
rect 4721 14977 4755 15011
rect 5917 14977 5951 15011
rect 7481 14977 7515 15011
rect 7757 14977 7791 15011
rect 8493 14977 8527 15011
rect 8585 14977 8619 15011
rect 9229 14977 9263 15011
rect 9413 14977 9447 15011
rect 3433 14909 3467 14943
rect 5825 14909 5859 14943
rect 9413 14841 9447 14875
rect 2237 14773 2271 14807
rect 4905 14773 4939 14807
rect 5549 14773 5583 14807
rect 5825 14773 5859 14807
rect 6745 14773 6779 14807
rect 7573 14773 7607 14807
rect 8585 14773 8619 14807
rect 2973 14569 3007 14603
rect 4353 14569 4387 14603
rect 10057 14501 10091 14535
rect 3157 14433 3191 14467
rect 5549 14433 5583 14467
rect 6285 14433 6319 14467
rect 1869 14365 1903 14399
rect 2145 14365 2179 14399
rect 3341 14365 3375 14399
rect 3433 14365 3467 14399
rect 4537 14365 4571 14399
rect 4721 14365 4755 14399
rect 4813 14365 4847 14399
rect 5733 14365 5767 14399
rect 5825 14365 5859 14399
rect 6469 14365 6503 14399
rect 6837 14365 6871 14399
rect 7849 14365 7883 14399
rect 8033 14365 8067 14399
rect 9137 14365 9171 14399
rect 9229 14365 9263 14399
rect 9413 14365 9447 14399
rect 10149 14365 10183 14399
rect 10793 14365 10827 14399
rect 10977 14365 11011 14399
rect 13277 14365 13311 14399
rect 13461 14365 13495 14399
rect 2329 14297 2363 14331
rect 10701 14297 10735 14331
rect 1961 14229 1995 14263
rect 5365 14229 5399 14263
rect 6745 14229 6779 14263
rect 7941 14229 7975 14263
rect 13461 14229 13495 14263
rect 4261 14025 4295 14059
rect 5273 14025 5307 14059
rect 7941 14025 7975 14059
rect 2145 13957 2179 13991
rect 3249 13957 3283 13991
rect 8493 13957 8527 13991
rect 12081 13957 12115 13991
rect 12541 13957 12575 13991
rect 12725 13957 12759 13991
rect 13461 13957 13495 13991
rect 14473 13957 14507 13991
rect 1909 13889 1943 13923
rect 2053 13889 2087 13923
rect 2329 13889 2363 13923
rect 3013 13889 3047 13923
rect 3157 13889 3191 13923
rect 3433 13889 3467 13923
rect 5089 13889 5123 13923
rect 6653 13889 6687 13923
rect 7021 13889 7055 13923
rect 7757 13889 7791 13923
rect 8677 13889 8711 13923
rect 9321 13889 9355 13923
rect 9505 13889 9539 13923
rect 10241 13889 10275 13923
rect 10333 13889 10367 13923
rect 11897 13889 11931 13923
rect 12909 13889 12943 13923
rect 13645 13889 13679 13923
rect 13737 13889 13771 13923
rect 14657 13889 14691 13923
rect 4077 13821 4111 13855
rect 4445 13821 4479 13855
rect 5457 13821 5491 13855
rect 7573 13821 7607 13855
rect 14289 13821 14323 13855
rect 8861 13753 8895 13787
rect 9597 13753 9631 13787
rect 10425 13753 10459 13787
rect 1777 13685 1811 13719
rect 2881 13685 2915 13719
rect 4629 13685 4663 13719
rect 5641 13685 5675 13719
rect 6929 13685 6963 13719
rect 11805 13685 11839 13719
rect 4077 13481 4111 13515
rect 6101 13481 6135 13515
rect 7481 13481 7515 13515
rect 12725 13481 12759 13515
rect 1593 13413 1627 13447
rect 5365 13413 5399 13447
rect 8217 13413 8251 13447
rect 6285 13345 6319 13379
rect 12173 13345 12207 13379
rect 1777 13277 1811 13311
rect 2421 13277 2455 13311
rect 2697 13277 2731 13311
rect 2841 13277 2875 13311
rect 4261 13277 4295 13311
rect 4353 13277 4387 13311
rect 4445 13277 4479 13311
rect 4537 13277 4571 13311
rect 5181 13277 5215 13311
rect 5457 13277 5491 13311
rect 6009 13277 6043 13311
rect 6929 13277 6963 13311
rect 7297 13277 7331 13311
rect 8309 13277 8343 13311
rect 8493 13277 8527 13311
rect 9597 13277 9631 13311
rect 9781 13277 9815 13311
rect 10149 13277 10183 13311
rect 10885 13277 10919 13311
rect 11069 13277 11103 13311
rect 11621 13277 11655 13311
rect 11989 13277 12023 13311
rect 12817 13277 12851 13311
rect 14381 13277 14415 13311
rect 14565 13277 14599 13311
rect 16405 13277 16439 13311
rect 16589 13277 16623 13311
rect 1961 13209 1995 13243
rect 2605 13209 2639 13243
rect 7941 13209 7975 13243
rect 13001 13209 13035 13243
rect 14657 13209 14691 13243
rect 2990 13141 3024 13175
rect 7113 13141 7147 13175
rect 10057 13141 10091 13175
rect 10701 13141 10735 13175
rect 11989 13141 12023 13175
rect 16405 13141 16439 13175
rect 2329 12937 2363 12971
rect 2421 12937 2455 12971
rect 10977 12937 11011 12971
rect 16221 12937 16255 12971
rect 4077 12869 4111 12903
rect 5181 12869 5215 12903
rect 7665 12869 7699 12903
rect 7757 12869 7791 12903
rect 13277 12869 13311 12903
rect 1961 12801 1995 12835
rect 3847 12801 3881 12835
rect 3985 12801 4019 12835
rect 4260 12801 4294 12835
rect 4353 12801 4387 12835
rect 5549 12801 5583 12835
rect 5641 12801 5675 12835
rect 5825 12801 5859 12835
rect 6653 12801 6687 12835
rect 6837 12801 6871 12835
rect 6929 12801 6963 12835
rect 7941 12801 7975 12835
rect 9229 12801 9263 12835
rect 10793 12801 10827 12835
rect 11069 12801 11103 12835
rect 11805 12801 11839 12835
rect 14289 12801 14323 12835
rect 14565 12801 14599 12835
rect 15209 12801 15243 12835
rect 15393 12801 15427 12835
rect 16037 12801 16071 12835
rect 16221 12801 16255 12835
rect 16957 12801 16991 12835
rect 17141 12801 17175 12835
rect 5457 12767 5491 12801
rect 2220 12733 2254 12767
rect 2513 12733 2547 12767
rect 5365 12733 5399 12767
rect 7205 12733 7239 12767
rect 9413 12733 9447 12767
rect 10057 12733 10091 12767
rect 10609 12733 10643 12767
rect 12725 12733 12759 12767
rect 3709 12665 3743 12699
rect 13553 12665 13587 12699
rect 15209 12665 15243 12699
rect 16957 12665 16991 12699
rect 1961 12597 1995 12631
rect 7113 12597 7147 12631
rect 8125 12597 8159 12631
rect 13737 12597 13771 12631
rect 14381 12597 14415 12631
rect 4261 12393 4295 12427
rect 6561 12393 6595 12427
rect 9321 12393 9355 12427
rect 10609 12393 10643 12427
rect 1869 12325 1903 12359
rect 4629 12325 4663 12359
rect 7665 12325 7699 12359
rect 14289 12325 14323 12359
rect 2125 12257 2159 12291
rect 2329 12257 2363 12291
rect 2973 12257 3007 12291
rect 7573 12257 7607 12291
rect 8125 12257 8159 12291
rect 9873 12257 9907 12291
rect 1869 12189 1903 12223
rect 2421 12189 2455 12223
rect 3157 12189 3191 12223
rect 3341 12189 3375 12223
rect 3433 12189 3467 12223
rect 4445 12189 4479 12223
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 5457 12189 5491 12223
rect 5549 12189 5583 12223
rect 6693 12189 6727 12223
rect 6837 12189 6871 12223
rect 7113 12189 7147 12223
rect 7941 12189 7975 12223
rect 9577 12189 9611 12223
rect 10333 12189 10367 12223
rect 11529 12189 11563 12223
rect 11621 12189 11655 12223
rect 12449 12189 12483 12223
rect 12725 12189 12759 12223
rect 14473 12189 14507 12223
rect 15209 12189 15243 12223
rect 15301 12189 15335 12223
rect 16129 12189 16163 12223
rect 16313 12189 16347 12223
rect 16957 12189 16991 12223
rect 17141 12189 17175 12223
rect 5273 12121 5307 12155
rect 5641 12121 5675 12155
rect 6929 12121 6963 12155
rect 9321 12121 9355 12155
rect 10977 12121 11011 12155
rect 14657 12121 14691 12155
rect 15485 12121 15519 12155
rect 16865 12121 16899 12155
rect 17693 12121 17727 12155
rect 17877 12121 17911 12155
rect 18061 12121 18095 12155
rect 2237 12053 2271 12087
rect 5825 12053 5859 12087
rect 9689 12053 9723 12087
rect 9781 12053 9815 12087
rect 10600 12053 10634 12087
rect 11805 12053 11839 12087
rect 13461 12053 13495 12087
rect 16129 12053 16163 12087
rect 2329 11849 2363 11883
rect 2697 11849 2731 11883
rect 5181 11849 5215 11883
rect 13737 11849 13771 11883
rect 2513 11781 2547 11815
rect 2605 11781 2639 11815
rect 2881 11781 2915 11815
rect 8401 11781 8435 11815
rect 10425 11781 10459 11815
rect 12449 11781 12483 11815
rect 13645 11781 13679 11815
rect 17969 11781 18003 11815
rect 3985 11713 4019 11747
rect 4143 11713 4177 11747
rect 4353 11713 4387 11747
rect 4629 11713 4663 11747
rect 5365 11713 5399 11747
rect 5641 11713 5675 11747
rect 5825 11713 5859 11747
rect 6561 11713 6595 11747
rect 6837 11713 6871 11747
rect 7113 11713 7147 11747
rect 8033 11713 8067 11747
rect 8953 11713 8987 11747
rect 9505 11713 9539 11747
rect 10241 11713 10275 11747
rect 10517 11713 10551 11747
rect 10661 11713 10695 11747
rect 12173 11713 12207 11747
rect 12266 11713 12300 11747
rect 12541 11713 12575 11747
rect 12679 11713 12713 11747
rect 14749 11713 14783 11747
rect 14933 11713 14967 11747
rect 15485 11713 15519 11747
rect 15669 11713 15703 11747
rect 16957 11713 16991 11747
rect 17141 11713 17175 11747
rect 18153 11713 18187 11747
rect 5457 11645 5491 11679
rect 6653 11645 6687 11679
rect 8125 11645 8159 11679
rect 8309 11645 8343 11679
rect 8493 11645 8527 11679
rect 9321 11645 9355 11679
rect 9781 11645 9815 11679
rect 13461 11645 13495 11679
rect 16865 11645 16899 11679
rect 5549 11577 5583 11611
rect 9045 11577 9079 11611
rect 14657 11577 14691 11611
rect 15485 11577 15519 11611
rect 17785 11577 17819 11611
rect 4353 11509 4387 11543
rect 7849 11509 7883 11543
rect 10793 11509 10827 11543
rect 12817 11509 12851 11543
rect 14105 11509 14139 11543
rect 11897 11305 11931 11339
rect 14289 11305 14323 11339
rect 3985 11237 4019 11271
rect 5181 11237 5215 11271
rect 5917 11237 5951 11271
rect 6469 11237 6503 11271
rect 10793 11237 10827 11271
rect 10885 11237 10919 11271
rect 14657 11237 14691 11271
rect 2493 11169 2527 11203
rect 2789 11169 2823 11203
rect 4629 11169 4663 11203
rect 8125 11169 8159 11203
rect 9965 11169 9999 11203
rect 10425 11169 10459 11203
rect 15209 11169 15243 11203
rect 2053 11101 2087 11135
rect 4353 11101 4387 11135
rect 4445 11101 4479 11135
rect 5181 11101 5215 11135
rect 6101 11101 6135 11135
rect 6469 11101 6503 11135
rect 7941 11101 7975 11135
rect 9229 11101 9263 11135
rect 9781 11101 9815 11135
rect 11529 11101 11563 11135
rect 11989 11101 12023 11135
rect 12725 11101 12759 11135
rect 12909 11101 12943 11135
rect 14289 11101 14323 11135
rect 14381 11101 14415 11135
rect 15301 11101 15335 11135
rect 15485 11101 15519 11135
rect 16405 11101 16439 11135
rect 16681 11101 16715 11135
rect 17325 11101 17359 11135
rect 17509 11101 17543 11135
rect 2237 11033 2271 11067
rect 2697 11033 2731 11067
rect 6745 11033 6779 11067
rect 9413 11033 9447 11067
rect 16773 11033 16807 11067
rect 17233 11033 17267 11067
rect 2605 10965 2639 10999
rect 7205 10965 7239 10999
rect 9321 10965 9355 10999
rect 13737 10965 13771 10999
rect 2973 10761 3007 10795
rect 3065 10761 3099 10795
rect 4169 10761 4203 10795
rect 5457 10761 5491 10795
rect 8861 10761 8895 10795
rect 14841 10761 14875 10795
rect 17969 10761 18003 10795
rect 2605 10693 2639 10727
rect 5365 10693 5399 10727
rect 10977 10693 11011 10727
rect 1777 10625 1811 10659
rect 1961 10625 1995 10659
rect 2835 10625 2869 10659
rect 3709 10625 3743 10659
rect 3985 10625 4019 10659
rect 5273 10625 5307 10659
rect 5825 10625 5859 10659
rect 12323 10625 12357 10659
rect 12725 10625 12759 10659
rect 13461 10625 13495 10659
rect 14933 10625 14967 10659
rect 15117 10625 15151 10659
rect 15669 10625 15703 10659
rect 15853 10625 15887 10659
rect 17969 10625 18003 10659
rect 3157 10557 3191 10591
rect 4261 10557 4295 10591
rect 5565 10557 5599 10591
rect 7120 10557 7154 10591
rect 10149 10557 10183 10591
rect 12633 10557 12667 10591
rect 13369 10557 13403 10591
rect 14289 10557 14323 10591
rect 17601 10557 17635 10591
rect 18153 10557 18187 10591
rect 1869 10489 1903 10523
rect 12081 10489 12115 10523
rect 15669 10489 15703 10523
rect 2421 10421 2455 10455
rect 3893 10421 3927 10455
rect 4445 10421 4479 10455
rect 6009 10421 6043 10455
rect 7376 10421 7410 10455
rect 10149 10149 10183 10183
rect 7757 10081 7791 10115
rect 15761 10081 15795 10115
rect 18107 10081 18141 10115
rect 1593 10013 1627 10047
rect 2145 10013 2179 10047
rect 3249 10013 3283 10047
rect 4077 10013 4111 10047
rect 5549 10013 5583 10047
rect 6377 10013 6411 10047
rect 7297 10013 7331 10047
rect 9321 10013 9355 10047
rect 9781 10013 9815 10047
rect 10701 10013 10735 10047
rect 12725 10013 12759 10047
rect 13093 10013 13127 10047
rect 14289 10013 14323 10047
rect 14473 10013 14507 10047
rect 14657 10013 14691 10047
rect 15485 10013 15519 10047
rect 17969 10013 18003 10047
rect 18337 10013 18371 10047
rect 1685 9945 1719 9979
rect 2697 9945 2731 9979
rect 2789 9945 2823 9979
rect 3985 9945 4019 9979
rect 6561 9945 6595 9979
rect 8217 9945 8251 9979
rect 8309 9945 8343 9979
rect 9137 9945 9171 9979
rect 9965 9945 9999 9979
rect 11713 9945 11747 9979
rect 7113 9877 7147 9911
rect 13737 9877 13771 9911
rect 17233 9877 17267 9911
rect 17969 9877 18003 9911
rect 5273 9673 5307 9707
rect 5365 9673 5399 9707
rect 12081 9673 12115 9707
rect 4169 9605 4203 9639
rect 4905 9605 4939 9639
rect 7021 9605 7055 9639
rect 8217 9605 8251 9639
rect 13461 9605 13495 9639
rect 17325 9605 17359 9639
rect 1685 9537 1719 9571
rect 1869 9537 1903 9571
rect 2329 9537 2363 9571
rect 3065 9537 3099 9571
rect 4077 9537 4111 9571
rect 5457 9537 5491 9571
rect 6561 9537 6595 9571
rect 7113 9537 7147 9571
rect 8953 9537 8987 9571
rect 9873 9537 9907 9571
rect 11989 9537 12023 9571
rect 14105 9537 14139 9571
rect 14315 9537 14349 9571
rect 15025 9537 15059 9571
rect 15117 9537 15151 9571
rect 15945 9537 15979 9571
rect 16129 9537 16163 9571
rect 17049 9537 17083 9571
rect 17877 9537 17911 9571
rect 18061 9537 18095 9571
rect 2973 9469 3007 9503
rect 3525 9469 3559 9503
rect 5164 9469 5198 9503
rect 7665 9469 7699 9503
rect 11897 9469 11931 9503
rect 14473 9469 14507 9503
rect 15853 9469 15887 9503
rect 16865 9469 16899 9503
rect 17417 9469 17451 9503
rect 2513 9401 2547 9435
rect 8125 9401 8159 9435
rect 10241 9401 10275 9435
rect 13001 9401 13035 9435
rect 13185 9401 13219 9435
rect 17969 9401 18003 9435
rect 4721 9333 4755 9367
rect 12449 9333 12483 9367
rect 14013 9333 14047 9367
rect 15301 9333 15335 9367
rect 17509 9129 17543 9163
rect 13369 9061 13403 9095
rect 9781 8993 9815 9027
rect 9873 8993 9907 9027
rect 11621 8993 11655 9027
rect 14289 8993 14323 9027
rect 18061 8993 18095 9027
rect 1593 8925 1627 8959
rect 2145 8925 2179 8959
rect 3249 8925 3283 8959
rect 4077 8925 4111 8959
rect 5549 8925 5583 8959
rect 6561 8925 6595 8959
rect 7297 8925 7331 8959
rect 7757 8925 7791 8959
rect 9321 8925 9355 8959
rect 10240 8925 10274 8959
rect 11161 8925 11195 8959
rect 16681 8925 16715 8959
rect 16865 8925 16899 8959
rect 17877 8925 17911 8959
rect 17969 8925 18003 8959
rect 1685 8857 1719 8891
rect 2697 8857 2731 8891
rect 2789 8857 2823 8891
rect 3985 8857 4019 8891
rect 6377 8857 6411 8891
rect 8217 8857 8251 8891
rect 8309 8857 8343 8891
rect 10425 8857 10459 8891
rect 11897 8857 11931 8891
rect 14565 8857 14599 8891
rect 7113 8789 7147 8823
rect 9229 8789 9263 8823
rect 10977 8789 11011 8823
rect 16037 8789 16071 8823
rect 16681 8789 16715 8823
rect 4169 8585 4203 8619
rect 5273 8585 5307 8619
rect 15025 8585 15059 8619
rect 16037 8585 16071 8619
rect 17877 8585 17911 8619
rect 18153 8585 18187 8619
rect 7021 8517 7055 8551
rect 8217 8517 8251 8551
rect 13553 8517 13587 8551
rect 17601 8517 17635 8551
rect 1685 8449 1719 8483
rect 1869 8449 1903 8483
rect 2329 8449 2363 8483
rect 3065 8449 3099 8483
rect 4077 8449 4111 8483
rect 4905 8449 4939 8483
rect 5135 8449 5169 8483
rect 5365 8449 5399 8483
rect 5457 8449 5491 8483
rect 6561 8449 6595 8483
rect 7113 8449 7147 8483
rect 7665 8449 7699 8483
rect 8953 8449 8987 8483
rect 9873 8449 9907 8483
rect 11713 8449 11747 8483
rect 12081 8449 12115 8483
rect 12173 8449 12207 8483
rect 15853 8449 15887 8483
rect 16129 8449 16163 8483
rect 17785 8449 17819 8483
rect 17969 8449 18003 8483
rect 2973 8381 3007 8415
rect 3525 8381 3559 8415
rect 11805 8381 11839 8415
rect 13277 8381 13311 8415
rect 2513 8313 2547 8347
rect 4721 8313 4755 8347
rect 8125 8313 8159 8347
rect 10241 8313 10275 8347
rect 15669 8313 15703 8347
rect 10057 8041 10091 8075
rect 13369 8041 13403 8075
rect 17325 8041 17359 8075
rect 10701 7973 10735 8007
rect 13001 7973 13035 8007
rect 14749 7973 14783 8007
rect 7757 7905 7791 7939
rect 12173 7905 12207 7939
rect 12449 7905 12483 7939
rect 15853 7905 15887 7939
rect 1593 7837 1627 7871
rect 2145 7837 2179 7871
rect 3249 7837 3283 7871
rect 4077 7837 4111 7871
rect 5549 7837 5583 7871
rect 6561 7837 6595 7871
rect 7297 7837 7331 7871
rect 9321 7837 9355 7871
rect 9781 7837 9815 7871
rect 12909 7837 12943 7871
rect 13185 7837 13219 7871
rect 14565 7837 14599 7871
rect 14841 7837 14875 7871
rect 15577 7837 15611 7871
rect 17877 7837 17911 7871
rect 18153 7837 18187 7871
rect 1685 7769 1719 7803
rect 2697 7769 2731 7803
rect 2789 7769 2823 7803
rect 3985 7769 4019 7803
rect 6377 7769 6411 7803
rect 8217 7769 8251 7803
rect 8309 7769 8343 7803
rect 9965 7769 9999 7803
rect 14381 7769 14415 7803
rect 7113 7701 7147 7735
rect 9229 7701 9263 7735
rect 17969 7701 18003 7735
rect 4169 7497 4203 7531
rect 5917 7497 5951 7531
rect 1685 7429 1719 7463
rect 3065 7429 3099 7463
rect 4077 7429 4111 7463
rect 7021 7429 7055 7463
rect 8217 7429 8251 7463
rect 17693 7429 17727 7463
rect 1869 7361 1903 7395
rect 2329 7361 2363 7395
rect 5273 7361 5307 7395
rect 6561 7361 6595 7395
rect 7113 7361 7147 7395
rect 7665 7361 7699 7395
rect 8953 7361 8987 7395
rect 9873 7361 9907 7395
rect 2973 7293 3007 7327
rect 3525 7293 3559 7327
rect 5457 7293 5491 7327
rect 5549 7293 5583 7327
rect 5641 7293 5675 7327
rect 5733 7293 5767 7327
rect 13737 7293 13771 7327
rect 14013 7293 14047 7327
rect 14473 7293 14507 7327
rect 14749 7293 14783 7327
rect 17785 7293 17819 7327
rect 17969 7293 18003 7327
rect 2513 7225 2547 7259
rect 8125 7225 8159 7259
rect 10241 7225 10275 7259
rect 12265 7225 12299 7259
rect 17325 7225 17359 7259
rect 16221 7157 16255 7191
rect 9873 6953 9907 6987
rect 11357 6953 11391 6987
rect 12725 6817 12759 6851
rect 14289 6817 14323 6851
rect 18337 6817 18371 6851
rect 1593 6749 1627 6783
rect 2145 6749 2179 6783
rect 3249 6749 3283 6783
rect 4077 6749 4111 6783
rect 5549 6749 5583 6783
rect 6561 6749 6595 6783
rect 7297 6749 7331 6783
rect 7757 6749 7791 6783
rect 9321 6749 9355 6783
rect 11621 6749 11655 6783
rect 12449 6749 12483 6783
rect 13369 6749 13403 6783
rect 13553 6749 13587 6783
rect 17509 6749 17543 6783
rect 17785 6749 17819 6783
rect 1685 6681 1719 6715
rect 2697 6681 2731 6715
rect 2789 6681 2823 6715
rect 3985 6681 4019 6715
rect 6377 6681 6411 6715
rect 8217 6681 8251 6715
rect 8309 6681 8343 6715
rect 13277 6681 13311 6715
rect 14565 6681 14599 6715
rect 7113 6613 7147 6647
rect 9229 6613 9263 6647
rect 12081 6613 12115 6647
rect 12541 6613 12575 6647
rect 16037 6613 16071 6647
rect 4169 6409 4203 6443
rect 5273 6341 5307 6375
rect 5917 6341 5951 6375
rect 7021 6341 7055 6375
rect 8217 6341 8251 6375
rect 13829 6341 13863 6375
rect 18337 6341 18371 6375
rect 1685 6273 1719 6307
rect 1869 6273 1903 6307
rect 2329 6273 2363 6307
rect 3065 6273 3099 6307
rect 4077 6273 4111 6307
rect 5457 6273 5491 6307
rect 5794 6273 5828 6307
rect 6561 6273 6595 6307
rect 7113 6273 7147 6307
rect 8953 6273 8987 6307
rect 9873 6273 9907 6307
rect 11161 6273 11195 6307
rect 14657 6273 14691 6307
rect 14841 6273 14875 6307
rect 15393 6273 15427 6307
rect 15761 6273 15795 6307
rect 15945 6273 15979 6307
rect 17325 6273 17359 6307
rect 2973 6205 3007 6239
rect 3525 6205 3559 6239
rect 5716 6205 5750 6239
rect 6009 6205 6043 6239
rect 7665 6205 7699 6239
rect 11069 6205 11103 6239
rect 12357 6205 12391 6239
rect 14105 6205 14139 6239
rect 15577 6205 15611 6239
rect 2513 6137 2547 6171
rect 8125 6137 8159 6171
rect 10241 6137 10275 6171
rect 14657 6137 14691 6171
rect 10333 5865 10367 5899
rect 14381 5865 14415 5899
rect 17049 5865 17083 5899
rect 2789 5797 2823 5831
rect 4077 5797 4111 5831
rect 18153 5797 18187 5831
rect 2697 5729 2731 5763
rect 7757 5729 7791 5763
rect 11805 5729 11839 5763
rect 13001 5729 13035 5763
rect 13185 5729 13219 5763
rect 14565 5729 14599 5763
rect 15301 5729 15335 5763
rect 15577 5729 15611 5763
rect 1593 5661 1627 5695
rect 2145 5661 2179 5695
rect 3249 5661 3283 5695
rect 4077 5661 4111 5695
rect 5549 5661 5583 5695
rect 6561 5661 6595 5695
rect 7297 5661 7331 5695
rect 9321 5661 9355 5695
rect 12081 5661 12115 5695
rect 14749 5661 14783 5695
rect 14841 5661 14875 5695
rect 17601 5661 17635 5695
rect 17831 5661 17865 5695
rect 1685 5593 1719 5627
rect 6377 5593 6411 5627
rect 8217 5593 8251 5627
rect 8309 5593 8343 5627
rect 9137 5593 9171 5627
rect 17969 5593 18003 5627
rect 7113 5525 7147 5559
rect 12541 5525 12575 5559
rect 12909 5525 12943 5559
rect 17785 5525 17819 5559
rect 4169 5321 4203 5355
rect 5641 5321 5675 5355
rect 5733 5321 5767 5355
rect 15761 5321 15795 5355
rect 3065 5253 3099 5287
rect 4077 5253 4111 5287
rect 7021 5253 7055 5287
rect 8217 5253 8251 5287
rect 11989 5253 12023 5287
rect 17877 5253 17911 5287
rect 18061 5253 18095 5287
rect 1685 5185 1719 5219
rect 1869 5185 1903 5219
rect 2329 5185 2363 5219
rect 3525 5185 3559 5219
rect 5273 5185 5307 5219
rect 5529 5185 5563 5219
rect 6561 5185 6595 5219
rect 7113 5185 7147 5219
rect 8953 5185 8987 5219
rect 9873 5185 9907 5219
rect 14013 5185 14047 5219
rect 16957 5185 16991 5219
rect 2973 5117 3007 5151
rect 5825 5117 5859 5151
rect 7665 5117 7699 5151
rect 11713 5117 11747 5151
rect 13461 5117 13495 5151
rect 14289 5117 14323 5151
rect 17233 5117 17267 5151
rect 2513 5049 2547 5083
rect 8125 5049 8159 5083
rect 10241 5049 10275 5083
rect 18245 5049 18279 5083
rect 5273 4981 5307 5015
rect 17049 4981 17083 5015
rect 18061 4981 18095 5015
rect 17141 4777 17175 4811
rect 12081 4709 12115 4743
rect 13369 4709 13403 4743
rect 14289 4709 14323 4743
rect 17785 4709 17819 4743
rect 1777 4641 1811 4675
rect 3249 4641 3283 4675
rect 7757 4641 7791 4675
rect 9229 4641 9263 4675
rect 11345 4641 11379 4675
rect 12725 4641 12759 4675
rect 15393 4641 15427 4675
rect 15669 4641 15703 4675
rect 18245 4641 18279 4675
rect 1593 4573 1627 4607
rect 2145 4573 2179 4607
rect 4077 4573 4111 4607
rect 5549 4573 5583 4607
rect 6561 4573 6595 4607
rect 7297 4573 7331 4607
rect 9321 4573 9355 4607
rect 11621 4573 11655 4607
rect 13553 4573 13587 4607
rect 13737 4573 13771 4607
rect 14564 4573 14598 4607
rect 14657 4573 14691 4607
rect 14749 4573 14783 4607
rect 14933 4573 14967 4607
rect 17693 4573 17727 4607
rect 18061 4573 18095 4607
rect 2697 4505 2731 4539
rect 2789 4505 2823 4539
rect 3985 4505 4019 4539
rect 6377 4505 6411 4539
rect 8217 4505 8251 4539
rect 8309 4505 8343 4539
rect 12541 4505 12575 4539
rect 7113 4437 7147 4471
rect 9873 4437 9907 4471
rect 12449 4437 12483 4471
rect 4169 4233 4203 4267
rect 12173 4233 12207 4267
rect 15301 4233 15335 4267
rect 1685 4165 1719 4199
rect 3065 4165 3099 4199
rect 4077 4165 4111 4199
rect 5181 4165 5215 4199
rect 7021 4165 7055 4199
rect 8217 4165 8251 4199
rect 1869 4097 1903 4131
rect 2329 4097 2363 4131
rect 3525 4097 3559 4131
rect 6561 4097 6595 4131
rect 7113 4097 7147 4131
rect 8953 4097 8987 4131
rect 9873 4097 9907 4131
rect 10977 4097 11011 4131
rect 11713 4097 11747 4131
rect 11897 4097 11931 4131
rect 13553 4097 13587 4131
rect 14013 4097 14047 4131
rect 17141 4097 17175 4131
rect 17325 4097 17359 4131
rect 18153 4097 18187 4131
rect 2973 4029 3007 4063
rect 5733 4029 5767 4063
rect 7665 4029 7699 4063
rect 12265 4029 12299 4063
rect 13277 4029 13311 4063
rect 15393 4029 15427 4063
rect 15577 4029 15611 4063
rect 2513 3961 2547 3995
rect 8125 3961 8159 3995
rect 10241 3961 10275 3995
rect 11069 3893 11103 3927
rect 14933 3893 14967 3927
rect 8309 3689 8343 3723
rect 10701 3689 10735 3723
rect 2789 3621 2823 3655
rect 4261 3621 4295 3655
rect 7757 3621 7791 3655
rect 9229 3621 9263 3655
rect 9781 3621 9815 3655
rect 13645 3621 13679 3655
rect 11897 3553 11931 3587
rect 17141 3553 17175 3587
rect 17785 3553 17819 3587
rect 17969 3553 18003 3587
rect 1593 3485 1627 3519
rect 2145 3485 2179 3519
rect 3249 3485 3283 3519
rect 4077 3485 4111 3519
rect 5549 3485 5583 3519
rect 6009 3485 6043 3519
rect 8493 3485 8527 3519
rect 9137 3485 9171 3519
rect 9599 3485 9633 3519
rect 10609 3485 10643 3519
rect 10885 3485 10919 3519
rect 11161 3485 11195 3519
rect 11437 3485 11471 3519
rect 14473 3485 14507 3519
rect 15393 3485 15427 3519
rect 17693 3485 17727 3519
rect 18153 3485 18187 3519
rect 1685 3417 1719 3451
rect 2697 3417 2731 3451
rect 6285 3417 6319 3451
rect 12173 3417 12207 3451
rect 14289 3417 14323 3451
rect 14841 3417 14875 3451
rect 15669 3417 15703 3451
rect 9597 3349 9631 3383
rect 14565 3349 14599 3383
rect 14657 3349 14691 3383
rect 4077 3145 4111 3179
rect 7021 3145 7055 3179
rect 8033 3145 8067 3179
rect 8401 3145 8435 3179
rect 8493 3145 8527 3179
rect 9413 3145 9447 3179
rect 13277 3145 13311 3179
rect 13737 3145 13771 3179
rect 2421 3077 2455 3111
rect 3985 3077 4019 3111
rect 5733 3077 5767 3111
rect 7297 3077 7331 3111
rect 9597 3077 9631 3111
rect 14749 3077 14783 3111
rect 18245 3077 18279 3111
rect 1593 3009 1627 3043
rect 3341 3009 3375 3043
rect 5181 3009 5215 3043
rect 6745 3009 6779 3043
rect 7849 3009 7883 3043
rect 8585 3009 8619 3043
rect 10057 3009 10091 3043
rect 11069 3009 11103 3043
rect 12173 3009 12207 3043
rect 13645 3009 13679 3043
rect 14473 3009 14507 3043
rect 17325 3009 17359 3043
rect 18061 3009 18095 3043
rect 2329 2941 2363 2975
rect 2881 2941 2915 2975
rect 6653 2941 6687 2975
rect 12265 2941 12299 2975
rect 12725 2941 12759 2975
rect 13829 2941 13863 2975
rect 17049 2941 17083 2975
rect 17877 2941 17911 2975
rect 1777 2873 1811 2907
rect 9229 2873 9263 2907
rect 16957 2873 16991 2907
rect 3433 2805 3467 2839
rect 9413 2805 9447 2839
rect 16221 2805 16255 2839
rect 1593 2601 1627 2635
rect 3065 2601 3099 2635
rect 6745 2601 6779 2635
rect 6929 2601 6963 2635
rect 7757 2601 7791 2635
rect 10885 2601 10919 2635
rect 12909 2601 12943 2635
rect 14565 2601 14599 2635
rect 16055 2601 16089 2635
rect 1593 2465 1627 2499
rect 4169 2465 4203 2499
rect 8217 2465 8251 2499
rect 9321 2465 9355 2499
rect 9413 2465 9447 2499
rect 11897 2465 11931 2499
rect 13093 2465 13127 2499
rect 16313 2465 16347 2499
rect 17417 2465 17451 2499
rect 1961 2397 1995 2431
rect 3157 2397 3191 2431
rect 3341 2397 3375 2431
rect 5365 2397 5399 2431
rect 7757 2397 7791 2431
rect 8125 2397 8159 2431
rect 9137 2397 9171 2431
rect 9505 2397 9539 2431
rect 9597 2397 9631 2431
rect 10333 2397 10367 2431
rect 10753 2397 10787 2431
rect 11989 2397 12023 2431
rect 12357 2397 12391 2431
rect 13277 2397 13311 2431
rect 13369 2397 13403 2431
rect 16865 2397 16899 2431
rect 17049 2397 17083 2431
rect 17877 2397 17911 2431
rect 18061 2397 18095 2431
rect 4721 2329 4755 2363
rect 6561 2329 6595 2363
rect 9781 2329 9815 2363
rect 10517 2329 10551 2363
rect 10609 2329 10643 2363
rect 18245 2329 18279 2363
rect 6745 2261 6779 2295
rect 7573 2261 7607 2295
rect 12265 2261 12299 2295
rect 17049 2261 17083 2295
<< metal1 >>
rect 1578 17484 1584 17536
rect 1636 17524 1642 17536
rect 7926 17524 7932 17536
rect 1636 17496 7932 17524
rect 1636 17484 1642 17496
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 1104 17434 18860 17456
rect 1104 17382 5502 17434
rect 5554 17382 5566 17434
rect 5618 17382 5630 17434
rect 5682 17382 5694 17434
rect 5746 17382 5758 17434
rect 5810 17382 5822 17434
rect 5874 17382 5886 17434
rect 5938 17382 5950 17434
rect 6002 17382 6014 17434
rect 6066 17382 6078 17434
rect 6130 17382 6142 17434
rect 6194 17382 6206 17434
rect 6258 17382 6270 17434
rect 6322 17382 6334 17434
rect 6386 17382 6398 17434
rect 6450 17382 6462 17434
rect 6514 17382 6526 17434
rect 6578 17382 6590 17434
rect 6642 17382 6654 17434
rect 6706 17382 13502 17434
rect 13554 17382 13566 17434
rect 13618 17382 13630 17434
rect 13682 17382 13694 17434
rect 13746 17382 13758 17434
rect 13810 17382 13822 17434
rect 13874 17382 13886 17434
rect 13938 17382 13950 17434
rect 14002 17382 14014 17434
rect 14066 17382 14078 17434
rect 14130 17382 14142 17434
rect 14194 17382 14206 17434
rect 14258 17382 14270 17434
rect 14322 17382 14334 17434
rect 14386 17382 14398 17434
rect 14450 17382 14462 17434
rect 14514 17382 14526 17434
rect 14578 17382 14590 17434
rect 14642 17382 14654 17434
rect 14706 17382 18860 17434
rect 1104 17360 18860 17382
rect 2314 17280 2320 17332
rect 2372 17320 2378 17332
rect 4430 17320 4436 17332
rect 2372 17292 4436 17320
rect 2372 17280 2378 17292
rect 4430 17280 4436 17292
rect 4488 17280 4494 17332
rect 566 17212 572 17264
rect 624 17252 630 17264
rect 2409 17255 2467 17261
rect 2409 17252 2421 17255
rect 624 17224 2421 17252
rect 624 17212 630 17224
rect 2409 17221 2421 17224
rect 2455 17221 2467 17255
rect 2409 17215 2467 17221
rect 2593 17255 2651 17261
rect 2593 17221 2605 17255
rect 2639 17252 2651 17255
rect 4157 17255 4215 17261
rect 2639 17224 4108 17252
rect 2639 17221 2651 17224
rect 2593 17215 2651 17221
rect 14 17144 20 17196
rect 72 17184 78 17196
rect 3053 17187 3111 17193
rect 3053 17184 3065 17187
rect 72 17156 3065 17184
rect 72 17144 78 17156
rect 3053 17153 3065 17156
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 3326 17144 3332 17196
rect 3384 17144 3390 17196
rect 4080 17184 4108 17224
rect 4157 17221 4169 17255
rect 4203 17252 4215 17255
rect 7558 17252 7564 17264
rect 4203 17224 7564 17252
rect 4203 17221 4215 17224
rect 4157 17215 4215 17221
rect 7558 17212 7564 17224
rect 7616 17212 7622 17264
rect 4338 17184 4344 17196
rect 4080 17156 4344 17184
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 4890 17144 4896 17196
rect 4948 17144 4954 17196
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17184 5135 17187
rect 9030 17184 9036 17196
rect 5123 17156 9036 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 750 17076 756 17128
rect 808 17116 814 17128
rect 2038 17116 2044 17128
rect 808 17088 2044 17116
rect 808 17076 814 17088
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 3421 17119 3479 17125
rect 3421 17085 3433 17119
rect 3467 17116 3479 17119
rect 5092 17116 5120 17147
rect 9030 17144 9036 17156
rect 9088 17144 9094 17196
rect 3467 17088 5120 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 1210 17008 1216 17060
rect 1268 17048 1274 17060
rect 1946 17048 1952 17060
rect 1268 17020 1952 17048
rect 1268 17008 1274 17020
rect 1946 17008 1952 17020
rect 2004 17008 2010 17060
rect 2225 17051 2283 17057
rect 2225 17017 2237 17051
rect 2271 17048 2283 17051
rect 3234 17048 3240 17060
rect 2271 17020 3240 17048
rect 2271 17017 2283 17020
rect 2225 17011 2283 17017
rect 3234 17008 3240 17020
rect 3292 17008 3298 17060
rect 3878 17008 3884 17060
rect 3936 17048 3942 17060
rect 3973 17051 4031 17057
rect 3973 17048 3985 17051
rect 3936 17020 3985 17048
rect 3936 17008 3942 17020
rect 3973 17017 3985 17020
rect 4019 17017 4031 17051
rect 3973 17011 4031 17017
rect 5077 17051 5135 17057
rect 5077 17017 5089 17051
rect 5123 17048 5135 17051
rect 11146 17048 11152 17060
rect 5123 17020 11152 17048
rect 5123 17017 5135 17020
rect 5077 17011 5135 17017
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 1302 16940 1308 16992
rect 1360 16980 1366 16992
rect 1762 16980 1768 16992
rect 1360 16952 1768 16980
rect 1360 16940 1366 16952
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 2409 16983 2467 16989
rect 2409 16949 2421 16983
rect 2455 16980 2467 16983
rect 4522 16980 4528 16992
rect 2455 16952 4528 16980
rect 2455 16949 2467 16952
rect 2409 16943 2467 16949
rect 4522 16940 4528 16952
rect 4580 16940 4586 16992
rect 1104 16890 18860 16912
rect 1104 16838 1502 16890
rect 1554 16838 1566 16890
rect 1618 16838 1630 16890
rect 1682 16838 1694 16890
rect 1746 16838 1758 16890
rect 1810 16838 1822 16890
rect 1874 16838 1886 16890
rect 1938 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 2270 16890
rect 2322 16838 2334 16890
rect 2386 16838 2398 16890
rect 2450 16838 2462 16890
rect 2514 16838 2526 16890
rect 2578 16838 2590 16890
rect 2642 16838 2654 16890
rect 2706 16838 9502 16890
rect 9554 16838 9566 16890
rect 9618 16838 9630 16890
rect 9682 16838 9694 16890
rect 9746 16838 9758 16890
rect 9810 16838 9822 16890
rect 9874 16838 9886 16890
rect 9938 16838 9950 16890
rect 10002 16838 10014 16890
rect 10066 16838 10078 16890
rect 10130 16838 10142 16890
rect 10194 16838 10206 16890
rect 10258 16838 10270 16890
rect 10322 16838 10334 16890
rect 10386 16838 10398 16890
rect 10450 16838 10462 16890
rect 10514 16838 10526 16890
rect 10578 16838 10590 16890
rect 10642 16838 10654 16890
rect 10706 16838 17502 16890
rect 17554 16838 17566 16890
rect 17618 16838 17630 16890
rect 17682 16838 17694 16890
rect 17746 16838 17758 16890
rect 17810 16838 17822 16890
rect 17874 16838 17886 16890
rect 17938 16838 17950 16890
rect 18002 16838 18014 16890
rect 18066 16838 18078 16890
rect 18130 16838 18142 16890
rect 18194 16838 18206 16890
rect 18258 16838 18270 16890
rect 18322 16838 18334 16890
rect 18386 16838 18398 16890
rect 18450 16838 18462 16890
rect 18514 16838 18526 16890
rect 18578 16838 18590 16890
rect 18642 16838 18654 16890
rect 18706 16838 18860 16890
rect 1104 16816 18860 16838
rect 6365 16711 6423 16717
rect 6365 16677 6377 16711
rect 6411 16708 6423 16711
rect 8478 16708 8484 16720
rect 6411 16680 8484 16708
rect 6411 16677 6423 16680
rect 6365 16671 6423 16677
rect 8478 16668 8484 16680
rect 8536 16668 8542 16720
rect 934 16532 940 16584
rect 992 16572 998 16584
rect 1581 16575 1639 16581
rect 1581 16572 1593 16575
rect 992 16544 1593 16572
rect 992 16532 998 16544
rect 1581 16541 1593 16544
rect 1627 16541 1639 16575
rect 1581 16535 1639 16541
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16541 1915 16575
rect 1857 16535 1915 16541
rect 2685 16575 2743 16581
rect 2685 16541 2697 16575
rect 2731 16572 2743 16575
rect 2774 16572 2780 16584
rect 2731 16544 2780 16572
rect 2731 16541 2743 16544
rect 2685 16535 2743 16541
rect 1872 16436 1900 16535
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16572 4215 16575
rect 4798 16572 4804 16584
rect 4203 16544 4804 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 5350 16532 5356 16584
rect 5408 16532 5414 16584
rect 5442 16532 5448 16584
rect 5500 16532 5506 16584
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16541 6331 16575
rect 6273 16535 6331 16541
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16572 6515 16575
rect 6730 16572 6736 16584
rect 6503 16544 6736 16572
rect 6503 16541 6515 16544
rect 6457 16535 6515 16541
rect 1946 16464 1952 16516
rect 2004 16464 2010 16516
rect 2409 16507 2467 16513
rect 2409 16473 2421 16507
rect 2455 16504 2467 16507
rect 2869 16507 2927 16513
rect 2455 16476 2825 16504
rect 2455 16473 2467 16476
rect 2409 16467 2467 16473
rect 2498 16436 2504 16448
rect 1872 16408 2504 16436
rect 2498 16396 2504 16408
rect 2556 16396 2562 16448
rect 2797 16436 2825 16476
rect 2869 16473 2881 16507
rect 2915 16504 2927 16507
rect 3602 16504 3608 16516
rect 2915 16476 3608 16504
rect 2915 16473 2927 16476
rect 2869 16467 2927 16473
rect 3602 16464 3608 16476
rect 3660 16464 3666 16516
rect 3970 16464 3976 16516
rect 4028 16464 4034 16516
rect 4338 16464 4344 16516
rect 4396 16504 4402 16516
rect 4982 16504 4988 16516
rect 4396 16476 4988 16504
rect 4396 16464 4402 16476
rect 4982 16464 4988 16476
rect 5040 16464 5046 16516
rect 6288 16504 6316 16535
rect 6730 16532 6736 16544
rect 6788 16532 6794 16584
rect 7374 16504 7380 16516
rect 6288 16476 7380 16504
rect 7374 16464 7380 16476
rect 7432 16464 7438 16516
rect 2958 16436 2964 16448
rect 2797 16408 2964 16436
rect 2958 16396 2964 16408
rect 3016 16396 3022 16448
rect 5537 16439 5595 16445
rect 5537 16405 5549 16439
rect 5583 16436 5595 16439
rect 12250 16436 12256 16448
rect 5583 16408 12256 16436
rect 5583 16405 5595 16408
rect 5537 16399 5595 16405
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 1104 16346 18860 16368
rect 1104 16294 5502 16346
rect 5554 16294 5566 16346
rect 5618 16294 5630 16346
rect 5682 16294 5694 16346
rect 5746 16294 5758 16346
rect 5810 16294 5822 16346
rect 5874 16294 5886 16346
rect 5938 16294 5950 16346
rect 6002 16294 6014 16346
rect 6066 16294 6078 16346
rect 6130 16294 6142 16346
rect 6194 16294 6206 16346
rect 6258 16294 6270 16346
rect 6322 16294 6334 16346
rect 6386 16294 6398 16346
rect 6450 16294 6462 16346
rect 6514 16294 6526 16346
rect 6578 16294 6590 16346
rect 6642 16294 6654 16346
rect 6706 16294 13502 16346
rect 13554 16294 13566 16346
rect 13618 16294 13630 16346
rect 13682 16294 13694 16346
rect 13746 16294 13758 16346
rect 13810 16294 13822 16346
rect 13874 16294 13886 16346
rect 13938 16294 13950 16346
rect 14002 16294 14014 16346
rect 14066 16294 14078 16346
rect 14130 16294 14142 16346
rect 14194 16294 14206 16346
rect 14258 16294 14270 16346
rect 14322 16294 14334 16346
rect 14386 16294 14398 16346
rect 14450 16294 14462 16346
rect 14514 16294 14526 16346
rect 14578 16294 14590 16346
rect 14642 16294 14654 16346
rect 14706 16294 18860 16346
rect 1104 16272 18860 16294
rect 2225 16167 2283 16173
rect 2225 16133 2237 16167
rect 2271 16164 2283 16167
rect 2498 16164 2504 16176
rect 2271 16136 2504 16164
rect 2271 16133 2283 16136
rect 2225 16127 2283 16133
rect 2498 16124 2504 16136
rect 2556 16164 2562 16176
rect 4433 16167 4491 16173
rect 2556 16136 3464 16164
rect 2556 16124 2562 16136
rect 3436 16108 3464 16136
rect 4433 16133 4445 16167
rect 4479 16133 4491 16167
rect 4433 16127 4491 16133
rect 382 16056 388 16108
rect 440 16096 446 16108
rect 2133 16099 2191 16105
rect 2133 16096 2145 16099
rect 440 16068 2145 16096
rect 440 16056 446 16068
rect 2133 16065 2145 16068
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 3050 16096 3056 16108
rect 2455 16068 3056 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 3050 16056 3056 16068
rect 3108 16056 3114 16108
rect 3418 16056 3424 16108
rect 3476 16056 3482 16108
rect 3510 16056 3516 16108
rect 3568 16056 3574 16108
rect 3694 16056 3700 16108
rect 3752 16096 3758 16108
rect 4448 16096 4476 16127
rect 4614 16124 4620 16176
rect 4672 16124 4678 16176
rect 5629 16167 5687 16173
rect 5629 16133 5641 16167
rect 5675 16164 5687 16167
rect 6270 16164 6276 16176
rect 5675 16136 6276 16164
rect 5675 16133 5687 16136
rect 5629 16127 5687 16133
rect 6270 16124 6276 16136
rect 6328 16124 6334 16176
rect 6733 16167 6791 16173
rect 6733 16133 6745 16167
rect 6779 16164 6791 16167
rect 9214 16164 9220 16176
rect 6779 16136 9220 16164
rect 6779 16133 6791 16136
rect 6733 16127 6791 16133
rect 9214 16124 9220 16136
rect 9272 16124 9278 16176
rect 3752 16068 4476 16096
rect 5813 16099 5871 16105
rect 3752 16056 3758 16068
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6822 16096 6828 16108
rect 5859 16068 6828 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 6917 16099 6975 16105
rect 6917 16065 6929 16099
rect 6963 16065 6975 16099
rect 6917 16059 6975 16065
rect 474 15988 480 16040
rect 532 16028 538 16040
rect 5258 16028 5264 16040
rect 532 16000 5264 16028
rect 532 15988 538 16000
rect 5258 15988 5264 16000
rect 5316 15988 5322 16040
rect 6932 16028 6960 16059
rect 7466 16056 7472 16108
rect 7524 16056 7530 16108
rect 7650 16056 7656 16108
rect 7708 16056 7714 16108
rect 9122 16028 9128 16040
rect 6932 16000 9128 16028
rect 9122 15988 9128 16000
rect 9180 15988 9186 16040
rect 1946 15920 1952 15972
rect 2004 15960 2010 15972
rect 2682 15960 2688 15972
rect 2004 15932 2688 15960
rect 2004 15920 2010 15932
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 3326 15920 3332 15972
rect 3384 15960 3390 15972
rect 3881 15963 3939 15969
rect 3881 15960 3893 15963
rect 3384 15932 3893 15960
rect 3384 15920 3390 15932
rect 3881 15929 3893 15932
rect 3927 15929 3939 15963
rect 3881 15923 3939 15929
rect 7653 15963 7711 15969
rect 7653 15929 7665 15963
rect 7699 15960 7711 15963
rect 12342 15960 12348 15972
rect 7699 15932 12348 15960
rect 7699 15929 7711 15932
rect 7653 15923 7711 15929
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 2593 15895 2651 15901
rect 2593 15861 2605 15895
rect 2639 15892 2651 15895
rect 3142 15892 3148 15904
rect 2639 15864 3148 15892
rect 2639 15861 2651 15864
rect 2593 15855 2651 15861
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 4522 15852 4528 15904
rect 4580 15892 4586 15904
rect 4617 15895 4675 15901
rect 4617 15892 4629 15895
rect 4580 15864 4629 15892
rect 4580 15852 4586 15864
rect 4617 15861 4629 15864
rect 4663 15861 4675 15895
rect 4617 15855 4675 15861
rect 4706 15852 4712 15904
rect 4764 15892 4770 15904
rect 4801 15895 4859 15901
rect 4801 15892 4813 15895
rect 4764 15864 4813 15892
rect 4764 15852 4770 15864
rect 4801 15861 4813 15864
rect 4847 15861 4859 15895
rect 4801 15855 4859 15861
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5537 15895 5595 15901
rect 5537 15892 5549 15895
rect 5040 15864 5549 15892
rect 5040 15852 5046 15864
rect 5537 15861 5549 15864
rect 5583 15861 5595 15895
rect 5537 15855 5595 15861
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 6730 15892 6736 15904
rect 6687 15864 6736 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 6730 15852 6736 15864
rect 6788 15892 6794 15904
rect 6914 15892 6920 15904
rect 6788 15864 6920 15892
rect 6788 15852 6794 15864
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 1104 15802 18860 15824
rect 1104 15750 1502 15802
rect 1554 15750 1566 15802
rect 1618 15750 1630 15802
rect 1682 15750 1694 15802
rect 1746 15750 1758 15802
rect 1810 15750 1822 15802
rect 1874 15750 1886 15802
rect 1938 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 2270 15802
rect 2322 15750 2334 15802
rect 2386 15750 2398 15802
rect 2450 15750 2462 15802
rect 2514 15750 2526 15802
rect 2578 15750 2590 15802
rect 2642 15750 2654 15802
rect 2706 15750 9502 15802
rect 9554 15750 9566 15802
rect 9618 15750 9630 15802
rect 9682 15750 9694 15802
rect 9746 15750 9758 15802
rect 9810 15750 9822 15802
rect 9874 15750 9886 15802
rect 9938 15750 9950 15802
rect 10002 15750 10014 15802
rect 10066 15750 10078 15802
rect 10130 15750 10142 15802
rect 10194 15750 10206 15802
rect 10258 15750 10270 15802
rect 10322 15750 10334 15802
rect 10386 15750 10398 15802
rect 10450 15750 10462 15802
rect 10514 15750 10526 15802
rect 10578 15750 10590 15802
rect 10642 15750 10654 15802
rect 10706 15750 17502 15802
rect 17554 15750 17566 15802
rect 17618 15750 17630 15802
rect 17682 15750 17694 15802
rect 17746 15750 17758 15802
rect 17810 15750 17822 15802
rect 17874 15750 17886 15802
rect 17938 15750 17950 15802
rect 18002 15750 18014 15802
rect 18066 15750 18078 15802
rect 18130 15750 18142 15802
rect 18194 15750 18206 15802
rect 18258 15750 18270 15802
rect 18322 15750 18334 15802
rect 18386 15750 18398 15802
rect 18450 15750 18462 15802
rect 18514 15750 18526 15802
rect 18578 15750 18590 15802
rect 18642 15750 18654 15802
rect 18706 15750 18860 15802
rect 1104 15728 18860 15750
rect 2590 15648 2596 15700
rect 2648 15688 2654 15700
rect 2866 15688 2872 15700
rect 2648 15660 2872 15688
rect 2648 15648 2654 15660
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 3326 15688 3332 15700
rect 2976 15660 3332 15688
rect 1578 15580 1584 15632
rect 1636 15620 1642 15632
rect 2976 15620 3004 15660
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 5350 15648 5356 15700
rect 5408 15648 5414 15700
rect 6178 15648 6184 15700
rect 6236 15648 6242 15700
rect 6270 15648 6276 15700
rect 6328 15688 6334 15700
rect 8202 15688 8208 15700
rect 6328 15660 8208 15688
rect 6328 15648 6334 15660
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 1636 15592 3004 15620
rect 3053 15623 3111 15629
rect 1636 15580 1642 15592
rect 3053 15589 3065 15623
rect 3099 15620 3111 15623
rect 3786 15620 3792 15632
rect 3099 15592 3792 15620
rect 3099 15589 3111 15592
rect 3053 15583 3111 15589
rect 3786 15580 3792 15592
rect 3844 15580 3850 15632
rect 4890 15620 4896 15632
rect 4172 15592 4896 15620
rect 290 15512 296 15564
rect 348 15552 354 15564
rect 4172 15552 4200 15592
rect 4890 15580 4896 15592
rect 4948 15620 4954 15632
rect 8570 15620 8576 15632
rect 4948 15592 8576 15620
rect 4948 15580 4954 15592
rect 8570 15580 8576 15592
rect 8628 15580 8634 15632
rect 348 15524 4016 15552
rect 348 15512 354 15524
rect 474 15444 480 15496
rect 532 15484 538 15496
rect 658 15484 664 15496
rect 532 15456 664 15484
rect 532 15444 538 15456
rect 658 15444 664 15456
rect 716 15444 722 15496
rect 1946 15444 1952 15496
rect 2004 15444 2010 15496
rect 2682 15444 2688 15496
rect 2740 15444 2746 15496
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3988 15493 4016 15524
rect 4080 15524 4200 15552
rect 4433 15555 4491 15561
rect 4080 15496 4108 15524
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 7098 15552 7104 15564
rect 4479 15524 7104 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 7098 15512 7104 15524
rect 7156 15512 7162 15564
rect 8386 15512 8392 15564
rect 8444 15552 8450 15564
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 8444 15524 9137 15552
rect 8444 15512 8450 15524
rect 9125 15521 9137 15524
rect 9171 15521 9183 15555
rect 19058 15552 19064 15564
rect 9125 15515 9183 15521
rect 9324 15524 19064 15552
rect 3053 15487 3111 15493
rect 3053 15484 3065 15487
rect 3016 15456 3065 15484
rect 3016 15444 3022 15456
rect 3053 15453 3065 15456
rect 3099 15453 3111 15487
rect 3053 15447 3111 15453
rect 3237 15487 3295 15493
rect 3237 15453 3249 15487
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 198 15376 204 15428
rect 256 15416 262 15428
rect 1673 15419 1731 15425
rect 1673 15416 1685 15419
rect 256 15388 1685 15416
rect 256 15376 262 15388
rect 1673 15385 1685 15388
rect 1719 15385 1731 15419
rect 1673 15379 1731 15385
rect 2133 15419 2191 15425
rect 2133 15385 2145 15419
rect 2179 15385 2191 15419
rect 3252 15416 3280 15447
rect 4062 15444 4068 15496
rect 4120 15444 4126 15496
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4212 15456 4261 15484
rect 4212 15444 4218 15456
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15484 5687 15487
rect 7558 15484 7564 15496
rect 5675 15456 7564 15484
rect 5675 15453 5687 15456
rect 5629 15447 5687 15453
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 9324 15493 9352 15524
rect 19058 15512 19064 15524
rect 19116 15512 19122 15564
rect 9309 15487 9367 15493
rect 8036 15456 9260 15484
rect 3418 15416 3424 15428
rect 3252 15388 3424 15416
rect 2133 15379 2191 15385
rect 658 15308 664 15360
rect 716 15348 722 15360
rect 1026 15348 1032 15360
rect 716 15320 1032 15348
rect 716 15308 722 15320
rect 1026 15308 1032 15320
rect 1084 15308 1090 15360
rect 1765 15351 1823 15357
rect 1765 15317 1777 15351
rect 1811 15348 1823 15351
rect 1854 15348 1860 15360
rect 1811 15320 1860 15348
rect 1811 15317 1823 15320
rect 1765 15311 1823 15317
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 2148 15348 2176 15379
rect 3418 15376 3424 15388
rect 3476 15416 3482 15428
rect 4080 15416 4108 15444
rect 3476 15388 4108 15416
rect 3476 15376 3482 15388
rect 5166 15376 5172 15428
rect 5224 15376 5230 15428
rect 6270 15376 6276 15428
rect 6328 15376 6334 15428
rect 6457 15419 6515 15425
rect 6457 15385 6469 15419
rect 6503 15416 6515 15419
rect 6730 15416 6736 15428
rect 6503 15388 6736 15416
rect 6503 15385 6515 15388
rect 6457 15379 6515 15385
rect 6730 15376 6736 15388
rect 6788 15376 6794 15428
rect 6917 15419 6975 15425
rect 6917 15385 6929 15419
rect 6963 15416 6975 15419
rect 7006 15416 7012 15428
rect 6963 15388 7012 15416
rect 6963 15385 6975 15388
rect 6917 15379 6975 15385
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 7101 15419 7159 15425
rect 7101 15385 7113 15419
rect 7147 15385 7159 15419
rect 7101 15379 7159 15385
rect 3326 15348 3332 15360
rect 2148 15320 3332 15348
rect 3326 15308 3332 15320
rect 3384 15308 3390 15360
rect 3878 15308 3884 15360
rect 3936 15348 3942 15360
rect 4246 15348 4252 15360
rect 3936 15320 4252 15348
rect 3936 15308 3942 15320
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 4522 15308 4528 15360
rect 4580 15348 4586 15360
rect 4982 15348 4988 15360
rect 4580 15320 4988 15348
rect 4580 15308 4586 15320
rect 4982 15308 4988 15320
rect 5040 15348 5046 15360
rect 5353 15351 5411 15357
rect 5353 15348 5365 15351
rect 5040 15320 5365 15348
rect 5040 15308 5046 15320
rect 5353 15317 5365 15320
rect 5399 15317 5411 15351
rect 7116 15348 7144 15379
rect 7282 15376 7288 15428
rect 7340 15416 7346 15428
rect 8036 15416 8064 15456
rect 7340 15388 8064 15416
rect 7340 15376 7346 15388
rect 8110 15376 8116 15428
rect 8168 15376 8174 15428
rect 8202 15376 8208 15428
rect 8260 15416 8266 15428
rect 8297 15419 8355 15425
rect 8297 15416 8309 15419
rect 8260 15388 8309 15416
rect 8260 15376 8266 15388
rect 8297 15385 8309 15388
rect 8343 15385 8355 15419
rect 8297 15379 8355 15385
rect 8481 15419 8539 15425
rect 8481 15385 8493 15419
rect 8527 15416 8539 15419
rect 8570 15416 8576 15428
rect 8527 15388 8576 15416
rect 8527 15385 8539 15388
rect 8481 15379 8539 15385
rect 8570 15376 8576 15388
rect 8628 15376 8634 15428
rect 8018 15348 8024 15360
rect 7116 15320 8024 15348
rect 5353 15311 5411 15317
rect 8018 15308 8024 15320
rect 8076 15308 8082 15360
rect 9232 15348 9260 15456
rect 9309 15453 9321 15487
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 12802 15348 12808 15360
rect 9232 15320 12808 15348
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 290 15240 296 15292
rect 348 15280 354 15292
rect 750 15280 756 15292
rect 348 15252 756 15280
rect 348 15240 354 15252
rect 750 15240 756 15252
rect 808 15240 814 15292
rect 1104 15258 18860 15280
rect 1104 15206 5502 15258
rect 5554 15206 5566 15258
rect 5618 15206 5630 15258
rect 5682 15206 5694 15258
rect 5746 15206 5758 15258
rect 5810 15206 5822 15258
rect 5874 15206 5886 15258
rect 5938 15206 5950 15258
rect 6002 15206 6014 15258
rect 6066 15206 6078 15258
rect 6130 15206 6142 15258
rect 6194 15206 6206 15258
rect 6258 15206 6270 15258
rect 6322 15206 6334 15258
rect 6386 15206 6398 15258
rect 6450 15206 6462 15258
rect 6514 15206 6526 15258
rect 6578 15206 6590 15258
rect 6642 15206 6654 15258
rect 6706 15206 13502 15258
rect 13554 15206 13566 15258
rect 13618 15206 13630 15258
rect 13682 15206 13694 15258
rect 13746 15206 13758 15258
rect 13810 15206 13822 15258
rect 13874 15206 13886 15258
rect 13938 15206 13950 15258
rect 14002 15206 14014 15258
rect 14066 15206 14078 15258
rect 14130 15206 14142 15258
rect 14194 15206 14206 15258
rect 14258 15206 14270 15258
rect 14322 15206 14334 15258
rect 14386 15206 14398 15258
rect 14450 15206 14462 15258
rect 14514 15206 14526 15258
rect 14578 15206 14590 15258
rect 14642 15206 14654 15258
rect 14706 15206 18860 15258
rect 1104 15184 18860 15206
rect 1854 15104 1860 15156
rect 1912 15144 1918 15156
rect 3418 15144 3424 15156
rect 1912 15116 3424 15144
rect 1912 15104 1918 15116
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 3605 15147 3663 15153
rect 3605 15113 3617 15147
rect 3651 15144 3663 15147
rect 3694 15144 3700 15156
rect 3651 15116 3700 15144
rect 3651 15113 3663 15116
rect 3605 15107 3663 15113
rect 3694 15104 3700 15116
rect 3752 15104 3758 15156
rect 6917 15147 6975 15153
rect 6917 15144 6929 15147
rect 3896 15116 6929 15144
rect 1302 15036 1308 15088
rect 1360 15076 1366 15088
rect 1765 15079 1823 15085
rect 1765 15076 1777 15079
rect 1360 15048 1777 15076
rect 1360 15036 1366 15048
rect 1765 15045 1777 15048
rect 1811 15045 1823 15079
rect 1765 15039 1823 15045
rect 2866 15036 2872 15088
rect 2924 15076 2930 15088
rect 3896 15076 3924 15116
rect 6917 15113 6929 15116
rect 6963 15113 6975 15147
rect 6917 15107 6975 15113
rect 4062 15076 4068 15088
rect 2924 15048 3924 15076
rect 3988 15048 4068 15076
rect 2924 15036 2930 15048
rect 3988 15017 4016 15048
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 4338 15036 4344 15088
rect 4396 15076 4402 15088
rect 4396 15048 6040 15076
rect 4396 15036 4402 15048
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 3605 15011 3663 15017
rect 2087 14980 3556 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 750 14900 756 14952
rect 808 14940 814 14952
rect 1578 14940 1584 14952
rect 808 14912 1584 14940
rect 808 14900 814 14912
rect 1578 14900 1584 14912
rect 1636 14900 1642 14952
rect 2958 14900 2964 14952
rect 3016 14940 3022 14952
rect 3421 14943 3479 14949
rect 3421 14940 3433 14943
rect 3016 14912 3433 14940
rect 3016 14900 3022 14912
rect 3421 14909 3433 14912
rect 3467 14909 3479 14943
rect 3421 14903 3479 14909
rect 1302 14832 1308 14884
rect 1360 14872 1366 14884
rect 1946 14872 1952 14884
rect 1360 14844 1952 14872
rect 1360 14832 1366 14844
rect 1946 14832 1952 14844
rect 2004 14832 2010 14884
rect 1026 14764 1032 14816
rect 1084 14804 1090 14816
rect 2225 14807 2283 14813
rect 2225 14804 2237 14807
rect 1084 14776 2237 14804
rect 1084 14764 1090 14776
rect 2225 14773 2237 14776
rect 2271 14773 2283 14807
rect 3436 14804 3464 14903
rect 3528 14872 3556 14980
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 3973 15011 4031 15017
rect 3973 14977 3985 15011
rect 4019 14977 4031 15011
rect 3973 14971 4031 14977
rect 3620 14940 3648 14971
rect 4246 14968 4252 15020
rect 4304 15008 4310 15020
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 4304 14980 4445 15008
rect 4304 14968 4310 14980
rect 4433 14977 4445 14980
rect 4479 14977 4491 15011
rect 4433 14971 4491 14977
rect 4522 14968 4528 15020
rect 4580 14968 4586 15020
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 5074 15008 5080 15020
rect 4755 14980 5080 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 4062 14940 4068 14952
rect 3620 14912 4068 14940
rect 4062 14900 4068 14912
rect 4120 14940 4126 14952
rect 4724 14940 4752 14971
rect 5074 14968 5080 14980
rect 5132 14968 5138 15020
rect 5166 14968 5172 15020
rect 5224 15008 5230 15020
rect 5905 15011 5963 15017
rect 5905 15008 5917 15011
rect 5224 14980 5917 15008
rect 5224 14968 5230 14980
rect 5905 14977 5917 14980
rect 5951 14977 5963 15011
rect 6012 15008 6040 15048
rect 6546 15036 6552 15088
rect 6604 15036 6610 15088
rect 6733 15079 6791 15085
rect 6733 15045 6745 15079
rect 6779 15045 6791 15079
rect 6733 15039 6791 15045
rect 6748 15008 6776 15039
rect 7282 15036 7288 15088
rect 7340 15076 7346 15088
rect 8202 15076 8208 15088
rect 7340 15048 8208 15076
rect 7340 15036 7346 15048
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 8294 15036 8300 15088
rect 8352 15076 8358 15088
rect 14734 15076 14740 15088
rect 8352 15048 8616 15076
rect 8352 15036 8358 15048
rect 6012 14980 6776 15008
rect 7469 15011 7527 15017
rect 5905 14971 5963 14977
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 7650 15008 7656 15020
rect 7515 14980 7656 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 4120 14912 4752 14940
rect 4120 14900 4126 14912
rect 4798 14900 4804 14952
rect 4856 14940 4862 14952
rect 5813 14943 5871 14949
rect 5813 14940 5825 14943
rect 4856 14912 5825 14940
rect 4856 14900 4862 14912
rect 5813 14909 5825 14912
rect 5859 14940 5871 14943
rect 5994 14940 6000 14952
rect 5859 14912 6000 14940
rect 5859 14909 5871 14912
rect 5813 14903 5871 14909
rect 5994 14900 6000 14912
rect 6052 14940 6058 14952
rect 7760 14940 7788 14971
rect 8018 14968 8024 15020
rect 8076 15008 8082 15020
rect 8588 15017 8616 15048
rect 9232 15048 14740 15076
rect 9232 15020 9260 15048
rect 14734 15036 14740 15048
rect 14792 15036 14798 15088
rect 8481 15011 8539 15017
rect 8481 15008 8493 15011
rect 8076 14980 8493 15008
rect 8076 14968 8082 14980
rect 8481 14977 8493 14980
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 8573 15011 8631 15017
rect 8573 14977 8585 15011
rect 8619 14977 8631 15011
rect 8573 14971 8631 14977
rect 7834 14940 7840 14952
rect 6052 14912 7840 14940
rect 6052 14900 6058 14912
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 8496 14940 8524 14971
rect 9214 14968 9220 15020
rect 9272 14968 9278 15020
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 8846 14940 8852 14952
rect 8496 14912 8852 14940
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9416 14940 9444 14971
rect 9180 14912 9444 14940
rect 9180 14900 9186 14912
rect 4246 14872 4252 14884
rect 3528 14844 4252 14872
rect 4246 14832 4252 14844
rect 4304 14832 4310 14884
rect 8754 14872 8760 14884
rect 4356 14844 8760 14872
rect 4356 14804 4384 14844
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 9398 14832 9404 14884
rect 9456 14832 9462 14884
rect 3436 14776 4384 14804
rect 2225 14767 2283 14773
rect 4890 14764 4896 14816
rect 4948 14764 4954 14816
rect 5534 14764 5540 14816
rect 5592 14764 5598 14816
rect 5810 14764 5816 14816
rect 5868 14764 5874 14816
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 6733 14807 6791 14813
rect 6733 14804 6745 14807
rect 6696 14776 6745 14804
rect 6696 14764 6702 14776
rect 6733 14773 6745 14776
rect 6779 14773 6791 14807
rect 6733 14767 6791 14773
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 7561 14807 7619 14813
rect 7561 14804 7573 14807
rect 7524 14776 7573 14804
rect 7524 14764 7530 14776
rect 7561 14773 7573 14776
rect 7607 14804 7619 14807
rect 8294 14804 8300 14816
rect 7607 14776 8300 14804
rect 7607 14773 7619 14776
rect 7561 14767 7619 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 8573 14807 8631 14813
rect 8573 14773 8585 14807
rect 8619 14804 8631 14807
rect 8938 14804 8944 14816
rect 8619 14776 8944 14804
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 1104 14714 18860 14736
rect 1104 14662 1502 14714
rect 1554 14662 1566 14714
rect 1618 14662 1630 14714
rect 1682 14662 1694 14714
rect 1746 14662 1758 14714
rect 1810 14662 1822 14714
rect 1874 14662 1886 14714
rect 1938 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 2270 14714
rect 2322 14662 2334 14714
rect 2386 14662 2398 14714
rect 2450 14662 2462 14714
rect 2514 14662 2526 14714
rect 2578 14662 2590 14714
rect 2642 14662 2654 14714
rect 2706 14662 9502 14714
rect 9554 14662 9566 14714
rect 9618 14662 9630 14714
rect 9682 14662 9694 14714
rect 9746 14662 9758 14714
rect 9810 14662 9822 14714
rect 9874 14662 9886 14714
rect 9938 14662 9950 14714
rect 10002 14662 10014 14714
rect 10066 14662 10078 14714
rect 10130 14662 10142 14714
rect 10194 14662 10206 14714
rect 10258 14662 10270 14714
rect 10322 14662 10334 14714
rect 10386 14662 10398 14714
rect 10450 14662 10462 14714
rect 10514 14662 10526 14714
rect 10578 14662 10590 14714
rect 10642 14662 10654 14714
rect 10706 14662 17502 14714
rect 17554 14662 17566 14714
rect 17618 14662 17630 14714
rect 17682 14662 17694 14714
rect 17746 14662 17758 14714
rect 17810 14662 17822 14714
rect 17874 14662 17886 14714
rect 17938 14662 17950 14714
rect 18002 14662 18014 14714
rect 18066 14662 18078 14714
rect 18130 14662 18142 14714
rect 18194 14662 18206 14714
rect 18258 14662 18270 14714
rect 18322 14662 18334 14714
rect 18386 14662 18398 14714
rect 18450 14662 18462 14714
rect 18514 14662 18526 14714
rect 18578 14662 18590 14714
rect 18642 14662 18654 14714
rect 18706 14662 18860 14714
rect 1104 14640 18860 14662
rect 2130 14560 2136 14612
rect 2188 14600 2194 14612
rect 2961 14603 3019 14609
rect 2961 14600 2973 14603
rect 2188 14572 2973 14600
rect 2188 14560 2194 14572
rect 2961 14569 2973 14572
rect 3007 14569 3019 14603
rect 2961 14563 3019 14569
rect 4338 14560 4344 14612
rect 4396 14560 4402 14612
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 4580 14572 4936 14600
rect 4580 14560 4586 14572
rect 4154 14532 4160 14544
rect 3160 14504 4160 14532
rect 3160 14473 3188 14504
rect 4154 14492 4160 14504
rect 4212 14532 4218 14544
rect 4798 14532 4804 14544
rect 4212 14504 4804 14532
rect 4212 14492 4218 14504
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14433 3203 14467
rect 4908 14464 4936 14572
rect 5074 14560 5080 14612
rect 5132 14600 5138 14612
rect 8018 14600 8024 14612
rect 5132 14572 8024 14600
rect 5132 14560 5138 14572
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 4982 14492 4988 14544
rect 5040 14532 5046 14544
rect 5810 14532 5816 14544
rect 5040 14504 5816 14532
rect 5040 14492 5046 14504
rect 5810 14492 5816 14504
rect 5868 14532 5874 14544
rect 8662 14532 8668 14544
rect 5868 14504 8668 14532
rect 5868 14492 5874 14504
rect 8662 14492 8668 14504
rect 8720 14532 8726 14544
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 8720 14504 10057 14532
rect 8720 14492 8726 14504
rect 10045 14501 10057 14504
rect 10091 14501 10103 14535
rect 10045 14495 10103 14501
rect 3145 14427 3203 14433
rect 4724 14436 4936 14464
rect 1210 14356 1216 14408
rect 1268 14396 1274 14408
rect 1857 14399 1915 14405
rect 1857 14396 1869 14399
rect 1268 14368 1869 14396
rect 1268 14356 1274 14368
rect 1857 14365 1869 14368
rect 1903 14365 1915 14399
rect 1857 14359 1915 14365
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2222 14396 2228 14408
rect 2179 14368 2228 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 2958 14356 2964 14408
rect 3016 14396 3022 14408
rect 3329 14399 3387 14405
rect 3329 14396 3341 14399
rect 3016 14368 3341 14396
rect 3016 14356 3022 14368
rect 3329 14365 3341 14368
rect 3375 14365 3387 14399
rect 3329 14359 3387 14365
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 3694 14396 3700 14408
rect 3467 14368 3700 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 750 14288 756 14340
rect 808 14328 814 14340
rect 2317 14331 2375 14337
rect 2317 14328 2329 14331
rect 808 14300 2329 14328
rect 808 14288 814 14300
rect 2317 14297 2329 14300
rect 2363 14297 2375 14331
rect 3344 14328 3372 14359
rect 3694 14356 3700 14368
rect 3752 14356 3758 14408
rect 4522 14356 4528 14408
rect 4580 14356 4586 14408
rect 4724 14405 4752 14436
rect 5442 14424 5448 14476
rect 5500 14464 5506 14476
rect 5537 14467 5595 14473
rect 5537 14464 5549 14467
rect 5500 14436 5549 14464
rect 5500 14424 5506 14436
rect 5537 14433 5549 14436
rect 5583 14433 5595 14467
rect 5537 14427 5595 14433
rect 5644 14436 5856 14464
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 4801 14399 4859 14405
rect 4801 14365 4813 14399
rect 4847 14396 4859 14399
rect 5074 14396 5080 14408
rect 4847 14368 5080 14396
rect 4847 14365 4859 14368
rect 4801 14359 4859 14365
rect 4724 14328 4752 14359
rect 5074 14356 5080 14368
rect 5132 14396 5138 14408
rect 5644 14396 5672 14436
rect 5132 14368 5672 14396
rect 5132 14356 5138 14368
rect 5718 14356 5724 14408
rect 5776 14356 5782 14408
rect 5828 14405 5856 14436
rect 6270 14424 6276 14476
rect 6328 14424 6334 14476
rect 7466 14464 7472 14476
rect 6380 14436 7472 14464
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14396 5871 14399
rect 6380 14396 6408 14436
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 7650 14424 7656 14476
rect 7708 14464 7714 14476
rect 13170 14464 13176 14476
rect 7708 14436 10180 14464
rect 7708 14424 7714 14436
rect 5859 14368 6408 14396
rect 5859 14365 5871 14368
rect 5813 14359 5871 14365
rect 6454 14356 6460 14408
rect 6512 14356 6518 14408
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14396 6883 14399
rect 7374 14396 7380 14408
rect 6871 14368 7380 14396
rect 6871 14365 6883 14368
rect 6825 14359 6883 14365
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 7834 14356 7840 14408
rect 7892 14356 7898 14408
rect 8036 14405 8064 14436
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14396 8079 14399
rect 8202 14396 8208 14408
rect 8067 14368 8208 14396
rect 8067 14365 8079 14368
rect 8021 14359 8079 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8754 14356 8760 14408
rect 8812 14396 8818 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 8812 14368 9137 14396
rect 8812 14356 8818 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9214 14356 9220 14408
rect 9272 14356 9278 14408
rect 10152 14405 10180 14436
rect 10980 14436 13176 14464
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14365 9459 14399
rect 9401 14359 9459 14365
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 5994 14328 6000 14340
rect 3344 14300 4752 14328
rect 5184 14300 6000 14328
rect 2317 14291 2375 14297
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14260 2007 14263
rect 2038 14260 2044 14272
rect 1995 14232 2044 14260
rect 1995 14229 2007 14232
rect 1949 14223 2007 14229
rect 2038 14220 2044 14232
rect 2096 14260 2102 14272
rect 2682 14260 2688 14272
rect 2096 14232 2688 14260
rect 2096 14220 2102 14232
rect 2682 14220 2688 14232
rect 2740 14260 2746 14272
rect 3418 14260 3424 14272
rect 2740 14232 3424 14260
rect 2740 14220 2746 14232
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 5184 14260 5212 14300
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 7282 14288 7288 14340
rect 7340 14328 7346 14340
rect 9416 14328 9444 14359
rect 10778 14356 10784 14408
rect 10836 14356 10842 14408
rect 10980 14405 11008 14436
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 15010 14464 15016 14476
rect 13280 14436 15016 14464
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 13280 14405 13308 14436
rect 15010 14424 15016 14436
rect 15068 14424 15074 14476
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 11848 14368 13277 14396
rect 11848 14356 11854 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14396 13507 14399
rect 15286 14396 15292 14408
rect 13495 14368 15292 14396
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 7340 14300 9444 14328
rect 10689 14331 10747 14337
rect 7340 14288 7346 14300
rect 10689 14297 10701 14331
rect 10735 14328 10747 14331
rect 10735 14300 11008 14328
rect 10735 14297 10747 14300
rect 10689 14291 10747 14297
rect 10980 14272 11008 14300
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 13464 14328 13492 14359
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 12492 14300 13492 14328
rect 12492 14288 12498 14300
rect 13538 14288 13544 14340
rect 13596 14328 13602 14340
rect 19794 14328 19800 14340
rect 13596 14300 19800 14328
rect 13596 14288 13602 14300
rect 19794 14288 19800 14300
rect 19852 14288 19858 14340
rect 4212 14232 5212 14260
rect 4212 14220 4218 14232
rect 5258 14220 5264 14272
rect 5316 14260 5322 14272
rect 5353 14263 5411 14269
rect 5353 14260 5365 14263
rect 5316 14232 5365 14260
rect 5316 14220 5322 14232
rect 5353 14229 5365 14232
rect 5399 14229 5411 14263
rect 5353 14223 5411 14229
rect 6733 14263 6791 14269
rect 6733 14229 6745 14263
rect 6779 14260 6791 14263
rect 6822 14260 6828 14272
rect 6779 14232 6828 14260
rect 6779 14229 6791 14232
rect 6733 14223 6791 14229
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7929 14263 7987 14269
rect 7929 14229 7941 14263
rect 7975 14260 7987 14263
rect 8018 14260 8024 14272
rect 7975 14232 8024 14260
rect 7975 14229 7987 14232
rect 7929 14223 7987 14229
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 8754 14220 8760 14272
rect 8812 14260 8818 14272
rect 9398 14260 9404 14272
rect 8812 14232 9404 14260
rect 8812 14220 8818 14232
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 10962 14220 10968 14272
rect 11020 14220 11026 14272
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14260 13507 14263
rect 18966 14260 18972 14272
rect 13495 14232 18972 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 18966 14220 18972 14232
rect 19024 14220 19030 14272
rect 1104 14170 18860 14192
rect 1104 14118 5502 14170
rect 5554 14118 5566 14170
rect 5618 14118 5630 14170
rect 5682 14118 5694 14170
rect 5746 14118 5758 14170
rect 5810 14118 5822 14170
rect 5874 14118 5886 14170
rect 5938 14118 5950 14170
rect 6002 14118 6014 14170
rect 6066 14118 6078 14170
rect 6130 14118 6142 14170
rect 6194 14118 6206 14170
rect 6258 14118 6270 14170
rect 6322 14118 6334 14170
rect 6386 14118 6398 14170
rect 6450 14118 6462 14170
rect 6514 14118 6526 14170
rect 6578 14118 6590 14170
rect 6642 14118 6654 14170
rect 6706 14118 13502 14170
rect 13554 14118 13566 14170
rect 13618 14118 13630 14170
rect 13682 14118 13694 14170
rect 13746 14118 13758 14170
rect 13810 14118 13822 14170
rect 13874 14118 13886 14170
rect 13938 14118 13950 14170
rect 14002 14118 14014 14170
rect 14066 14118 14078 14170
rect 14130 14118 14142 14170
rect 14194 14118 14206 14170
rect 14258 14118 14270 14170
rect 14322 14118 14334 14170
rect 14386 14118 14398 14170
rect 14450 14118 14462 14170
rect 14514 14118 14526 14170
rect 14578 14118 14590 14170
rect 14642 14118 14654 14170
rect 14706 14118 18860 14170
rect 1104 14096 18860 14118
rect 1210 14016 1216 14068
rect 1268 14056 1274 14068
rect 3050 14056 3056 14068
rect 1268 14028 3056 14056
rect 1268 14016 1274 14028
rect 3050 14016 3056 14028
rect 3108 14056 3114 14068
rect 3108 14028 3280 14056
rect 3108 14016 3114 14028
rect 566 13988 572 14000
rect 492 13960 572 13988
rect 492 13784 520 13960
rect 566 13948 572 13960
rect 624 13948 630 14000
rect 1302 13948 1308 14000
rect 1360 13988 1366 14000
rect 2130 13988 2136 14000
rect 1360 13960 2136 13988
rect 1360 13948 1366 13960
rect 2130 13948 2136 13960
rect 2188 13948 2194 14000
rect 2866 13988 2872 14000
rect 2332 13960 2872 13988
rect 1118 13880 1124 13932
rect 1176 13920 1182 13932
rect 1897 13923 1955 13929
rect 1897 13920 1909 13923
rect 1176 13892 1909 13920
rect 1176 13880 1182 13892
rect 1897 13889 1909 13892
rect 1943 13889 1955 13923
rect 1897 13883 1955 13889
rect 2038 13880 2044 13932
rect 2096 13880 2102 13932
rect 2332 13929 2360 13960
rect 2866 13948 2872 13960
rect 2924 13948 2930 14000
rect 3252 13997 3280 14028
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 4249 14059 4307 14065
rect 4249 14056 4261 14059
rect 3476 14028 4261 14056
rect 3476 14016 3482 14028
rect 4249 14025 4261 14028
rect 4295 14025 4307 14059
rect 4249 14019 4307 14025
rect 4522 14016 4528 14068
rect 4580 14056 4586 14068
rect 5261 14059 5319 14065
rect 5261 14056 5273 14059
rect 4580 14028 5273 14056
rect 4580 14016 4586 14028
rect 5261 14025 5273 14028
rect 5307 14025 5319 14059
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 5261 14019 5319 14025
rect 6012 14028 7941 14056
rect 3237 13991 3295 13997
rect 3237 13957 3249 13991
rect 3283 13957 3295 13991
rect 3237 13951 3295 13957
rect 4430 13948 4436 14000
rect 4488 13988 4494 14000
rect 5902 13988 5908 14000
rect 4488 13960 5908 13988
rect 4488 13948 4494 13960
rect 5902 13948 5908 13960
rect 5960 13948 5966 14000
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13889 2375 13923
rect 3001 13923 3059 13929
rect 3001 13920 3013 13923
rect 2317 13883 2375 13889
rect 2608 13892 3013 13920
rect 566 13812 572 13864
rect 624 13852 630 13864
rect 624 13824 1256 13852
rect 624 13812 630 13824
rect 1228 13784 1256 13824
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 1578 13852 1584 13864
rect 1360 13824 1584 13852
rect 1360 13812 1366 13824
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 2608 13784 2636 13892
rect 3001 13889 3013 13892
rect 3047 13889 3059 13923
rect 3001 13883 3059 13889
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13920 3479 13923
rect 3970 13920 3976 13932
rect 3467 13892 3976 13920
rect 3467 13889 3479 13892
rect 3421 13883 3479 13889
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 3160 13852 3188 13883
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 4263 13892 4660 13920
rect 2740 13824 3188 13852
rect 4065 13855 4123 13861
rect 2740 13812 2746 13824
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4154 13852 4160 13864
rect 4111 13824 4160 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 4263 13784 4291 13892
rect 4433 13855 4491 13861
rect 4433 13821 4445 13855
rect 4479 13821 4491 13855
rect 4433 13815 4491 13821
rect 492 13756 612 13784
rect 1228 13756 2636 13784
rect 2700 13756 4291 13784
rect 584 13376 612 13756
rect 1210 13676 1216 13728
rect 1268 13716 1274 13728
rect 1765 13719 1823 13725
rect 1765 13716 1777 13719
rect 1268 13688 1777 13716
rect 1268 13676 1274 13688
rect 1765 13685 1777 13688
rect 1811 13685 1823 13719
rect 1765 13679 1823 13685
rect 1854 13676 1860 13728
rect 1912 13716 1918 13728
rect 2700 13716 2728 13756
rect 4448 13728 4476 13815
rect 4632 13784 4660 13892
rect 5074 13880 5080 13932
rect 5132 13880 5138 13932
rect 6012 13920 6040 14028
rect 7929 14025 7941 14028
rect 7975 14025 7987 14059
rect 9490 14056 9496 14068
rect 7929 14019 7987 14025
rect 8036 14028 9496 14056
rect 7282 13988 7288 14000
rect 6932 13960 7288 13988
rect 5167 13892 6040 13920
rect 4798 13812 4804 13864
rect 4856 13852 4862 13864
rect 5167 13852 5195 13892
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 6512 13892 6653 13920
rect 6512 13880 6518 13892
rect 6641 13889 6653 13892
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 4856 13824 5195 13852
rect 5445 13855 5503 13861
rect 4856 13812 4862 13824
rect 5445 13821 5457 13855
rect 5491 13821 5503 13855
rect 6932 13852 6960 13960
rect 7282 13948 7288 13960
rect 7340 13948 7346 14000
rect 8036 13988 8064 14028
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 15194 14056 15200 14068
rect 12544 14028 15200 14056
rect 7668 13960 8064 13988
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 7466 13920 7472 13932
rect 7055 13892 7472 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 5445 13815 5503 13821
rect 6656 13824 6960 13852
rect 5460 13784 5488 13815
rect 6656 13796 6684 13824
rect 7190 13812 7196 13864
rect 7248 13852 7254 13864
rect 7561 13855 7619 13861
rect 7561 13852 7573 13855
rect 7248 13824 7573 13852
rect 7248 13812 7254 13824
rect 7561 13821 7573 13824
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 6638 13784 6644 13796
rect 4632 13756 6644 13784
rect 1912 13688 2728 13716
rect 2869 13719 2927 13725
rect 1912 13676 1918 13688
rect 2869 13685 2881 13719
rect 2915 13716 2927 13719
rect 3050 13716 3056 13728
rect 2915 13688 3056 13716
rect 2915 13685 2927 13688
rect 2869 13679 2927 13685
rect 3050 13676 3056 13688
rect 3108 13676 3114 13728
rect 4430 13676 4436 13728
rect 4488 13676 4494 13728
rect 4632 13725 4660 13756
rect 6638 13744 6644 13756
rect 6696 13744 6702 13796
rect 7668 13784 7696 13960
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 8260 13960 8493 13988
rect 8260 13948 8266 13960
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 8570 13948 8576 14000
rect 8628 13988 8634 14000
rect 9030 13988 9036 14000
rect 8628 13960 9036 13988
rect 8628 13948 8634 13960
rect 9030 13948 9036 13960
rect 9088 13988 9094 14000
rect 9088 13960 10272 13988
rect 9088 13948 9094 13960
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 7760 13852 7788 13883
rect 7834 13880 7840 13932
rect 7892 13920 7898 13932
rect 8665 13923 8723 13929
rect 8665 13920 8677 13923
rect 7892 13892 8677 13920
rect 7892 13880 7898 13892
rect 8665 13889 8677 13892
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 9309 13923 9367 13929
rect 9309 13889 9321 13923
rect 9355 13889 9367 13923
rect 9309 13883 9367 13889
rect 7760 13824 8064 13852
rect 6748 13756 7696 13784
rect 4617 13719 4675 13725
rect 4617 13685 4629 13719
rect 4663 13685 4675 13719
rect 4617 13679 4675 13685
rect 5626 13676 5632 13728
rect 5684 13716 5690 13728
rect 6748 13716 6776 13756
rect 5684 13688 6776 13716
rect 5684 13676 5690 13688
rect 6914 13676 6920 13728
rect 6972 13676 6978 13728
rect 7926 13676 7932 13728
rect 7984 13716 7990 13728
rect 8036 13716 8064 13824
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 9324 13852 9352 13883
rect 9490 13880 9496 13932
rect 9548 13880 9554 13932
rect 10244 13929 10272 13960
rect 11974 13948 11980 14000
rect 12032 13988 12038 14000
rect 12544 13997 12572 14028
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 12069 13991 12127 13997
rect 12069 13988 12081 13991
rect 12032 13960 12081 13988
rect 12032 13948 12038 13960
rect 12069 13957 12081 13960
rect 12115 13957 12127 13991
rect 12069 13951 12127 13957
rect 12529 13991 12587 13997
rect 12529 13957 12541 13991
rect 12575 13957 12587 13991
rect 12529 13951 12587 13957
rect 12713 13991 12771 13997
rect 12713 13957 12725 13991
rect 12759 13988 12771 13991
rect 12986 13988 12992 14000
rect 12759 13960 12992 13988
rect 12759 13957 12771 13960
rect 12713 13951 12771 13957
rect 12986 13948 12992 13960
rect 13044 13948 13050 14000
rect 13354 13948 13360 14000
rect 13412 13988 13418 14000
rect 13449 13991 13507 13997
rect 13449 13988 13461 13991
rect 13412 13960 13461 13988
rect 13412 13948 13418 13960
rect 13449 13957 13461 13960
rect 13495 13957 13507 13991
rect 14461 13991 14519 13997
rect 13449 13951 13507 13957
rect 13648 13960 14228 13988
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13889 10287 13923
rect 10229 13883 10287 13889
rect 8352 13824 9352 13852
rect 10244 13852 10272 13883
rect 10318 13880 10324 13932
rect 10376 13920 10382 13932
rect 11790 13920 11796 13932
rect 10376 13892 11796 13920
rect 10376 13880 10382 13892
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 11931 13892 12756 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12728 13864 12756 13892
rect 12894 13880 12900 13932
rect 12952 13880 12958 13932
rect 13648 13929 13676 13960
rect 13633 13923 13691 13929
rect 13633 13889 13645 13923
rect 13679 13889 13691 13923
rect 13633 13883 13691 13889
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 12434 13852 12440 13864
rect 10244 13824 12440 13852
rect 8352 13812 8358 13824
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12710 13812 12716 13864
rect 12768 13812 12774 13864
rect 13078 13812 13084 13864
rect 13136 13852 13142 13864
rect 13740 13852 13768 13883
rect 13136 13824 13768 13852
rect 13136 13812 13142 13824
rect 8846 13744 8852 13796
rect 8904 13744 8910 13796
rect 9585 13787 9643 13793
rect 9585 13753 9597 13787
rect 9631 13753 9643 13787
rect 9585 13747 9643 13753
rect 10413 13787 10471 13793
rect 10413 13753 10425 13787
rect 10459 13784 10471 13787
rect 14200 13784 14228 13960
rect 14461 13957 14473 13991
rect 14507 13988 14519 13991
rect 14826 13988 14832 14000
rect 14507 13960 14832 13988
rect 14507 13957 14519 13960
rect 14461 13951 14519 13957
rect 14826 13948 14832 13960
rect 14884 13948 14890 14000
rect 14918 13948 14924 14000
rect 14976 13988 14982 14000
rect 19334 13988 19340 14000
rect 14976 13960 19340 13988
rect 14976 13948 14982 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13920 14703 13923
rect 19886 13920 19892 13932
rect 14691 13892 19892 13920
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 19886 13880 19892 13892
rect 19944 13880 19950 13932
rect 14277 13855 14335 13861
rect 14277 13821 14289 13855
rect 14323 13852 14335 13855
rect 19610 13852 19616 13864
rect 14323 13824 19616 13852
rect 14323 13821 14335 13824
rect 14277 13815 14335 13821
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 14918 13784 14924 13796
rect 10459 13756 12354 13784
rect 14200 13756 14924 13784
rect 10459 13753 10471 13756
rect 10413 13747 10471 13753
rect 7984 13688 8064 13716
rect 7984 13676 7990 13688
rect 8570 13676 8576 13728
rect 8628 13716 8634 13728
rect 9600 13716 9628 13747
rect 8628 13688 9628 13716
rect 8628 13676 8634 13688
rect 11790 13676 11796 13728
rect 11848 13676 11854 13728
rect 12326 13716 12354 13756
rect 14918 13744 14924 13756
rect 14976 13744 14982 13796
rect 16298 13716 16304 13728
rect 12326 13688 16304 13716
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 1104 13626 18860 13648
rect 1104 13574 1502 13626
rect 1554 13574 1566 13626
rect 1618 13574 1630 13626
rect 1682 13574 1694 13626
rect 1746 13574 1758 13626
rect 1810 13574 1822 13626
rect 1874 13574 1886 13626
rect 1938 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 2270 13626
rect 2322 13574 2334 13626
rect 2386 13574 2398 13626
rect 2450 13574 2462 13626
rect 2514 13574 2526 13626
rect 2578 13574 2590 13626
rect 2642 13574 2654 13626
rect 2706 13574 9502 13626
rect 9554 13574 9566 13626
rect 9618 13574 9630 13626
rect 9682 13574 9694 13626
rect 9746 13574 9758 13626
rect 9810 13574 9822 13626
rect 9874 13574 9886 13626
rect 9938 13574 9950 13626
rect 10002 13574 10014 13626
rect 10066 13574 10078 13626
rect 10130 13574 10142 13626
rect 10194 13574 10206 13626
rect 10258 13574 10270 13626
rect 10322 13574 10334 13626
rect 10386 13574 10398 13626
rect 10450 13574 10462 13626
rect 10514 13574 10526 13626
rect 10578 13574 10590 13626
rect 10642 13574 10654 13626
rect 10706 13574 17502 13626
rect 17554 13574 17566 13626
rect 17618 13574 17630 13626
rect 17682 13574 17694 13626
rect 17746 13574 17758 13626
rect 17810 13574 17822 13626
rect 17874 13574 17886 13626
rect 17938 13574 17950 13626
rect 18002 13574 18014 13626
rect 18066 13574 18078 13626
rect 18130 13574 18142 13626
rect 18194 13574 18206 13626
rect 18258 13574 18270 13626
rect 18322 13574 18334 13626
rect 18386 13574 18398 13626
rect 18450 13574 18462 13626
rect 18514 13574 18526 13626
rect 18578 13574 18590 13626
rect 18642 13574 18654 13626
rect 18706 13574 18860 13626
rect 1104 13552 18860 13574
rect 658 13472 664 13524
rect 716 13512 722 13524
rect 2222 13512 2228 13524
rect 716 13484 2228 13512
rect 716 13472 722 13484
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 2372 13484 4077 13512
rect 2372 13472 2378 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4982 13512 4988 13524
rect 4065 13475 4123 13481
rect 4356 13484 4988 13512
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 2866 13444 2872 13456
rect 1627 13416 2872 13444
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 2866 13404 2872 13416
rect 2924 13404 2930 13456
rect 2884 13376 2912 13404
rect 584 13348 2452 13376
rect 2884 13348 3740 13376
rect 2424 13320 2452 13348
rect 1762 13268 1768 13320
rect 1820 13268 1826 13320
rect 2406 13268 2412 13320
rect 2464 13268 2470 13320
rect 2498 13268 2504 13320
rect 2556 13308 2562 13320
rect 2866 13317 2872 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2556 13280 2697 13308
rect 2556 13268 2562 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 2829 13311 2872 13317
rect 2829 13277 2841 13311
rect 2829 13271 2872 13277
rect 2866 13268 2872 13271
rect 2924 13268 2930 13320
rect 1946 13200 1952 13252
rect 2004 13200 2010 13252
rect 2590 13200 2596 13252
rect 2648 13200 2654 13252
rect 3712 13240 3740 13348
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 4356 13317 4384 13484
rect 4982 13472 4988 13484
rect 5040 13472 5046 13524
rect 5166 13472 5172 13524
rect 5224 13512 5230 13524
rect 5442 13512 5448 13524
rect 5224 13484 5448 13512
rect 5224 13472 5230 13484
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 6089 13515 6147 13521
rect 6089 13512 6101 13515
rect 5592 13484 6101 13512
rect 5592 13472 5598 13484
rect 6089 13481 6101 13484
rect 6135 13512 6147 13515
rect 6822 13512 6828 13524
rect 6135 13484 6828 13512
rect 6135 13481 6147 13484
rect 6089 13475 6147 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 7524 13484 9168 13512
rect 7524 13472 7530 13484
rect 4798 13444 4804 13456
rect 4540 13416 4804 13444
rect 4540 13317 4568 13416
rect 4798 13404 4804 13416
rect 4856 13404 4862 13456
rect 5350 13404 5356 13456
rect 5408 13444 5414 13456
rect 5626 13444 5632 13456
rect 5408 13416 5632 13444
rect 5408 13404 5414 13416
rect 5626 13404 5632 13416
rect 5684 13404 5690 13456
rect 6273 13379 6331 13385
rect 6273 13376 6285 13379
rect 5532 13348 6285 13376
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 4212 13280 4261 13308
rect 4212 13268 4218 13280
rect 4249 13277 4261 13280
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 4341 13311 4399 13317
rect 4341 13277 4353 13311
rect 4387 13277 4399 13311
rect 4341 13271 4399 13277
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13277 4491 13311
rect 4433 13271 4491 13277
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 4448 13240 4476 13271
rect 3712 13212 4476 13240
rect 4540 13240 4568 13271
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 4856 13280 5181 13308
rect 4856 13268 4862 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 5532 13308 5560 13348
rect 6273 13345 6285 13348
rect 6319 13376 6331 13379
rect 7484 13376 7512 13472
rect 8202 13404 8208 13456
rect 8260 13404 8266 13456
rect 8754 13444 8760 13456
rect 8312 13416 8760 13444
rect 6319 13348 7512 13376
rect 6319 13345 6331 13348
rect 6273 13339 6331 13345
rect 7834 13336 7840 13388
rect 7892 13376 7898 13388
rect 8018 13376 8024 13388
rect 7892 13348 8024 13376
rect 7892 13336 7898 13348
rect 8018 13336 8024 13348
rect 8076 13336 8082 13388
rect 5491 13280 5560 13308
rect 5997 13311 6055 13317
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 5997 13277 6009 13311
rect 6043 13308 6055 13311
rect 6454 13308 6460 13320
rect 6043 13280 6460 13308
rect 6043 13277 6055 13280
rect 5997 13271 6055 13277
rect 5074 13240 5080 13252
rect 4540 13212 5080 13240
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 5184 13240 5212 13271
rect 6012 13240 6040 13271
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 8312 13317 8340 13416
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 9140 13444 9168 13484
rect 9214 13472 9220 13524
rect 9272 13512 9278 13524
rect 12434 13512 12440 13524
rect 9272 13484 12440 13512
rect 9272 13472 9278 13484
rect 12434 13472 12440 13484
rect 12492 13512 12498 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 12492 13484 12725 13512
rect 12492 13472 12498 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 12713 13475 12771 13481
rect 12618 13444 12624 13456
rect 9140 13416 12624 13444
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 12158 13376 12164 13388
rect 11848 13348 12164 13376
rect 11848 13336 11854 13348
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 15102 13376 15108 13388
rect 14384 13348 15108 13376
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6696 13280 6929 13308
rect 6696 13268 6702 13280
rect 6917 13277 6929 13280
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13308 7343 13311
rect 8297 13311 8355 13317
rect 7331 13280 8248 13308
rect 7331 13277 7343 13280
rect 7285 13271 7343 13277
rect 5184 13212 6040 13240
rect 6472 13240 6500 13268
rect 7300 13240 7328 13271
rect 6472 13212 7328 13240
rect 7834 13200 7840 13252
rect 7892 13240 7898 13252
rect 7929 13243 7987 13249
rect 7929 13240 7941 13243
rect 7892 13212 7941 13240
rect 7892 13200 7898 13212
rect 7929 13209 7941 13212
rect 7975 13209 7987 13243
rect 8220 13240 8248 13280
rect 8297 13277 8309 13311
rect 8343 13277 8355 13311
rect 8297 13271 8355 13277
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13308 8539 13311
rect 8754 13308 8760 13320
rect 8527 13280 8760 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 9582 13268 9588 13320
rect 9640 13268 9646 13320
rect 9766 13268 9772 13320
rect 9824 13268 9830 13320
rect 10134 13268 10140 13320
rect 10192 13268 10198 13320
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 10873 13311 10931 13317
rect 10873 13308 10885 13311
rect 10468 13280 10885 13308
rect 10468 13268 10474 13280
rect 10873 13277 10885 13280
rect 10919 13277 10931 13311
rect 10873 13271 10931 13277
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13308 11115 13311
rect 11238 13308 11244 13320
rect 11103 13280 11244 13308
rect 11103 13277 11115 13280
rect 11057 13271 11115 13277
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 11606 13268 11612 13320
rect 11664 13268 11670 13320
rect 11977 13311 12035 13317
rect 11977 13277 11989 13311
rect 12023 13308 12035 13311
rect 12023 13280 12112 13308
rect 12023 13277 12035 13280
rect 11977 13271 12035 13277
rect 8220 13212 9628 13240
rect 7929 13203 7987 13209
rect 474 13132 480 13184
rect 532 13172 538 13184
rect 2866 13172 2872 13184
rect 532 13144 2872 13172
rect 532 13132 538 13144
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 2978 13175 3036 13181
rect 2978 13141 2990 13175
rect 3024 13172 3036 13175
rect 4154 13172 4160 13184
rect 3024 13144 4160 13172
rect 3024 13141 3036 13144
rect 2978 13135 3036 13141
rect 4154 13132 4160 13144
rect 4212 13132 4218 13184
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 7101 13175 7159 13181
rect 7101 13172 7113 13175
rect 5500 13144 7113 13172
rect 5500 13132 5506 13144
rect 7101 13141 7113 13144
rect 7147 13172 7159 13175
rect 7282 13172 7288 13184
rect 7147 13144 7288 13172
rect 7147 13141 7159 13144
rect 7101 13135 7159 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 9600 13172 9628 13212
rect 9950 13172 9956 13184
rect 9600 13144 9956 13172
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 10045 13175 10103 13181
rect 10045 13141 10057 13175
rect 10091 13172 10103 13175
rect 10594 13172 10600 13184
rect 10091 13144 10600 13172
rect 10091 13141 10103 13144
rect 10045 13135 10103 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 10689 13175 10747 13181
rect 10689 13141 10701 13175
rect 10735 13172 10747 13175
rect 10778 13172 10784 13184
rect 10735 13144 10784 13172
rect 10735 13141 10747 13144
rect 10689 13135 10747 13141
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 11974 13132 11980 13184
rect 12032 13132 12038 13184
rect 12084 13172 12112 13280
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 14384 13317 14412 13348
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 16206 13376 16212 13388
rect 15344 13348 16212 13376
rect 15344 13336 15350 13348
rect 16206 13336 16212 13348
rect 16264 13376 16270 13388
rect 16264 13348 16620 13376
rect 16264 13336 16270 13348
rect 12805 13311 12863 13317
rect 12805 13308 12817 13311
rect 12676 13280 12817 13308
rect 12676 13268 12682 13280
rect 12805 13277 12817 13280
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13308 14611 13311
rect 14734 13308 14740 13320
rect 14599 13280 14740 13308
rect 14599 13277 14611 13280
rect 14553 13271 14611 13277
rect 14734 13268 14740 13280
rect 14792 13308 14798 13320
rect 14918 13308 14924 13320
rect 14792 13280 14924 13308
rect 14792 13268 14798 13280
rect 14918 13268 14924 13280
rect 14976 13268 14982 13320
rect 16390 13268 16396 13320
rect 16448 13268 16454 13320
rect 16592 13317 16620 13348
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13308 16635 13311
rect 17126 13308 17132 13320
rect 16623 13280 17132 13308
rect 16623 13277 16635 13280
rect 16577 13271 16635 13277
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 12989 13243 13047 13249
rect 12989 13240 13001 13243
rect 12768 13212 13001 13240
rect 12768 13200 12774 13212
rect 12989 13209 13001 13212
rect 13035 13209 13047 13243
rect 12989 13203 13047 13209
rect 14645 13243 14703 13249
rect 14645 13209 14657 13243
rect 14691 13240 14703 13243
rect 15930 13240 15936 13252
rect 14691 13212 15936 13240
rect 14691 13209 14703 13212
rect 14645 13203 14703 13209
rect 15930 13200 15936 13212
rect 15988 13200 15994 13252
rect 13354 13172 13360 13184
rect 12084 13144 13360 13172
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 16393 13175 16451 13181
rect 16393 13172 16405 13175
rect 15436 13144 16405 13172
rect 15436 13132 15442 13144
rect 16393 13141 16405 13144
rect 16439 13141 16451 13175
rect 16393 13135 16451 13141
rect 1104 13082 18860 13104
rect 14 12996 20 13048
rect 72 13036 78 13048
rect 474 13036 480 13048
rect 72 13008 480 13036
rect 72 12996 78 13008
rect 474 12996 480 13008
rect 532 12996 538 13048
rect 1104 13030 5502 13082
rect 5554 13030 5566 13082
rect 5618 13030 5630 13082
rect 5682 13030 5694 13082
rect 5746 13030 5758 13082
rect 5810 13030 5822 13082
rect 5874 13030 5886 13082
rect 5938 13030 5950 13082
rect 6002 13030 6014 13082
rect 6066 13030 6078 13082
rect 6130 13030 6142 13082
rect 6194 13030 6206 13082
rect 6258 13030 6270 13082
rect 6322 13030 6334 13082
rect 6386 13030 6398 13082
rect 6450 13030 6462 13082
rect 6514 13030 6526 13082
rect 6578 13030 6590 13082
rect 6642 13030 6654 13082
rect 6706 13030 13502 13082
rect 13554 13030 13566 13082
rect 13618 13030 13630 13082
rect 13682 13030 13694 13082
rect 13746 13030 13758 13082
rect 13810 13030 13822 13082
rect 13874 13030 13886 13082
rect 13938 13030 13950 13082
rect 14002 13030 14014 13082
rect 14066 13030 14078 13082
rect 14130 13030 14142 13082
rect 14194 13030 14206 13082
rect 14258 13030 14270 13082
rect 14322 13030 14334 13082
rect 14386 13030 14398 13082
rect 14450 13030 14462 13082
rect 14514 13030 14526 13082
rect 14578 13030 14590 13082
rect 14642 13030 14654 13082
rect 14706 13030 18860 13082
rect 1104 13008 18860 13030
rect 1302 12968 1308 12980
rect 32 12940 1308 12968
rect 32 12912 60 12940
rect 1302 12928 1308 12940
rect 1360 12928 1366 12980
rect 2314 12928 2320 12980
rect 2372 12928 2378 12980
rect 2409 12971 2467 12977
rect 2409 12937 2421 12971
rect 2455 12968 2467 12971
rect 2682 12968 2688 12980
rect 2455 12940 2688 12968
rect 2455 12937 2467 12940
rect 2409 12931 2467 12937
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 2832 12940 4108 12968
rect 2832 12928 2838 12940
rect 14 12860 20 12912
rect 72 12860 78 12912
rect 106 12860 112 12912
rect 164 12900 170 12912
rect 164 12872 2774 12900
rect 164 12860 170 12872
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 1964 12696 1992 12795
rect 2406 12792 2412 12844
rect 2464 12832 2470 12844
rect 2746 12832 2774 12872
rect 3510 12860 3516 12912
rect 3568 12900 3574 12912
rect 3694 12900 3700 12912
rect 3568 12872 3700 12900
rect 3568 12860 3574 12872
rect 3694 12860 3700 12872
rect 3752 12860 3758 12912
rect 4080 12909 4108 12940
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 6178 12968 6184 12980
rect 4212 12940 6184 12968
rect 4212 12928 4218 12940
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 6932 12940 8156 12968
rect 4065 12903 4123 12909
rect 4065 12869 4077 12903
rect 4111 12900 4123 12903
rect 4430 12900 4436 12912
rect 4111 12872 4436 12900
rect 4111 12869 4123 12872
rect 4065 12863 4123 12869
rect 4430 12860 4436 12872
rect 4488 12860 4494 12912
rect 4982 12860 4988 12912
rect 5040 12900 5046 12912
rect 5169 12903 5227 12909
rect 5169 12900 5181 12903
rect 5040 12872 5181 12900
rect 5040 12860 5046 12872
rect 5169 12869 5181 12872
rect 5215 12869 5227 12903
rect 6932 12900 6960 12940
rect 5169 12863 5227 12869
rect 5644 12872 6960 12900
rect 3835 12835 3893 12841
rect 3835 12832 3847 12835
rect 2464 12804 2636 12832
rect 2746 12804 3847 12832
rect 2464 12792 2470 12804
rect 2222 12773 2228 12776
rect 2208 12767 2228 12773
rect 2208 12733 2220 12767
rect 2208 12727 2228 12733
rect 2222 12724 2228 12727
rect 2280 12724 2286 12776
rect 2314 12724 2320 12776
rect 2372 12764 2378 12776
rect 2501 12767 2559 12773
rect 2501 12764 2513 12767
rect 2372 12736 2513 12764
rect 2372 12724 2378 12736
rect 2501 12733 2513 12736
rect 2547 12733 2559 12767
rect 2608 12764 2636 12804
rect 3835 12801 3847 12804
rect 3881 12801 3893 12835
rect 3835 12795 3893 12801
rect 3973 12835 4031 12841
rect 3973 12801 3985 12835
rect 4019 12801 4031 12835
rect 4246 12832 4252 12844
rect 4207 12804 4252 12832
rect 3973 12795 4031 12801
rect 2774 12764 2780 12776
rect 2608 12736 2780 12764
rect 2501 12727 2559 12733
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 3234 12764 3240 12776
rect 2924 12736 3240 12764
rect 2924 12724 2930 12736
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3988 12764 4016 12795
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 4338 12792 4344 12844
rect 4396 12792 4402 12844
rect 5353 12767 5411 12773
rect 5353 12764 5365 12767
rect 3620 12736 4016 12764
rect 5276 12736 5365 12764
rect 2590 12696 2596 12708
rect 1044 12668 2596 12696
rect 1044 12424 1072 12668
rect 2590 12656 2596 12668
rect 2648 12696 2654 12708
rect 3620 12696 3648 12736
rect 5276 12708 5304 12736
rect 5353 12733 5365 12736
rect 5399 12733 5411 12767
rect 5442 12758 5448 12810
rect 5500 12758 5506 12810
rect 5534 12792 5540 12844
rect 5592 12792 5598 12844
rect 5644 12841 5672 12872
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 6730 12832 6736 12844
rect 6687 12804 6736 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 5828 12764 5856 12795
rect 6730 12792 6736 12804
rect 6788 12792 6794 12844
rect 6822 12792 6828 12844
rect 6880 12792 6886 12844
rect 6932 12841 6960 12872
rect 7190 12860 7196 12912
rect 7248 12860 7254 12912
rect 7558 12860 7564 12912
rect 7616 12900 7622 12912
rect 7653 12903 7711 12909
rect 7653 12900 7665 12903
rect 7616 12872 7665 12900
rect 7616 12860 7622 12872
rect 7653 12869 7665 12872
rect 7699 12869 7711 12903
rect 7653 12863 7711 12869
rect 7745 12903 7803 12909
rect 7745 12869 7757 12903
rect 7791 12900 7803 12903
rect 8128 12900 8156 12940
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 8352 12940 10977 12968
rect 8352 12928 8358 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 12618 12968 12624 12980
rect 10965 12931 11023 12937
rect 11808 12940 12624 12968
rect 8846 12900 8852 12912
rect 7791 12872 8064 12900
rect 8128 12872 8852 12900
rect 7791 12869 7803 12872
rect 7745 12863 7803 12869
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12801 6975 12835
rect 7208 12832 7236 12860
rect 6917 12795 6975 12801
rect 7024 12804 7236 12832
rect 5994 12764 6000 12776
rect 5828 12736 6000 12764
rect 5353 12727 5411 12733
rect 5994 12724 6000 12736
rect 6052 12764 6058 12776
rect 7024 12764 7052 12804
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7760 12832 7788 12863
rect 7432 12804 7788 12832
rect 7432 12792 7438 12804
rect 7926 12792 7932 12844
rect 7984 12792 7990 12844
rect 8036 12832 8064 12872
rect 8846 12860 8852 12872
rect 8904 12860 8910 12912
rect 9950 12860 9956 12912
rect 10008 12900 10014 12912
rect 11808 12900 11836 12940
rect 12618 12928 12624 12940
rect 12676 12968 12682 12980
rect 13170 12968 13176 12980
rect 12676 12940 13176 12968
rect 12676 12928 12682 12940
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 16209 12971 16267 12977
rect 16209 12937 16221 12971
rect 16255 12968 16267 12971
rect 19242 12968 19248 12980
rect 16255 12940 19248 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 10008 12872 11836 12900
rect 10008 12860 10014 12872
rect 8036 12804 8340 12832
rect 6052 12736 7052 12764
rect 6052 12724 6058 12736
rect 7190 12724 7196 12776
rect 7248 12764 7254 12776
rect 8202 12764 8208 12776
rect 7248 12736 8208 12764
rect 7248 12724 7254 12736
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8312 12764 8340 12804
rect 8662 12792 8668 12844
rect 8720 12832 8726 12844
rect 9217 12835 9275 12841
rect 9217 12832 9229 12835
rect 8720 12804 9229 12832
rect 8720 12792 8726 12804
rect 9217 12801 9229 12804
rect 9263 12832 9275 12835
rect 9490 12832 9496 12844
rect 9263 12804 9496 12832
rect 9263 12801 9275 12804
rect 9217 12795 9275 12801
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 9582 12792 9588 12844
rect 9640 12832 9646 12844
rect 9640 12804 10640 12832
rect 9640 12792 9646 12804
rect 9030 12764 9036 12776
rect 8312 12736 9036 12764
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 9401 12767 9459 12773
rect 9401 12733 9413 12767
rect 9447 12733 9459 12767
rect 9401 12727 9459 12733
rect 2648 12668 3648 12696
rect 2648 12656 2654 12668
rect 1486 12588 1492 12640
rect 1544 12628 1550 12640
rect 1854 12628 1860 12640
rect 1544 12600 1860 12628
rect 1544 12588 1550 12600
rect 1854 12588 1860 12600
rect 1912 12588 1918 12640
rect 1949 12631 2007 12637
rect 1949 12597 1961 12631
rect 1995 12628 2007 12631
rect 2958 12628 2964 12640
rect 1995 12600 2964 12628
rect 1995 12597 2007 12600
rect 1949 12591 2007 12597
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 3620 12628 3648 12668
rect 3697 12699 3755 12705
rect 3697 12665 3709 12699
rect 3743 12696 3755 12699
rect 5166 12696 5172 12708
rect 3743 12668 5172 12696
rect 3743 12665 3755 12668
rect 3697 12659 3755 12665
rect 5166 12656 5172 12668
rect 5224 12656 5230 12708
rect 5258 12656 5264 12708
rect 5316 12696 5322 12708
rect 6546 12696 6552 12708
rect 5316 12668 6552 12696
rect 5316 12656 5322 12668
rect 6546 12656 6552 12668
rect 6604 12656 6610 12708
rect 6638 12656 6644 12708
rect 6696 12696 6702 12708
rect 6914 12696 6920 12708
rect 6696 12668 6920 12696
rect 6696 12656 6702 12668
rect 6914 12656 6920 12668
rect 6972 12656 6978 12708
rect 9214 12696 9220 12708
rect 7484 12668 9220 12696
rect 5902 12628 5908 12640
rect 3620 12600 5908 12628
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 7101 12631 7159 12637
rect 7101 12628 7113 12631
rect 6420 12600 7113 12628
rect 6420 12588 6426 12600
rect 7101 12597 7113 12600
rect 7147 12628 7159 12631
rect 7484 12628 7512 12668
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 9416 12696 9444 12727
rect 9766 12724 9772 12776
rect 9824 12764 9830 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 9824 12736 10057 12764
rect 9824 12724 9830 12736
rect 10045 12733 10057 12736
rect 10091 12764 10103 12767
rect 10502 12764 10508 12776
rect 10091 12736 10508 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 10612 12773 10640 12804
rect 10778 12792 10784 12844
rect 10836 12792 10842 12844
rect 11054 12792 11060 12844
rect 11112 12792 11118 12844
rect 11808 12841 11836 12872
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 13265 12903 13323 12909
rect 13265 12900 13277 12903
rect 12124 12872 13277 12900
rect 12124 12860 12130 12872
rect 13265 12869 13277 12872
rect 13311 12869 13323 12903
rect 15470 12900 15476 12912
rect 13265 12863 13323 12869
rect 15212 12872 15476 12900
rect 11888 12844 11940 12850
rect 11793 12835 11851 12841
rect 11793 12801 11805 12835
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 14277 12835 14335 12841
rect 14277 12832 14289 12835
rect 12952 12804 14289 12832
rect 12952 12792 12958 12804
rect 14277 12801 14289 12804
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 11888 12786 11940 12792
rect 10597 12767 10655 12773
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 11330 12764 11336 12776
rect 10643 12736 11336 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 10410 12696 10416 12708
rect 9416 12668 10416 12696
rect 10410 12656 10416 12668
rect 10468 12696 10474 12708
rect 11900 12696 11928 12786
rect 12710 12724 12716 12776
rect 12768 12724 12774 12776
rect 12986 12724 12992 12776
rect 13044 12764 13050 12776
rect 14568 12764 14596 12795
rect 15010 12792 15016 12844
rect 15068 12832 15074 12844
rect 15212 12841 15240 12872
rect 15470 12860 15476 12872
rect 15528 12900 15534 12912
rect 16390 12900 16396 12912
rect 15528 12872 16396 12900
rect 15528 12860 15534 12872
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 15068 12804 15209 12832
rect 15068 12792 15074 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 15197 12795 15255 12801
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 16040 12841 16068 12872
rect 16390 12860 16396 12872
rect 16448 12900 16454 12912
rect 16448 12872 16988 12900
rect 16448 12860 16454 12872
rect 15381 12835 15439 12841
rect 15381 12832 15393 12835
rect 15344 12804 15393 12832
rect 15344 12792 15350 12804
rect 15381 12801 15393 12804
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 16206 12792 16212 12844
rect 16264 12792 16270 12844
rect 16960 12841 16988 12872
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 17126 12792 17132 12844
rect 17184 12792 17190 12844
rect 16850 12764 16856 12776
rect 13044 12736 16856 12764
rect 13044 12724 13050 12736
rect 16850 12724 16856 12736
rect 16908 12724 16914 12776
rect 10468 12668 11928 12696
rect 10468 12656 10474 12668
rect 13446 12656 13452 12708
rect 13504 12696 13510 12708
rect 13541 12699 13599 12705
rect 13541 12696 13553 12699
rect 13504 12668 13553 12696
rect 13504 12656 13510 12668
rect 13541 12665 13553 12668
rect 13587 12665 13599 12699
rect 13541 12659 13599 12665
rect 15197 12699 15255 12705
rect 15197 12665 15209 12699
rect 15243 12665 15255 12699
rect 15197 12659 15255 12665
rect 16945 12699 17003 12705
rect 16945 12665 16957 12699
rect 16991 12696 17003 12699
rect 19518 12696 19524 12708
rect 16991 12668 19524 12696
rect 16991 12665 17003 12668
rect 16945 12659 17003 12665
rect 7147 12600 7512 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7650 12588 7656 12640
rect 7708 12628 7714 12640
rect 8113 12631 8171 12637
rect 8113 12628 8125 12631
rect 7708 12600 8125 12628
rect 7708 12588 7714 12600
rect 8113 12597 8125 12600
rect 8159 12597 8171 12631
rect 8113 12591 8171 12597
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 10870 12628 10876 12640
rect 10652 12600 10876 12628
rect 10652 12588 10658 12600
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 13170 12588 13176 12640
rect 13228 12628 13234 12640
rect 13725 12631 13783 12637
rect 13725 12628 13737 12631
rect 13228 12600 13737 12628
rect 13228 12588 13234 12600
rect 13725 12597 13737 12600
rect 13771 12597 13783 12631
rect 13725 12591 13783 12597
rect 14366 12588 14372 12640
rect 14424 12588 14430 12640
rect 15212 12628 15240 12659
rect 19518 12656 19524 12668
rect 19576 12656 19582 12708
rect 19702 12628 19708 12640
rect 15212 12600 19708 12628
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 1104 12538 18860 12560
rect 1104 12486 1502 12538
rect 1554 12486 1566 12538
rect 1618 12486 1630 12538
rect 1682 12486 1694 12538
rect 1746 12486 1758 12538
rect 1810 12486 1822 12538
rect 1874 12486 1886 12538
rect 1938 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 2270 12538
rect 2322 12486 2334 12538
rect 2386 12486 2398 12538
rect 2450 12486 2462 12538
rect 2514 12486 2526 12538
rect 2578 12486 2590 12538
rect 2642 12486 2654 12538
rect 2706 12486 9502 12538
rect 9554 12486 9566 12538
rect 9618 12486 9630 12538
rect 9682 12486 9694 12538
rect 9746 12486 9758 12538
rect 9810 12486 9822 12538
rect 9874 12486 9886 12538
rect 9938 12486 9950 12538
rect 10002 12486 10014 12538
rect 10066 12486 10078 12538
rect 10130 12486 10142 12538
rect 10194 12486 10206 12538
rect 10258 12486 10270 12538
rect 10322 12486 10334 12538
rect 10386 12486 10398 12538
rect 10450 12486 10462 12538
rect 10514 12486 10526 12538
rect 10578 12486 10590 12538
rect 10642 12486 10654 12538
rect 10706 12486 17502 12538
rect 17554 12486 17566 12538
rect 17618 12486 17630 12538
rect 17682 12486 17694 12538
rect 17746 12486 17758 12538
rect 17810 12486 17822 12538
rect 17874 12486 17886 12538
rect 17938 12486 17950 12538
rect 18002 12486 18014 12538
rect 18066 12486 18078 12538
rect 18130 12486 18142 12538
rect 18194 12486 18206 12538
rect 18258 12486 18270 12538
rect 18322 12486 18334 12538
rect 18386 12486 18398 12538
rect 18450 12486 18462 12538
rect 18514 12486 18526 12538
rect 18578 12486 18590 12538
rect 18642 12486 18654 12538
rect 18706 12486 18860 12538
rect 1104 12464 18860 12486
rect 1762 12424 1768 12436
rect 1044 12396 1768 12424
rect 1762 12384 1768 12396
rect 1820 12384 1826 12436
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 2924 12396 3096 12424
rect 2924 12384 2930 12396
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 2498 12356 2504 12368
rect 1903 12328 2504 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 2498 12316 2504 12328
rect 2556 12316 2562 12368
rect 842 12248 848 12300
rect 900 12288 906 12300
rect 2113 12291 2171 12297
rect 2113 12288 2125 12291
rect 900 12260 2125 12288
rect 900 12248 906 12260
rect 2113 12257 2125 12260
rect 2159 12257 2171 12291
rect 2113 12251 2171 12257
rect 2314 12248 2320 12300
rect 2372 12288 2378 12300
rect 2961 12291 3019 12297
rect 2961 12288 2973 12291
rect 2372 12260 2973 12288
rect 2372 12248 2378 12260
rect 2961 12257 2973 12260
rect 3007 12257 3019 12291
rect 2961 12251 3019 12257
rect 1762 12180 1768 12232
rect 1820 12220 1826 12232
rect 1857 12223 1915 12229
rect 1857 12220 1869 12223
rect 1820 12192 1869 12220
rect 1820 12180 1826 12192
rect 1857 12189 1869 12192
rect 1903 12189 1915 12223
rect 1857 12183 1915 12189
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 3068 12220 3096 12396
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4212 12396 4261 12424
rect 4212 12384 4218 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4890 12424 4896 12436
rect 4249 12387 4307 12393
rect 4540 12396 4896 12424
rect 4540 12356 4568 12396
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 5166 12384 5172 12436
rect 5224 12424 5230 12436
rect 6270 12424 6276 12436
rect 5224 12396 6276 12424
rect 5224 12384 5230 12396
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 6549 12427 6607 12433
rect 6549 12393 6561 12427
rect 6595 12424 6607 12427
rect 8018 12424 8024 12436
rect 6595 12396 8024 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 8018 12384 8024 12396
rect 8076 12384 8082 12436
rect 8662 12424 8668 12436
rect 8312 12396 8668 12424
rect 3344 12328 4568 12356
rect 4617 12359 4675 12365
rect 2455 12192 3096 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 3142 12180 3148 12232
rect 3200 12180 3206 12232
rect 3344 12229 3372 12328
rect 4172 12300 4200 12328
rect 4617 12325 4629 12359
rect 4663 12356 4675 12359
rect 5534 12356 5540 12368
rect 4663 12328 5540 12356
rect 4663 12325 4675 12328
rect 4617 12319 4675 12325
rect 5534 12316 5540 12328
rect 5592 12316 5598 12368
rect 5626 12316 5632 12368
rect 5684 12356 5690 12368
rect 7190 12356 7196 12368
rect 5684 12328 7196 12356
rect 5684 12316 5690 12328
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 7653 12359 7711 12365
rect 7653 12325 7665 12359
rect 7699 12356 7711 12359
rect 7926 12356 7932 12368
rect 7699 12328 7932 12356
rect 7699 12325 7711 12328
rect 7653 12319 7711 12325
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 8202 12356 8208 12368
rect 8036 12328 8208 12356
rect 4154 12248 4160 12300
rect 4212 12248 4218 12300
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 4304 12260 4752 12288
rect 4304 12248 4310 12260
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3418 12180 3424 12232
rect 3476 12180 3482 12232
rect 4430 12180 4436 12232
rect 4488 12180 4494 12232
rect 4724 12229 4752 12260
rect 5074 12248 5080 12300
rect 5132 12288 5138 12300
rect 5132 12260 5580 12288
rect 5132 12248 5138 12260
rect 5552 12232 5580 12260
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 7282 12288 7288 12300
rect 5960 12260 7288 12288
rect 5960 12248 5966 12260
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4540 12152 4568 12183
rect 4890 12180 4896 12232
rect 4948 12220 4954 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 4948 12192 5457 12220
rect 4948 12180 4954 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 5810 12180 5816 12232
rect 5868 12220 5874 12232
rect 6840 12229 6868 12260
rect 7282 12248 7288 12260
rect 7340 12288 7346 12300
rect 7561 12291 7619 12297
rect 7561 12288 7573 12291
rect 7340 12260 7573 12288
rect 7340 12248 7346 12260
rect 7561 12257 7573 12260
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 6681 12223 6739 12229
rect 6681 12220 6693 12223
rect 5868 12192 6693 12220
rect 5868 12180 5874 12192
rect 6681 12189 6693 12192
rect 6727 12189 6739 12223
rect 6681 12183 6739 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 7101 12223 7159 12229
rect 7101 12220 7113 12223
rect 7064 12192 7113 12220
rect 7064 12180 7070 12192
rect 7101 12189 7113 12192
rect 7147 12189 7159 12223
rect 7929 12223 7987 12229
rect 7101 12183 7159 12189
rect 5166 12152 5172 12164
rect 4540 12124 5172 12152
rect 5166 12112 5172 12124
rect 5224 12112 5230 12164
rect 5261 12155 5319 12161
rect 5261 12121 5273 12155
rect 5307 12121 5319 12155
rect 5261 12115 5319 12121
rect 2222 12044 2228 12096
rect 2280 12044 2286 12096
rect 3878 12044 3884 12096
rect 3936 12084 3942 12096
rect 4246 12084 4252 12096
rect 3936 12056 4252 12084
rect 3936 12044 3942 12056
rect 4246 12044 4252 12056
rect 4304 12084 4310 12096
rect 5276 12084 5304 12115
rect 5350 12112 5356 12164
rect 5408 12152 5414 12164
rect 5629 12155 5687 12161
rect 5629 12152 5641 12155
rect 5408 12124 5641 12152
rect 5408 12112 5414 12124
rect 5629 12121 5641 12124
rect 5675 12121 5687 12155
rect 5629 12115 5687 12121
rect 6270 12112 6276 12164
rect 6328 12152 6334 12164
rect 6917 12155 6975 12161
rect 6328 12124 6868 12152
rect 6328 12112 6334 12124
rect 4304 12056 5304 12084
rect 5813 12087 5871 12093
rect 4304 12044 4310 12056
rect 5813 12053 5825 12087
rect 5859 12084 5871 12087
rect 6730 12084 6736 12096
rect 5859 12056 6736 12084
rect 5859 12053 5871 12056
rect 5813 12047 5871 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 6840 12084 6868 12124
rect 6917 12121 6929 12155
rect 6963 12152 6975 12155
rect 7282 12152 7288 12198
rect 6963 12146 7288 12152
rect 7340 12146 7346 12198
rect 7929 12189 7941 12223
rect 7975 12220 7987 12223
rect 8036 12220 8064 12328
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 8113 12291 8171 12297
rect 8113 12257 8125 12291
rect 8159 12288 8171 12291
rect 8312 12288 8340 12396
rect 8662 12384 8668 12396
rect 8720 12424 8726 12436
rect 9214 12424 9220 12436
rect 8720 12396 9220 12424
rect 8720 12384 8726 12396
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 9309 12427 9367 12433
rect 9309 12393 9321 12427
rect 9355 12424 9367 12427
rect 10410 12424 10416 12436
rect 9355 12396 10416 12424
rect 9355 12393 9367 12396
rect 9309 12387 9367 12393
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 10594 12384 10600 12436
rect 10652 12424 10658 12436
rect 11330 12424 11336 12436
rect 10652 12396 11336 12424
rect 10652 12384 10658 12396
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 11698 12424 11704 12436
rect 11480 12396 11704 12424
rect 11480 12384 11486 12396
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 13446 12424 13452 12436
rect 13096 12396 13452 12424
rect 10042 12316 10048 12368
rect 10100 12356 10106 12368
rect 11238 12356 11244 12368
rect 10100 12328 11244 12356
rect 10100 12316 10106 12328
rect 11238 12316 11244 12328
rect 11296 12316 11302 12368
rect 13096 12356 13124 12396
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 11440 12328 13124 12356
rect 9398 12288 9404 12300
rect 8159 12260 8340 12288
rect 8772 12260 9404 12288
rect 8159 12257 8171 12260
rect 8113 12251 8171 12257
rect 7975 12192 8064 12220
rect 7975 12189 7987 12192
rect 7929 12183 7987 12189
rect 6963 12124 7328 12146
rect 6963 12121 6975 12124
rect 6917 12115 6975 12121
rect 7742 12112 7748 12164
rect 7800 12152 7806 12164
rect 8772 12152 8800 12260
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 9861 12291 9919 12297
rect 9861 12257 9873 12291
rect 9907 12288 9919 12291
rect 10226 12288 10232 12300
rect 9907 12260 10232 12288
rect 9907 12257 9919 12260
rect 9861 12251 9919 12257
rect 10226 12248 10232 12260
rect 10284 12288 10290 12300
rect 10594 12288 10600 12300
rect 10284 12260 10600 12288
rect 10284 12248 10290 12260
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 8938 12180 8944 12232
rect 8996 12220 9002 12232
rect 9565 12223 9623 12229
rect 8996 12192 9444 12220
rect 8996 12180 9002 12192
rect 7800 12124 8800 12152
rect 7800 12112 7806 12124
rect 8846 12112 8852 12164
rect 8904 12152 8910 12164
rect 9309 12155 9367 12161
rect 9309 12152 9321 12155
rect 8904 12124 9321 12152
rect 8904 12112 8910 12124
rect 9309 12121 9321 12124
rect 9355 12121 9367 12155
rect 9309 12115 9367 12121
rect 7282 12084 7288 12096
rect 6840 12056 7288 12084
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 9416 12084 9444 12192
rect 9565 12189 9577 12223
rect 9611 12220 9623 12223
rect 9611 12189 9628 12220
rect 9565 12183 9628 12189
rect 9600 12152 9628 12183
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 9732 12192 10333 12220
rect 9732 12180 9738 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 11440 12220 11468 12328
rect 13354 12316 13360 12368
rect 13412 12356 13418 12368
rect 14277 12359 14335 12365
rect 14277 12356 14289 12359
rect 13412 12328 14289 12356
rect 13412 12316 13418 12328
rect 14277 12325 14289 12328
rect 14323 12356 14335 12359
rect 16022 12356 16028 12368
rect 14323 12328 16028 12356
rect 14323 12325 14335 12328
rect 14277 12319 14335 12325
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 14366 12288 14372 12300
rect 12584 12260 14372 12288
rect 12584 12248 12590 12260
rect 14366 12248 14372 12260
rect 14424 12288 14430 12300
rect 17218 12288 17224 12300
rect 14424 12260 15332 12288
rect 14424 12248 14430 12260
rect 10468 12192 11468 12220
rect 11517 12223 11575 12229
rect 10468 12180 10474 12192
rect 11517 12189 11529 12223
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12220 11667 12223
rect 11882 12220 11888 12232
rect 11655 12192 11888 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 9858 12152 9864 12164
rect 9600 12124 9864 12152
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 10965 12155 11023 12161
rect 10965 12152 10977 12155
rect 10560 12124 10977 12152
rect 10560 12112 10566 12124
rect 10965 12121 10977 12124
rect 11011 12121 11023 12155
rect 11532 12152 11560 12183
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 11974 12180 11980 12232
rect 12032 12220 12038 12232
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 12032 12192 12449 12220
rect 12032 12180 12038 12192
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12710 12180 12716 12232
rect 12768 12180 12774 12232
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12220 14519 12223
rect 14507 12192 15148 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 12618 12152 12624 12164
rect 11532 12124 12624 12152
rect 10965 12115 11023 12121
rect 12618 12112 12624 12124
rect 12676 12112 12682 12164
rect 14645 12155 14703 12161
rect 14645 12121 14657 12155
rect 14691 12152 14703 12155
rect 14826 12152 14832 12164
rect 14691 12124 14832 12152
rect 14691 12121 14703 12124
rect 14645 12115 14703 12121
rect 14826 12112 14832 12124
rect 14884 12112 14890 12164
rect 15120 12152 15148 12192
rect 15194 12180 15200 12232
rect 15252 12180 15258 12232
rect 15304 12229 15332 12260
rect 15948 12260 17224 12288
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12189 15347 12223
rect 15948 12220 15976 12260
rect 17218 12248 17224 12260
rect 17276 12248 17282 12300
rect 15289 12183 15347 12189
rect 15396 12192 15976 12220
rect 16117 12223 16175 12229
rect 15396 12152 15424 12192
rect 16117 12189 16129 12223
rect 16163 12220 16175 12223
rect 16206 12220 16212 12232
rect 16163 12192 16212 12220
rect 16163 12189 16175 12192
rect 16117 12183 16175 12189
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12220 16359 12223
rect 16390 12220 16396 12232
rect 16347 12192 16396 12220
rect 16347 12189 16359 12192
rect 16301 12183 16359 12189
rect 16390 12180 16396 12192
rect 16448 12220 16454 12232
rect 16942 12220 16948 12232
rect 16448 12192 16948 12220
rect 16448 12180 16454 12192
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 17126 12180 17132 12232
rect 17184 12180 17190 12232
rect 15120 12124 15424 12152
rect 15473 12155 15531 12161
rect 15473 12121 15485 12155
rect 15519 12152 15531 12155
rect 15654 12152 15660 12164
rect 15519 12124 15660 12152
rect 15519 12121 15531 12124
rect 15473 12115 15531 12121
rect 15654 12112 15660 12124
rect 15712 12152 15718 12164
rect 16574 12152 16580 12164
rect 15712 12124 16580 12152
rect 15712 12112 15718 12124
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 16758 12112 16764 12164
rect 16816 12152 16822 12164
rect 16853 12155 16911 12161
rect 16853 12152 16865 12155
rect 16816 12124 16865 12152
rect 16816 12112 16822 12124
rect 16853 12121 16865 12124
rect 16899 12121 16911 12155
rect 16853 12115 16911 12121
rect 17310 12112 17316 12164
rect 17368 12152 17374 12164
rect 17681 12155 17739 12161
rect 17681 12152 17693 12155
rect 17368 12124 17693 12152
rect 17368 12112 17374 12124
rect 17681 12121 17693 12124
rect 17727 12121 17739 12155
rect 17681 12115 17739 12121
rect 17862 12112 17868 12164
rect 17920 12112 17926 12164
rect 18049 12155 18107 12161
rect 18049 12121 18061 12155
rect 18095 12152 18107 12155
rect 18782 12152 18788 12164
rect 18095 12124 18788 12152
rect 18095 12121 18107 12124
rect 18049 12115 18107 12121
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 9677 12087 9735 12093
rect 9677 12084 9689 12087
rect 7616 12056 9689 12084
rect 7616 12044 7622 12056
rect 9677 12053 9689 12056
rect 9723 12053 9735 12087
rect 9677 12047 9735 12053
rect 9769 12087 9827 12093
rect 9769 12053 9781 12087
rect 9815 12084 9827 12087
rect 10588 12087 10646 12093
rect 10588 12084 10600 12087
rect 9815 12056 10600 12084
rect 9815 12053 9827 12056
rect 9769 12047 9827 12053
rect 10588 12053 10600 12056
rect 10634 12084 10646 12087
rect 10870 12084 10876 12096
rect 10634 12056 10876 12084
rect 10634 12053 10646 12056
rect 10588 12047 10646 12053
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 11514 12044 11520 12096
rect 11572 12084 11578 12096
rect 11793 12087 11851 12093
rect 11793 12084 11805 12087
rect 11572 12056 11805 12084
rect 11572 12044 11578 12056
rect 11793 12053 11805 12056
rect 11839 12053 11851 12087
rect 11793 12047 11851 12053
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 12986 12084 12992 12096
rect 12492 12056 12992 12084
rect 12492 12044 12498 12056
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 13354 12044 13360 12096
rect 13412 12084 13418 12096
rect 13449 12087 13507 12093
rect 13449 12084 13461 12087
rect 13412 12056 13461 12084
rect 13412 12044 13418 12056
rect 13449 12053 13461 12056
rect 13495 12053 13507 12087
rect 13449 12047 13507 12053
rect 14918 12044 14924 12096
rect 14976 12084 14982 12096
rect 15378 12084 15384 12096
rect 14976 12056 15384 12084
rect 14976 12044 14982 12056
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 16114 12044 16120 12096
rect 16172 12044 16178 12096
rect 1104 11994 18860 12016
rect 1104 11942 5502 11994
rect 5554 11942 5566 11994
rect 5618 11942 5630 11994
rect 5682 11942 5694 11994
rect 5746 11942 5758 11994
rect 5810 11942 5822 11994
rect 5874 11942 5886 11994
rect 5938 11942 5950 11994
rect 6002 11942 6014 11994
rect 6066 11942 6078 11994
rect 6130 11942 6142 11994
rect 6194 11942 6206 11994
rect 6258 11942 6270 11994
rect 6322 11942 6334 11994
rect 6386 11942 6398 11994
rect 6450 11942 6462 11994
rect 6514 11942 6526 11994
rect 6578 11942 6590 11994
rect 6642 11942 6654 11994
rect 6706 11942 13502 11994
rect 13554 11942 13566 11994
rect 13618 11942 13630 11994
rect 13682 11942 13694 11994
rect 13746 11942 13758 11994
rect 13810 11942 13822 11994
rect 13874 11942 13886 11994
rect 13938 11942 13950 11994
rect 14002 11942 14014 11994
rect 14066 11942 14078 11994
rect 14130 11942 14142 11994
rect 14194 11942 14206 11994
rect 14258 11942 14270 11994
rect 14322 11942 14334 11994
rect 14386 11942 14398 11994
rect 14450 11942 14462 11994
rect 14514 11942 14526 11994
rect 14578 11942 14590 11994
rect 14642 11942 14654 11994
rect 14706 11942 18860 11994
rect 1104 11920 18860 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 2317 11883 2375 11889
rect 2317 11880 2329 11883
rect 1452 11852 2329 11880
rect 1452 11840 1458 11852
rect 2317 11849 2329 11852
rect 2363 11849 2375 11883
rect 2317 11843 2375 11849
rect 2685 11883 2743 11889
rect 2685 11849 2697 11883
rect 2731 11880 2743 11883
rect 2731 11852 3096 11880
rect 2731 11849 2743 11852
rect 2685 11843 2743 11849
rect 2406 11772 2412 11824
rect 2464 11812 2470 11824
rect 2501 11815 2559 11821
rect 2501 11812 2513 11815
rect 2464 11784 2513 11812
rect 2464 11772 2470 11784
rect 2501 11781 2513 11784
rect 2547 11781 2559 11815
rect 2501 11775 2559 11781
rect 2590 11772 2596 11824
rect 2648 11772 2654 11824
rect 2866 11772 2872 11824
rect 2924 11772 2930 11824
rect 3068 11812 3096 11852
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 3878 11880 3884 11892
rect 3200 11852 3884 11880
rect 3200 11840 3206 11852
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 4614 11840 4620 11892
rect 4672 11880 4678 11892
rect 5169 11883 5227 11889
rect 5169 11880 5181 11883
rect 4672 11852 5181 11880
rect 4672 11840 4678 11852
rect 5169 11849 5181 11852
rect 5215 11849 5227 11883
rect 10042 11880 10048 11892
rect 5169 11843 5227 11849
rect 6564 11852 8156 11880
rect 3068 11784 3372 11812
rect 3344 11744 3372 11784
rect 3418 11772 3424 11824
rect 3476 11812 3482 11824
rect 6362 11812 6368 11824
rect 3476 11784 6368 11812
rect 3476 11772 3482 11784
rect 3786 11744 3792 11756
rect 3344 11716 3792 11744
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 4131 11747 4189 11753
rect 4131 11713 4143 11747
rect 4177 11744 4189 11747
rect 4246 11744 4252 11756
rect 4177 11716 4252 11744
rect 4177 11713 4189 11716
rect 4131 11707 4189 11713
rect 3988 11676 4016 11707
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 4356 11753 4384 11784
rect 5184 11756 5212 11784
rect 6362 11772 6368 11784
rect 6420 11772 6426 11824
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11744 4675 11747
rect 4663 11716 4752 11744
rect 4663 11713 4675 11716
rect 4617 11707 4675 11713
rect 4430 11676 4436 11688
rect 3988 11648 4436 11676
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 3510 11568 3516 11620
rect 3568 11608 3574 11620
rect 4724 11608 4752 11716
rect 4798 11704 4804 11756
rect 4856 11704 4862 11756
rect 5166 11704 5172 11756
rect 5224 11704 5230 11756
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 5353 11747 5411 11753
rect 5353 11744 5365 11747
rect 5316 11716 5365 11744
rect 5316 11704 5322 11716
rect 5353 11713 5365 11716
rect 5399 11744 5411 11747
rect 5399 11716 5580 11744
rect 5399 11713 5411 11716
rect 5353 11707 5411 11713
rect 4816 11676 4844 11704
rect 5445 11679 5503 11685
rect 5445 11676 5457 11679
rect 4816 11648 5457 11676
rect 5445 11645 5457 11648
rect 5491 11645 5503 11679
rect 5552 11676 5580 11716
rect 5626 11704 5632 11756
rect 5684 11704 5690 11756
rect 5810 11704 5816 11756
rect 5868 11704 5874 11756
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6564 11753 6592 11852
rect 7190 11812 7196 11824
rect 6840 11784 7196 11812
rect 6840 11753 6868 11784
rect 7190 11772 7196 11784
rect 7248 11772 7254 11824
rect 7834 11812 7840 11824
rect 7668 11784 7840 11812
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 5960 11716 6561 11744
rect 5960 11704 5966 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 5920 11676 5948 11704
rect 5552 11648 5948 11676
rect 5445 11639 5503 11645
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 6641 11679 6699 11685
rect 6641 11676 6653 11679
rect 6052 11648 6653 11676
rect 6052 11636 6058 11648
rect 6641 11645 6653 11648
rect 6687 11645 6699 11679
rect 7116 11676 7144 11707
rect 7558 11704 7564 11756
rect 7616 11704 7622 11756
rect 7190 11676 7196 11688
rect 7116 11648 7196 11676
rect 6641 11639 6699 11645
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 5258 11608 5264 11620
rect 3568 11580 4660 11608
rect 4724 11580 5264 11608
rect 3568 11568 3574 11580
rect 4632 11552 4660 11580
rect 5258 11568 5264 11580
rect 5316 11568 5322 11620
rect 5537 11611 5595 11617
rect 5537 11577 5549 11611
rect 5583 11608 5595 11611
rect 5583 11580 5617 11608
rect 5583 11577 5595 11580
rect 5537 11571 5595 11577
rect 1302 11500 1308 11552
rect 1360 11540 1366 11552
rect 1762 11540 1768 11552
rect 1360 11512 1768 11540
rect 1360 11500 1366 11512
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4028 11512 4353 11540
rect 4028 11500 4034 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 5552 11540 5580 11571
rect 6454 11568 6460 11620
rect 6512 11608 6518 11620
rect 7006 11608 7012 11620
rect 6512 11580 7012 11608
rect 6512 11568 6518 11580
rect 7006 11568 7012 11580
rect 7064 11568 7070 11620
rect 7576 11540 7604 11704
rect 7668 11552 7696 11784
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11713 8079 11747
rect 8128 11744 8156 11852
rect 8588 11852 10048 11880
rect 8389 11815 8447 11821
rect 8389 11781 8401 11815
rect 8435 11812 8447 11815
rect 8588 11812 8616 11852
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10244 11852 10456 11880
rect 9674 11812 9680 11824
rect 8435 11784 8616 11812
rect 8864 11784 9680 11812
rect 8435 11781 8447 11784
rect 8389 11775 8447 11781
rect 8128 11716 8524 11744
rect 8021 11707 8079 11713
rect 8036 11608 8064 11707
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11645 8171 11679
rect 8113 11639 8171 11645
rect 7760 11580 8064 11608
rect 8128 11608 8156 11639
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8496 11685 8524 11716
rect 8864 11740 8892 11784
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 9766 11772 9772 11824
rect 9824 11812 9830 11824
rect 10244 11812 10272 11852
rect 10428 11821 10456 11852
rect 10502 11840 10508 11892
rect 10560 11880 10566 11892
rect 11606 11880 11612 11892
rect 10560 11852 11612 11880
rect 10560 11840 10566 11852
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 12986 11880 12992 11892
rect 12452 11852 12992 11880
rect 9824 11784 10272 11812
rect 10413 11815 10471 11821
rect 9824 11772 9830 11784
rect 10413 11781 10425 11815
rect 10459 11781 10471 11815
rect 10413 11775 10471 11781
rect 10778 11772 10784 11824
rect 10836 11812 10842 11824
rect 11882 11812 11888 11824
rect 10836 11784 11888 11812
rect 10836 11772 10842 11784
rect 11882 11772 11888 11784
rect 11940 11812 11946 11824
rect 12452 11821 12480 11852
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13725 11883 13783 11889
rect 13725 11880 13737 11883
rect 13412 11852 13737 11880
rect 13412 11840 13418 11852
rect 13725 11849 13737 11852
rect 13771 11849 13783 11883
rect 13725 11843 13783 11849
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 14826 11880 14832 11892
rect 14608 11852 14832 11880
rect 14608 11840 14614 11852
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 12437 11815 12495 11821
rect 11940 11784 12297 11812
rect 11940 11772 11946 11784
rect 8941 11747 8999 11753
rect 8941 11740 8953 11747
rect 8864 11713 8953 11740
rect 8987 11713 8999 11747
rect 8864 11712 8999 11713
rect 8941 11707 8999 11712
rect 9398 11704 9404 11756
rect 9456 11744 9462 11756
rect 9493 11747 9551 11753
rect 9493 11744 9505 11747
rect 9456 11716 9505 11744
rect 9456 11704 9462 11716
rect 9493 11713 9505 11716
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 8297 11679 8355 11685
rect 8297 11676 8309 11679
rect 8260 11648 8309 11676
rect 8260 11636 8266 11648
rect 8297 11645 8309 11648
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 8481 11679 8539 11685
rect 8481 11645 8493 11679
rect 8527 11676 8539 11679
rect 9309 11679 9367 11685
rect 8527 11648 9168 11676
rect 8527 11645 8539 11648
rect 8481 11639 8539 11645
rect 8570 11608 8576 11620
rect 8128 11580 8576 11608
rect 7760 11552 7788 11580
rect 8570 11568 8576 11580
rect 8628 11568 8634 11620
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9033 11611 9091 11617
rect 9033 11608 9045 11611
rect 8996 11580 9045 11608
rect 8996 11568 9002 11580
rect 9033 11577 9045 11580
rect 9079 11577 9091 11611
rect 9140 11608 9168 11648
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 9582 11676 9588 11688
rect 9355 11648 9588 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 9766 11636 9772 11688
rect 9824 11636 9830 11688
rect 10244 11676 10272 11707
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 10686 11753 10692 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10376 11716 10517 11744
rect 10376 11704 10382 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 10649 11747 10692 11753
rect 10649 11713 10661 11747
rect 10744 11744 10750 11756
rect 12269 11753 12297 11784
rect 12437 11781 12449 11815
rect 12483 11781 12495 11815
rect 13170 11812 13176 11824
rect 12437 11775 12495 11781
rect 12544 11784 13176 11812
rect 12544 11753 12572 11784
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 13262 11772 13268 11824
rect 13320 11812 13326 11824
rect 13633 11815 13691 11821
rect 13633 11812 13645 11815
rect 13320 11784 13645 11812
rect 13320 11772 13326 11784
rect 13633 11781 13645 11784
rect 13679 11781 13691 11815
rect 15378 11812 15384 11824
rect 13633 11775 13691 11781
rect 14936 11784 15384 11812
rect 12710 11753 12716 11756
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 10744 11716 12173 11744
rect 10649 11707 10692 11713
rect 10686 11704 10692 11707
rect 10744 11704 10750 11716
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 12254 11747 12312 11753
rect 12254 11713 12266 11747
rect 12300 11713 12312 11747
rect 12254 11707 12312 11713
rect 12529 11747 12587 11753
rect 12529 11713 12541 11747
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 12667 11747 12716 11753
rect 12667 11713 12679 11747
rect 12713 11713 12716 11747
rect 12667 11707 12716 11713
rect 10870 11676 10876 11688
rect 10244 11648 10876 11676
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 12176 11676 12204 11707
rect 12710 11704 12716 11707
rect 12768 11704 12774 11756
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 13280 11744 13308 11772
rect 14936 11753 14964 11784
rect 15378 11772 15384 11784
rect 15436 11812 15442 11824
rect 17957 11815 18015 11821
rect 15436 11784 15700 11812
rect 15436 11772 15442 11784
rect 13044 11716 13308 11744
rect 14737 11747 14795 11753
rect 13044 11704 13050 11716
rect 14737 11713 14749 11747
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 13449 11679 13507 11685
rect 12176 11648 12572 11676
rect 12544 11620 12572 11648
rect 13449 11645 13461 11679
rect 13495 11645 13507 11679
rect 14752 11676 14780 11707
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15672 11753 15700 11784
rect 17957 11781 17969 11815
rect 18003 11812 18015 11815
rect 18966 11812 18972 11824
rect 18003 11784 18972 11812
rect 18003 11781 18015 11784
rect 17957 11775 18015 11781
rect 18966 11772 18972 11784
rect 19024 11772 19030 11824
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11744 15715 11747
rect 16206 11744 16212 11756
rect 15703 11716 16212 11744
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 16942 11704 16948 11756
rect 17000 11704 17006 11756
rect 17126 11704 17132 11756
rect 17184 11704 17190 11756
rect 17402 11704 17408 11756
rect 17460 11744 17466 11756
rect 18141 11747 18199 11753
rect 18141 11744 18153 11747
rect 17460 11716 18153 11744
rect 17460 11704 17466 11716
rect 18141 11713 18153 11716
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 15194 11676 15200 11688
rect 14752 11648 15200 11676
rect 13449 11639 13507 11645
rect 9140 11580 12480 11608
rect 9033 11571 9091 11577
rect 4672 11512 7604 11540
rect 4672 11500 4678 11512
rect 7650 11500 7656 11552
rect 7708 11500 7714 11552
rect 7742 11500 7748 11552
rect 7800 11500 7806 11552
rect 7837 11543 7895 11549
rect 7837 11509 7849 11543
rect 7883 11540 7895 11543
rect 9398 11540 9404 11552
rect 7883 11512 9404 11540
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 10781 11543 10839 11549
rect 10781 11509 10793 11543
rect 10827 11540 10839 11543
rect 11146 11540 11152 11552
rect 10827 11512 11152 11540
rect 10827 11509 10839 11512
rect 10781 11503 10839 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 12452 11540 12480 11580
rect 12526 11568 12532 11620
rect 12584 11608 12590 11620
rect 13464 11608 13492 11639
rect 15194 11636 15200 11648
rect 15252 11676 15258 11688
rect 15488 11676 15516 11704
rect 15252 11648 15516 11676
rect 15252 11636 15258 11648
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 16853 11679 16911 11685
rect 16853 11676 16865 11679
rect 16540 11648 16865 11676
rect 16540 11636 16546 11648
rect 16853 11645 16865 11648
rect 16899 11645 16911 11679
rect 16853 11639 16911 11645
rect 14274 11608 14280 11620
rect 12584 11580 14280 11608
rect 12584 11568 12590 11580
rect 14274 11568 14280 11580
rect 14332 11568 14338 11620
rect 14645 11611 14703 11617
rect 14645 11577 14657 11611
rect 14691 11608 14703 11611
rect 14826 11608 14832 11620
rect 14691 11580 14832 11608
rect 14691 11577 14703 11580
rect 14645 11571 14703 11577
rect 14826 11568 14832 11580
rect 14884 11568 14890 11620
rect 15473 11611 15531 11617
rect 15473 11577 15485 11611
rect 15519 11608 15531 11611
rect 15562 11608 15568 11620
rect 15519 11580 15568 11608
rect 15519 11577 15531 11580
rect 15473 11571 15531 11577
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 15838 11568 15844 11620
rect 15896 11608 15902 11620
rect 17773 11611 17831 11617
rect 17773 11608 17785 11611
rect 15896 11580 17785 11608
rect 15896 11568 15902 11580
rect 17773 11577 17785 11580
rect 17819 11577 17831 11611
rect 17773 11571 17831 11577
rect 12710 11540 12716 11552
rect 12452 11512 12716 11540
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 12802 11500 12808 11552
rect 12860 11500 12866 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 14093 11543 14151 11549
rect 14093 11540 14105 11543
rect 13320 11512 14105 11540
rect 13320 11500 13326 11512
rect 14093 11509 14105 11512
rect 14139 11509 14151 11543
rect 14093 11503 14151 11509
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 17862 11540 17868 11552
rect 16632 11512 17868 11540
rect 16632 11500 16638 11512
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 1104 11450 18860 11472
rect 1104 11398 1502 11450
rect 1554 11398 1566 11450
rect 1618 11398 1630 11450
rect 1682 11398 1694 11450
rect 1746 11398 1758 11450
rect 1810 11398 1822 11450
rect 1874 11398 1886 11450
rect 1938 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 2270 11450
rect 2322 11398 2334 11450
rect 2386 11398 2398 11450
rect 2450 11398 2462 11450
rect 2514 11398 2526 11450
rect 2578 11398 2590 11450
rect 2642 11398 2654 11450
rect 2706 11398 9502 11450
rect 9554 11398 9566 11450
rect 9618 11398 9630 11450
rect 9682 11398 9694 11450
rect 9746 11398 9758 11450
rect 9810 11398 9822 11450
rect 9874 11398 9886 11450
rect 9938 11398 9950 11450
rect 10002 11398 10014 11450
rect 10066 11398 10078 11450
rect 10130 11398 10142 11450
rect 10194 11398 10206 11450
rect 10258 11398 10270 11450
rect 10322 11398 10334 11450
rect 10386 11398 10398 11450
rect 10450 11398 10462 11450
rect 10514 11398 10526 11450
rect 10578 11398 10590 11450
rect 10642 11398 10654 11450
rect 10706 11398 17502 11450
rect 17554 11398 17566 11450
rect 17618 11398 17630 11450
rect 17682 11398 17694 11450
rect 17746 11398 17758 11450
rect 17810 11398 17822 11450
rect 17874 11398 17886 11450
rect 17938 11398 17950 11450
rect 18002 11398 18014 11450
rect 18066 11398 18078 11450
rect 18130 11398 18142 11450
rect 18194 11398 18206 11450
rect 18258 11398 18270 11450
rect 18322 11398 18334 11450
rect 18386 11398 18398 11450
rect 18450 11398 18462 11450
rect 18514 11398 18526 11450
rect 18578 11398 18590 11450
rect 18642 11398 18654 11450
rect 18706 11398 18860 11450
rect 1104 11376 18860 11398
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 3418 11336 3424 11348
rect 1820 11308 3424 11336
rect 1820 11296 1826 11308
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 7374 11336 7380 11348
rect 7064 11308 7380 11336
rect 7064 11296 7070 11308
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 9122 11336 9128 11348
rect 8260 11308 9128 11336
rect 8260 11296 8266 11308
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 9214 11296 9220 11348
rect 9272 11336 9278 11348
rect 9490 11336 9496 11348
rect 9272 11308 9496 11336
rect 9272 11296 9278 11308
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 11885 11339 11943 11345
rect 11885 11336 11897 11339
rect 10796 11308 11897 11336
rect 3973 11271 4031 11277
rect 3973 11268 3985 11271
rect 2792 11240 3985 11268
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 2792 11209 2820 11240
rect 3973 11237 3985 11240
rect 4019 11237 4031 11271
rect 3973 11231 4031 11237
rect 4430 11228 4436 11280
rect 4488 11268 4494 11280
rect 4798 11268 4804 11280
rect 4488 11240 4804 11268
rect 4488 11228 4494 11240
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 5166 11228 5172 11280
rect 5224 11228 5230 11280
rect 5902 11228 5908 11280
rect 5960 11228 5966 11280
rect 6454 11268 6460 11280
rect 6012 11240 6460 11268
rect 2481 11203 2539 11209
rect 2481 11200 2493 11203
rect 1452 11172 2493 11200
rect 1452 11160 1458 11172
rect 2481 11169 2493 11172
rect 2527 11169 2539 11203
rect 2481 11163 2539 11169
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11169 2835 11203
rect 2777 11163 2835 11169
rect 4614 11160 4620 11212
rect 4672 11160 4678 11212
rect 6012 11200 6040 11240
rect 6454 11228 6460 11240
rect 6512 11228 6518 11280
rect 7190 11228 7196 11280
rect 7248 11268 7254 11280
rect 7926 11268 7932 11280
rect 7248 11240 7932 11268
rect 7248 11228 7254 11240
rect 7926 11228 7932 11240
rect 7984 11228 7990 11280
rect 10796 11277 10824 11308
rect 11885 11305 11897 11308
rect 11931 11336 11943 11339
rect 12066 11336 12072 11348
rect 11931 11308 12072 11336
rect 11931 11305 11943 11308
rect 11885 11299 11943 11305
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 14274 11296 14280 11348
rect 14332 11296 14338 11348
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 15654 11336 15660 11348
rect 15528 11308 15660 11336
rect 15528 11296 15534 11308
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 10781 11271 10839 11277
rect 10781 11237 10793 11271
rect 10827 11237 10839 11271
rect 10781 11231 10839 11237
rect 10873 11271 10931 11277
rect 10873 11237 10885 11271
rect 10919 11268 10931 11271
rect 10919 11240 12297 11268
rect 10919 11237 10931 11240
rect 10873 11231 10931 11237
rect 4724 11172 6040 11200
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2866 11132 2872 11144
rect 2087 11104 2872 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4341 11135 4399 11141
rect 4341 11132 4353 11135
rect 4120 11104 4353 11132
rect 4120 11092 4126 11104
rect 4341 11101 4353 11104
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11132 4491 11135
rect 4724 11132 4752 11172
rect 4479 11104 4752 11132
rect 4479 11101 4491 11104
rect 4433 11095 4491 11101
rect 4798 11092 4804 11144
rect 4856 11132 4862 11144
rect 5169 11135 5227 11141
rect 5169 11132 5181 11135
rect 4856 11104 5181 11132
rect 4856 11092 4862 11104
rect 5169 11101 5181 11104
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 7208 11132 7236 11228
rect 7742 11160 7748 11212
rect 7800 11200 7806 11212
rect 8113 11203 8171 11209
rect 7800 11172 8064 11200
rect 7800 11160 7806 11172
rect 6503 11104 7236 11132
rect 7929 11135 7987 11141
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 8036 11132 8064 11172
rect 8113 11169 8125 11203
rect 8159 11200 8171 11203
rect 8570 11200 8576 11212
rect 8159 11172 8576 11200
rect 8159 11169 8171 11172
rect 8113 11163 8171 11169
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 9950 11160 9956 11212
rect 10008 11160 10014 11212
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10686 11200 10692 11212
rect 10459 11172 10692 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 11054 11200 11060 11212
rect 10980 11172 11060 11200
rect 8846 11132 8852 11144
rect 8036 11104 8852 11132
rect 7929 11095 7987 11101
rect 1302 11024 1308 11076
rect 1360 11064 1366 11076
rect 2222 11064 2228 11076
rect 1360 11036 2228 11064
rect 1360 11024 1366 11036
rect 2222 11024 2228 11036
rect 2280 11024 2286 11076
rect 2685 11067 2743 11073
rect 2685 11033 2697 11067
rect 2731 11064 2743 11067
rect 2731 11036 4292 11064
rect 2731 11033 2743 11036
rect 2685 11027 2743 11033
rect 2593 10999 2651 11005
rect 2593 10965 2605 10999
rect 2639 10996 2651 10999
rect 3602 10996 3608 11008
rect 2639 10968 3608 10996
rect 2639 10965 2651 10968
rect 2593 10959 2651 10965
rect 3602 10956 3608 10968
rect 3660 10956 3666 11008
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 4154 10996 4160 11008
rect 4028 10968 4160 10996
rect 4028 10956 4034 10968
rect 4154 10956 4160 10968
rect 4212 10956 4218 11008
rect 4264 10996 4292 11036
rect 4614 11024 4620 11076
rect 4672 11064 4678 11076
rect 6104 11064 6132 11095
rect 4672 11036 6132 11064
rect 4672 11024 4678 11036
rect 6362 11024 6368 11076
rect 6420 11064 6426 11076
rect 6733 11067 6791 11073
rect 6733 11064 6745 11067
rect 6420 11036 6745 11064
rect 6420 11024 6426 11036
rect 6733 11033 6745 11036
rect 6779 11064 6791 11067
rect 7558 11064 7564 11076
rect 6779 11036 7564 11064
rect 6779 11033 6791 11036
rect 6733 11027 6791 11033
rect 7558 11024 7564 11036
rect 7616 11064 7622 11076
rect 7944 11064 7972 11095
rect 8846 11092 8852 11104
rect 8904 11092 8910 11144
rect 9214 11092 9220 11144
rect 9272 11092 9278 11144
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 9858 11132 9864 11144
rect 9815 11104 9864 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 7616 11036 7972 11064
rect 7616 11024 7622 11036
rect 4706 10996 4712 11008
rect 4264 10968 4712 10996
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 7193 10999 7251 11005
rect 7193 10965 7205 10999
rect 7239 10996 7251 10999
rect 7374 10996 7380 11008
rect 7239 10968 7380 10996
rect 7239 10965 7251 10968
rect 7193 10959 7251 10965
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 7944 10996 7972 11036
rect 8018 11024 8024 11076
rect 8076 11064 8082 11076
rect 9401 11067 9459 11073
rect 8076 11036 8984 11064
rect 8076 11024 8082 11036
rect 8956 11008 8984 11036
rect 9401 11033 9413 11067
rect 9447 11064 9459 11067
rect 9490 11064 9496 11076
rect 9447 11036 9496 11064
rect 9447 11033 9459 11036
rect 9401 11027 9459 11033
rect 9490 11024 9496 11036
rect 9548 11024 9554 11076
rect 10686 11024 10692 11076
rect 10744 11064 10750 11076
rect 10980 11064 11008 11172
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 12269 11200 12297 11240
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 14645 11271 14703 11277
rect 14645 11268 14657 11271
rect 12400 11240 14657 11268
rect 12400 11228 12406 11240
rect 14645 11237 14657 11240
rect 14691 11237 14703 11271
rect 14645 11231 14703 11237
rect 12269 11172 14320 11200
rect 11514 11092 11520 11144
rect 11572 11092 11578 11144
rect 11977 11135 12035 11141
rect 11977 11101 11989 11135
rect 12023 11132 12035 11135
rect 12158 11132 12164 11144
rect 12023 11104 12164 11132
rect 12023 11101 12035 11104
rect 11977 11095 12035 11101
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 14292 11141 14320 11172
rect 14458 11160 14464 11212
rect 14516 11200 14522 11212
rect 15197 11203 15255 11209
rect 15197 11200 15209 11203
rect 14516 11172 15209 11200
rect 14516 11160 14522 11172
rect 15197 11169 15209 11172
rect 15243 11169 15255 11203
rect 15197 11163 15255 11169
rect 17126 11160 17132 11212
rect 17184 11200 17190 11212
rect 17184 11172 17540 11200
rect 17184 11160 17190 11172
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12268 11104 12725 11132
rect 10744 11036 11008 11064
rect 10744 11024 10750 11036
rect 11606 11024 11612 11076
rect 11664 11064 11670 11076
rect 12268 11064 12296 11104
rect 12713 11101 12725 11104
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11101 12955 11135
rect 12897 11095 12955 11101
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 12912 11064 12940 11095
rect 11664 11036 12296 11064
rect 12728 11036 12940 11064
rect 11664 11024 11670 11036
rect 12728 11008 12756 11036
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 14384 11064 14412 11095
rect 14642 11092 14648 11144
rect 14700 11132 14706 11144
rect 15102 11132 15108 11144
rect 14700 11104 15108 11132
rect 14700 11092 14706 11104
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 13228 11036 14412 11064
rect 13228 11024 13234 11036
rect 14550 11024 14556 11076
rect 14608 11064 14614 11076
rect 14608 11036 15148 11064
rect 14608 11024 14614 11036
rect 8110 10996 8116 11008
rect 7944 10968 8116 10996
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 8938 10956 8944 11008
rect 8996 10956 9002 11008
rect 9030 10956 9036 11008
rect 9088 10996 9094 11008
rect 9309 10999 9367 11005
rect 9309 10996 9321 10999
rect 9088 10968 9321 10996
rect 9088 10956 9094 10968
rect 9309 10965 9321 10968
rect 9355 10965 9367 10999
rect 9309 10959 9367 10965
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 11882 10996 11888 11008
rect 9824 10968 11888 10996
rect 9824 10956 9830 10968
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 12710 10956 12716 11008
rect 12768 10956 12774 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13725 10999 13783 11005
rect 13725 10996 13737 10999
rect 13412 10968 13737 10996
rect 13412 10956 13418 10968
rect 13725 10965 13737 10968
rect 13771 10965 13783 10999
rect 15120 10996 15148 11036
rect 15194 11024 15200 11076
rect 15252 11064 15258 11076
rect 15304 11064 15332 11095
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 15473 11135 15531 11141
rect 15473 11132 15485 11135
rect 15436 11104 15485 11132
rect 15436 11092 15442 11104
rect 15473 11101 15485 11104
rect 15519 11132 15531 11135
rect 16393 11135 16451 11141
rect 16393 11132 16405 11135
rect 15519 11104 16405 11132
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 16393 11101 16405 11104
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 16942 11132 16948 11144
rect 16715 11104 16948 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 16942 11092 16948 11104
rect 17000 11132 17006 11144
rect 17512 11141 17540 11172
rect 17313 11135 17371 11141
rect 17313 11132 17325 11135
rect 17000 11104 17325 11132
rect 17000 11092 17006 11104
rect 17313 11101 17325 11104
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 17497 11135 17555 11141
rect 17497 11101 17509 11135
rect 17543 11101 17555 11135
rect 17497 11095 17555 11101
rect 15252 11036 15332 11064
rect 16761 11067 16819 11073
rect 15252 11024 15258 11036
rect 16761 11033 16773 11067
rect 16807 11064 16819 11067
rect 16850 11064 16856 11076
rect 16807 11036 16856 11064
rect 16807 11033 16819 11036
rect 16761 11027 16819 11033
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 17034 11024 17040 11076
rect 17092 11064 17098 11076
rect 17221 11067 17279 11073
rect 17221 11064 17233 11067
rect 17092 11036 17233 11064
rect 17092 11024 17098 11036
rect 17221 11033 17233 11036
rect 17267 11033 17279 11067
rect 17221 11027 17279 11033
rect 17126 10996 17132 11008
rect 15120 10968 17132 10996
rect 13725 10959 13783 10965
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 1104 10906 18860 10928
rect 1104 10854 5502 10906
rect 5554 10854 5566 10906
rect 5618 10854 5630 10906
rect 5682 10854 5694 10906
rect 5746 10854 5758 10906
rect 5810 10854 5822 10906
rect 5874 10854 5886 10906
rect 5938 10854 5950 10906
rect 6002 10854 6014 10906
rect 6066 10854 6078 10906
rect 6130 10854 6142 10906
rect 6194 10854 6206 10906
rect 6258 10854 6270 10906
rect 6322 10854 6334 10906
rect 6386 10854 6398 10906
rect 6450 10854 6462 10906
rect 6514 10854 6526 10906
rect 6578 10854 6590 10906
rect 6642 10854 6654 10906
rect 6706 10854 13502 10906
rect 13554 10854 13566 10906
rect 13618 10854 13630 10906
rect 13682 10854 13694 10906
rect 13746 10854 13758 10906
rect 13810 10854 13822 10906
rect 13874 10854 13886 10906
rect 13938 10854 13950 10906
rect 14002 10854 14014 10906
rect 14066 10854 14078 10906
rect 14130 10854 14142 10906
rect 14194 10854 14206 10906
rect 14258 10854 14270 10906
rect 14322 10854 14334 10906
rect 14386 10854 14398 10906
rect 14450 10854 14462 10906
rect 14514 10854 14526 10906
rect 14578 10854 14590 10906
rect 14642 10854 14654 10906
rect 14706 10854 18860 10906
rect 1104 10832 18860 10854
rect 1118 10752 1124 10804
rect 1176 10792 1182 10804
rect 2961 10795 3019 10801
rect 2961 10792 2973 10795
rect 1176 10764 2973 10792
rect 1176 10752 1182 10764
rect 2961 10761 2973 10764
rect 3007 10761 3019 10795
rect 2961 10755 3019 10761
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 3970 10792 3976 10804
rect 3099 10764 3976 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 290 10684 296 10736
rect 348 10724 354 10736
rect 348 10696 2084 10724
rect 348 10684 354 10696
rect 1762 10616 1768 10668
rect 1820 10616 1826 10668
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10625 2007 10659
rect 2056 10656 2084 10696
rect 2222 10684 2228 10736
rect 2280 10724 2286 10736
rect 2593 10727 2651 10733
rect 2593 10724 2605 10727
rect 2280 10696 2605 10724
rect 2280 10684 2286 10696
rect 2593 10693 2605 10696
rect 2639 10693 2651 10727
rect 2976 10724 3004 10755
rect 3970 10752 3976 10764
rect 4028 10792 4034 10804
rect 4157 10795 4215 10801
rect 4157 10792 4169 10795
rect 4028 10764 4169 10792
rect 4028 10752 4034 10764
rect 4157 10761 4169 10764
rect 4203 10761 4215 10795
rect 4157 10755 4215 10761
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 4890 10792 4896 10804
rect 4672 10764 4896 10792
rect 4672 10752 4678 10764
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5445 10795 5503 10801
rect 5445 10761 5457 10795
rect 5491 10792 5503 10795
rect 7466 10792 7472 10804
rect 5491 10764 7472 10792
rect 5491 10761 5503 10764
rect 5445 10755 5503 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8168 10764 8861 10792
rect 8168 10752 8174 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 2976 10696 3096 10724
rect 2593 10687 2651 10693
rect 2823 10659 2881 10665
rect 2823 10656 2835 10659
rect 2056 10628 2835 10656
rect 1949 10619 2007 10625
rect 2823 10625 2835 10628
rect 2869 10625 2881 10659
rect 2823 10619 2881 10625
rect 1964 10588 1992 10619
rect 1964 10560 2524 10588
rect 1854 10480 1860 10532
rect 1912 10480 1918 10532
rect 1394 10412 1400 10464
rect 1452 10452 1458 10464
rect 2409 10455 2467 10461
rect 2409 10452 2421 10455
rect 1452 10424 2421 10452
rect 1452 10412 1458 10424
rect 2409 10421 2421 10424
rect 2455 10421 2467 10455
rect 2496 10452 2524 10560
rect 3068 10520 3096 10696
rect 3602 10684 3608 10736
rect 3660 10724 3666 10736
rect 4522 10724 4528 10736
rect 3660 10696 4528 10724
rect 3660 10684 3666 10696
rect 4522 10684 4528 10696
rect 4580 10724 4586 10736
rect 5353 10727 5411 10733
rect 5353 10724 5365 10727
rect 4580 10696 5365 10724
rect 4580 10684 4586 10696
rect 5353 10693 5365 10696
rect 5399 10693 5411 10727
rect 8864 10724 8892 10755
rect 9214 10752 9220 10804
rect 9272 10792 9278 10804
rect 9674 10792 9680 10804
rect 9272 10764 9680 10792
rect 9272 10752 9278 10764
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 14829 10795 14887 10801
rect 14829 10792 14841 10795
rect 9784 10764 14841 10792
rect 9582 10724 9588 10736
rect 8864 10696 9588 10724
rect 5353 10687 5411 10693
rect 9582 10684 9588 10696
rect 9640 10684 9646 10736
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3476 10628 3709 10656
rect 3476 10616 3482 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3844 10628 3985 10656
rect 3844 10616 3850 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4706 10616 4712 10668
rect 4764 10656 4770 10668
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 4764 10628 5273 10656
rect 4764 10616 4770 10628
rect 5261 10625 5273 10628
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5500 10628 5825 10656
rect 5500 10616 5506 10628
rect 5813 10625 5825 10628
rect 5859 10625 5871 10659
rect 9784 10656 9812 10764
rect 14829 10761 14841 10764
rect 14875 10761 14887 10795
rect 14829 10755 14887 10761
rect 17957 10795 18015 10801
rect 17957 10761 17969 10795
rect 18003 10792 18015 10795
rect 19242 10792 19248 10804
rect 18003 10764 19248 10792
rect 18003 10761 18015 10764
rect 17957 10755 18015 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 10965 10727 11023 10733
rect 10965 10693 10977 10727
rect 11011 10724 11023 10727
rect 11330 10724 11336 10736
rect 11011 10696 11336 10724
rect 11011 10693 11023 10696
rect 10965 10687 11023 10693
rect 11330 10684 11336 10696
rect 11388 10684 11394 10736
rect 11514 10684 11520 10736
rect 11572 10724 11578 10736
rect 12066 10724 12072 10736
rect 11572 10696 12072 10724
rect 11572 10684 11578 10696
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 15194 10724 15200 10736
rect 14936 10696 15200 10724
rect 12342 10665 12348 10668
rect 8510 10628 9812 10656
rect 12311 10659 12348 10665
rect 5813 10619 5871 10625
rect 3145 10591 3203 10597
rect 3145 10557 3157 10591
rect 3191 10588 3203 10591
rect 3878 10588 3884 10600
rect 3191 10560 3884 10588
rect 3191 10557 3203 10560
rect 3145 10551 3203 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 4338 10588 4344 10600
rect 4295 10560 4344 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 4338 10548 4344 10560
rect 4396 10588 4402 10600
rect 4982 10588 4988 10600
rect 4396 10560 4988 10588
rect 4396 10548 4402 10560
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 5534 10548 5540 10600
rect 5592 10597 5598 10600
rect 5592 10591 5611 10597
rect 5599 10557 5611 10591
rect 5592 10551 5611 10557
rect 5592 10548 5598 10551
rect 7098 10548 7104 10600
rect 7156 10597 7162 10600
rect 7156 10551 7166 10597
rect 7156 10548 7162 10551
rect 8662 10548 8668 10600
rect 8720 10588 8726 10600
rect 8846 10588 8852 10600
rect 8720 10560 8852 10588
rect 8720 10548 8726 10560
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9306 10548 9312 10600
rect 9364 10588 9370 10600
rect 10060 10588 10088 10642
rect 12311 10625 12323 10659
rect 12311 10619 12348 10625
rect 12342 10616 12348 10619
rect 12400 10616 12406 10668
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 12713 10659 12771 10665
rect 12713 10656 12725 10659
rect 12584 10628 12725 10656
rect 12584 10616 12590 10628
rect 12713 10625 12725 10628
rect 12759 10625 12771 10659
rect 12713 10619 12771 10625
rect 12802 10616 12808 10668
rect 12860 10656 12866 10668
rect 14936 10665 14964 10696
rect 15194 10684 15200 10696
rect 15252 10684 15258 10736
rect 15396 10696 15884 10724
rect 15396 10668 15424 10696
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 12860 10628 13461 10656
rect 12860 10616 12866 10628
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10656 15163 10659
rect 15378 10656 15384 10668
rect 15151 10628 15384 10656
rect 15151 10625 15163 10628
rect 15105 10619 15163 10625
rect 9364 10560 10088 10588
rect 10137 10591 10195 10597
rect 9364 10548 9370 10560
rect 10137 10557 10149 10591
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 6546 10520 6552 10532
rect 3068 10492 6552 10520
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 9950 10480 9956 10532
rect 10008 10520 10014 10532
rect 10152 10520 10180 10551
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 12158 10588 12164 10600
rect 10928 10560 12164 10588
rect 10928 10548 10934 10560
rect 12158 10548 12164 10560
rect 12216 10548 12222 10600
rect 12618 10548 12624 10600
rect 12676 10548 12682 10600
rect 13354 10548 13360 10600
rect 13412 10548 13418 10600
rect 14274 10548 14280 10600
rect 14332 10548 14338 10600
rect 14458 10548 14464 10600
rect 14516 10588 14522 10600
rect 14936 10588 14964 10619
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 15856 10665 15884 10696
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10656 15899 10659
rect 16206 10656 16212 10668
rect 15887 10628 16212 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 15672 10588 15700 10619
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 16390 10616 16396 10668
rect 16448 10656 16454 10668
rect 17957 10659 18015 10665
rect 17957 10656 17969 10659
rect 16448 10628 17969 10656
rect 16448 10616 16454 10628
rect 17957 10625 17969 10628
rect 18003 10625 18015 10659
rect 17957 10619 18015 10625
rect 14516 10560 15700 10588
rect 14516 10548 14522 10560
rect 16942 10548 16948 10600
rect 17000 10588 17006 10600
rect 17218 10588 17224 10600
rect 17000 10560 17224 10588
rect 17000 10548 17006 10560
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 17402 10548 17408 10600
rect 17460 10588 17466 10600
rect 17589 10591 17647 10597
rect 17589 10588 17601 10591
rect 17460 10560 17601 10588
rect 17460 10548 17466 10560
rect 17589 10557 17601 10560
rect 17635 10557 17647 10591
rect 17589 10551 17647 10557
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10588 18199 10591
rect 18874 10588 18880 10600
rect 18187 10560 18880 10588
rect 18187 10557 18199 10560
rect 18141 10551 18199 10557
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 11422 10520 11428 10532
rect 10008 10492 11428 10520
rect 10008 10480 10014 10492
rect 11422 10480 11428 10492
rect 11480 10480 11486 10532
rect 11882 10480 11888 10532
rect 11940 10520 11946 10532
rect 12069 10523 12127 10529
rect 12069 10520 12081 10523
rect 11940 10492 12081 10520
rect 11940 10480 11946 10492
rect 12069 10489 12081 10492
rect 12115 10489 12127 10523
rect 12636 10520 12664 10548
rect 12636 10492 13400 10520
rect 12069 10483 12127 10489
rect 13372 10464 13400 10492
rect 15654 10480 15660 10532
rect 15712 10480 15718 10532
rect 3142 10452 3148 10464
rect 2496 10424 3148 10452
rect 2409 10415 2467 10421
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3881 10455 3939 10461
rect 3881 10421 3893 10455
rect 3927 10452 3939 10455
rect 3970 10452 3976 10464
rect 3927 10424 3976 10452
rect 3927 10421 3939 10424
rect 3881 10415 3939 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 5258 10452 5264 10464
rect 4479 10424 5264 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 6822 10452 6828 10464
rect 6043 10424 6828 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7374 10461 7380 10464
rect 7364 10455 7380 10461
rect 7364 10421 7376 10455
rect 7364 10415 7380 10421
rect 7374 10412 7380 10415
rect 7432 10412 7438 10464
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 8478 10452 8484 10464
rect 7984 10424 8484 10452
rect 7984 10412 7990 10424
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 9766 10452 9772 10464
rect 8720 10424 9772 10452
rect 8720 10412 8726 10424
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 12618 10452 12624 10464
rect 10192 10424 12624 10452
rect 10192 10412 10198 10424
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 13354 10412 13360 10464
rect 13412 10412 13418 10464
rect 15010 10412 15016 10464
rect 15068 10452 15074 10464
rect 16022 10452 16028 10464
rect 15068 10424 16028 10452
rect 15068 10412 15074 10424
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 17218 10452 17224 10464
rect 16356 10424 17224 10452
rect 16356 10412 16362 10424
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 1104 10362 18860 10384
rect 1104 10310 1502 10362
rect 1554 10310 1566 10362
rect 1618 10310 1630 10362
rect 1682 10310 1694 10362
rect 1746 10310 1758 10362
rect 1810 10310 1822 10362
rect 1874 10310 1886 10362
rect 1938 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 2270 10362
rect 2322 10310 2334 10362
rect 2386 10310 2398 10362
rect 2450 10310 2462 10362
rect 2514 10310 2526 10362
rect 2578 10310 2590 10362
rect 2642 10310 2654 10362
rect 2706 10310 9502 10362
rect 9554 10310 9566 10362
rect 9618 10310 9630 10362
rect 9682 10310 9694 10362
rect 9746 10310 9758 10362
rect 9810 10310 9822 10362
rect 9874 10310 9886 10362
rect 9938 10310 9950 10362
rect 10002 10310 10014 10362
rect 10066 10310 10078 10362
rect 10130 10310 10142 10362
rect 10194 10310 10206 10362
rect 10258 10310 10270 10362
rect 10322 10310 10334 10362
rect 10386 10310 10398 10362
rect 10450 10310 10462 10362
rect 10514 10310 10526 10362
rect 10578 10310 10590 10362
rect 10642 10310 10654 10362
rect 10706 10310 17502 10362
rect 17554 10310 17566 10362
rect 17618 10310 17630 10362
rect 17682 10310 17694 10362
rect 17746 10310 17758 10362
rect 17810 10310 17822 10362
rect 17874 10310 17886 10362
rect 17938 10310 17950 10362
rect 18002 10310 18014 10362
rect 18066 10310 18078 10362
rect 18130 10310 18142 10362
rect 18194 10310 18206 10362
rect 18258 10310 18270 10362
rect 18322 10310 18334 10362
rect 18386 10310 18398 10362
rect 18450 10310 18462 10362
rect 18514 10310 18526 10362
rect 18578 10310 18590 10362
rect 18642 10310 18654 10362
rect 18706 10310 18860 10362
rect 1104 10288 18860 10310
rect 2590 10208 2596 10260
rect 2648 10248 2654 10260
rect 2866 10248 2872 10260
rect 2648 10220 2872 10248
rect 2648 10208 2654 10220
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 4890 10248 4896 10260
rect 3200 10220 4896 10248
rect 3200 10208 3206 10220
rect 4890 10208 4896 10220
rect 4948 10208 4954 10260
rect 4982 10208 4988 10260
rect 5040 10248 5046 10260
rect 10502 10248 10508 10260
rect 5040 10220 10508 10248
rect 5040 10208 5046 10220
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 12158 10248 12164 10260
rect 10888 10220 12164 10248
rect 3326 10140 3332 10192
rect 3384 10180 3390 10192
rect 10137 10183 10195 10189
rect 3384 10152 5580 10180
rect 3384 10140 3390 10152
rect 2314 10112 2320 10124
rect 1596 10084 2320 10112
rect 1596 10053 1624 10084
rect 2314 10072 2320 10084
rect 2372 10112 2378 10124
rect 2372 10084 4108 10112
rect 2372 10072 2378 10084
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10044 2191 10047
rect 2866 10044 2872 10056
rect 2179 10016 2872 10044
rect 2179 10013 2191 10016
rect 2133 10007 2191 10013
rect 2866 10004 2872 10016
rect 2924 10044 2930 10056
rect 3142 10044 3148 10056
rect 2924 10016 3148 10044
rect 2924 10004 2930 10016
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 3326 10044 3332 10056
rect 3283 10016 3332 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 4080 10053 4108 10084
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 5442 10044 5448 10056
rect 4764 10016 5448 10044
rect 4764 10004 4770 10016
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5552 10053 5580 10152
rect 10137 10149 10149 10183
rect 10183 10180 10195 10183
rect 10888 10180 10916 10220
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 14642 10208 14648 10260
rect 14700 10248 14706 10260
rect 16298 10248 16304 10260
rect 14700 10220 16304 10248
rect 14700 10208 14706 10220
rect 16298 10208 16304 10220
rect 16356 10208 16362 10260
rect 17126 10208 17132 10260
rect 17184 10248 17190 10260
rect 17494 10248 17500 10260
rect 17184 10220 17500 10248
rect 17184 10208 17190 10220
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 10183 10152 10916 10180
rect 11164 10152 13124 10180
rect 10183 10149 10195 10152
rect 10137 10143 10195 10149
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7745 10115 7803 10121
rect 7745 10112 7757 10115
rect 6972 10084 7757 10112
rect 6972 10072 6978 10084
rect 7745 10081 7757 10084
rect 7791 10081 7803 10115
rect 8570 10112 8576 10124
rect 7745 10075 7803 10081
rect 7852 10084 8576 10112
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10044 6423 10047
rect 7282 10044 7288 10056
rect 6411 10016 7288 10044
rect 6411 10013 6423 10016
rect 6365 10007 6423 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 1026 9936 1032 9988
rect 1084 9936 1090 9988
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 2406 9976 2412 9988
rect 1719 9948 2412 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 2406 9936 2412 9948
rect 2464 9936 2470 9988
rect 2682 9936 2688 9988
rect 2740 9936 2746 9988
rect 2777 9979 2835 9985
rect 2777 9945 2789 9979
rect 2823 9976 2835 9979
rect 3973 9979 4031 9985
rect 3973 9976 3985 9979
rect 2823 9948 3985 9976
rect 2823 9945 2835 9948
rect 2777 9939 2835 9945
rect 3973 9945 3985 9948
rect 4019 9976 4031 9979
rect 6549 9979 6607 9985
rect 6549 9976 6561 9979
rect 4019 9948 6561 9976
rect 4019 9945 4031 9948
rect 3973 9939 4031 9945
rect 6549 9945 6561 9948
rect 6595 9976 6607 9979
rect 7852 9976 7880 10084
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 9122 10072 9128 10124
rect 9180 10112 9186 10124
rect 11164 10112 11192 10152
rect 9180 10084 11192 10112
rect 13096 10112 13124 10152
rect 17218 10140 17224 10192
rect 17276 10180 17282 10192
rect 18690 10180 18696 10192
rect 17276 10152 18696 10180
rect 17276 10140 17282 10152
rect 18690 10140 18696 10152
rect 18748 10140 18754 10192
rect 15010 10112 15016 10124
rect 13096 10084 15016 10112
rect 9180 10072 9186 10084
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 8220 10016 9321 10044
rect 6595 9948 7880 9976
rect 6595 9945 6607 9948
rect 6549 9939 6607 9945
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 8220 9985 8248 10016
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 9766 10004 9772 10056
rect 9824 10004 9830 10056
rect 10704 10053 10732 10084
rect 11336 10056 11388 10062
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 12526 10004 12532 10056
rect 12584 10044 12590 10056
rect 13096 10053 13124 10084
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 15378 10112 15384 10124
rect 15120 10084 15384 10112
rect 12713 10047 12771 10053
rect 12713 10044 12725 10047
rect 12584 10016 12725 10044
rect 12584 10004 12590 10016
rect 12713 10013 12725 10016
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10013 13139 10047
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13081 10007 13139 10013
rect 13188 10016 14289 10044
rect 11336 9998 11388 10004
rect 8205 9979 8263 9985
rect 8205 9976 8217 9979
rect 8168 9948 8217 9976
rect 8168 9936 8174 9948
rect 8205 9945 8217 9948
rect 8251 9945 8263 9979
rect 8205 9939 8263 9945
rect 8297 9979 8355 9985
rect 8297 9945 8309 9979
rect 8343 9945 8355 9979
rect 8297 9939 8355 9945
rect 1044 9908 1072 9936
rect 1210 9908 1216 9920
rect 1044 9880 1216 9908
rect 1210 9868 1216 9880
rect 1268 9868 1274 9920
rect 4982 9868 4988 9920
rect 5040 9908 5046 9920
rect 6638 9908 6644 9920
rect 5040 9880 6644 9908
rect 5040 9868 5046 9880
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 7101 9911 7159 9917
rect 7101 9877 7113 9911
rect 7147 9908 7159 9911
rect 8312 9908 8340 9939
rect 9122 9936 9128 9988
rect 9180 9936 9186 9988
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9945 10011 9979
rect 9953 9939 10011 9945
rect 7147 9880 8340 9908
rect 9968 9908 9996 9939
rect 10870 9936 10876 9988
rect 10928 9976 10934 9988
rect 11238 9976 11244 9988
rect 10928 9948 11244 9976
rect 10928 9936 10934 9948
rect 11238 9936 11244 9948
rect 11296 9936 11302 9988
rect 11698 9936 11704 9988
rect 11756 9936 11762 9988
rect 12066 9936 12072 9988
rect 12124 9976 12130 9988
rect 13188 9976 13216 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14458 10004 14464 10056
rect 14516 10004 14522 10056
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10044 14703 10047
rect 15120 10044 15148 10084
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15749 10115 15807 10121
rect 15749 10081 15761 10115
rect 15795 10112 15807 10115
rect 17126 10112 17132 10124
rect 15795 10084 17132 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 18095 10115 18153 10121
rect 18095 10081 18107 10115
rect 18141 10112 18153 10115
rect 18782 10112 18788 10124
rect 18141 10084 18788 10112
rect 18141 10081 18153 10084
rect 18095 10075 18153 10081
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 14691 10016 15148 10044
rect 14691 10013 14703 10016
rect 14645 10007 14703 10013
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 15252 10016 15485 10044
rect 15252 10004 15258 10016
rect 15473 10013 15485 10016
rect 15519 10013 15531 10047
rect 17957 10047 18015 10053
rect 17957 10044 17969 10047
rect 15473 10007 15531 10013
rect 17144 10016 17969 10044
rect 17034 9976 17040 9988
rect 12124 9948 13216 9976
rect 16974 9948 17040 9976
rect 12124 9936 12130 9948
rect 17034 9936 17040 9948
rect 17092 9936 17098 9988
rect 11054 9908 11060 9920
rect 9968 9880 11060 9908
rect 7147 9877 7159 9880
rect 7101 9871 7159 9877
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 13262 9868 13268 9920
rect 13320 9908 13326 9920
rect 13725 9911 13783 9917
rect 13725 9908 13737 9911
rect 13320 9880 13737 9908
rect 13320 9868 13326 9880
rect 13725 9877 13737 9880
rect 13771 9877 13783 9911
rect 13725 9871 13783 9877
rect 14826 9868 14832 9920
rect 14884 9908 14890 9920
rect 15286 9908 15292 9920
rect 14884 9880 15292 9908
rect 14884 9868 14890 9880
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 15930 9868 15936 9920
rect 15988 9908 15994 9920
rect 16390 9908 16396 9920
rect 15988 9880 16396 9908
rect 15988 9868 15994 9880
rect 16390 9868 16396 9880
rect 16448 9908 16454 9920
rect 17144 9908 17172 10016
rect 17957 10013 17969 10016
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 17402 9936 17408 9988
rect 17460 9976 17466 9988
rect 18340 9976 18368 10007
rect 18782 9976 18788 9988
rect 17460 9948 18788 9976
rect 17460 9936 17466 9948
rect 18782 9936 18788 9948
rect 18840 9936 18846 9988
rect 16448 9880 17172 9908
rect 16448 9868 16454 9880
rect 17218 9868 17224 9920
rect 17276 9868 17282 9920
rect 17957 9911 18015 9917
rect 17957 9877 17969 9911
rect 18003 9908 18015 9911
rect 18046 9908 18052 9920
rect 18003 9880 18052 9908
rect 18003 9877 18015 9880
rect 17957 9871 18015 9877
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 290 9800 296 9852
rect 348 9840 354 9852
rect 842 9840 848 9852
rect 348 9812 848 9840
rect 348 9800 354 9812
rect 842 9800 848 9812
rect 900 9800 906 9852
rect 1104 9818 18860 9840
rect 1104 9766 5502 9818
rect 5554 9766 5566 9818
rect 5618 9766 5630 9818
rect 5682 9766 5694 9818
rect 5746 9766 5758 9818
rect 5810 9766 5822 9818
rect 5874 9766 5886 9818
rect 5938 9766 5950 9818
rect 6002 9766 6014 9818
rect 6066 9766 6078 9818
rect 6130 9766 6142 9818
rect 6194 9766 6206 9818
rect 6258 9766 6270 9818
rect 6322 9766 6334 9818
rect 6386 9766 6398 9818
rect 6450 9766 6462 9818
rect 6514 9766 6526 9818
rect 6578 9766 6590 9818
rect 6642 9766 6654 9818
rect 6706 9766 13502 9818
rect 13554 9766 13566 9818
rect 13618 9766 13630 9818
rect 13682 9766 13694 9818
rect 13746 9766 13758 9818
rect 13810 9766 13822 9818
rect 13874 9766 13886 9818
rect 13938 9766 13950 9818
rect 14002 9766 14014 9818
rect 14066 9766 14078 9818
rect 14130 9766 14142 9818
rect 14194 9766 14206 9818
rect 14258 9766 14270 9818
rect 14322 9766 14334 9818
rect 14386 9766 14398 9818
rect 14450 9766 14462 9818
rect 14514 9766 14526 9818
rect 14578 9766 14590 9818
rect 14642 9766 14654 9818
rect 14706 9766 18860 9818
rect 1104 9744 18860 9766
rect 106 9664 112 9716
rect 164 9704 170 9716
rect 3970 9704 3976 9716
rect 164 9676 3976 9704
rect 164 9664 170 9676
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 5074 9664 5080 9716
rect 5132 9704 5138 9716
rect 5261 9707 5319 9713
rect 5261 9704 5273 9707
rect 5132 9676 5273 9704
rect 5132 9664 5138 9676
rect 5261 9673 5273 9676
rect 5307 9673 5319 9707
rect 5261 9667 5319 9673
rect 5350 9664 5356 9716
rect 5408 9664 5414 9716
rect 6914 9704 6920 9716
rect 6564 9676 6920 9704
rect 2682 9596 2688 9648
rect 2740 9636 2746 9648
rect 4157 9639 4215 9645
rect 4157 9636 4169 9639
rect 2740 9608 4169 9636
rect 2740 9596 2746 9608
rect 4157 9605 4169 9608
rect 4203 9605 4215 9639
rect 4157 9599 4215 9605
rect 4522 9596 4528 9648
rect 4580 9636 4586 9648
rect 4706 9636 4712 9648
rect 4580 9608 4712 9636
rect 4580 9596 4586 9608
rect 4706 9596 4712 9608
rect 4764 9636 4770 9648
rect 4893 9639 4951 9645
rect 4893 9636 4905 9639
rect 4764 9608 4905 9636
rect 4764 9596 4770 9608
rect 4893 9605 4905 9608
rect 4939 9605 4951 9639
rect 4893 9599 4951 9605
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 2314 9568 2320 9580
rect 1903 9540 2320 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 566 9460 572 9512
rect 624 9500 630 9512
rect 1026 9500 1032 9512
rect 624 9472 1032 9500
rect 624 9460 630 9472
rect 1026 9460 1032 9472
rect 1084 9460 1090 9512
rect 1688 9500 1716 9531
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 2464 9540 3065 9568
rect 2464 9528 2470 9540
rect 3053 9537 3065 9540
rect 3099 9568 3111 9571
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3099 9540 4077 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 6564 9577 6592 9676
rect 6914 9664 6920 9676
rect 6972 9664 6978 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 11330 9704 11336 9716
rect 10836 9676 11336 9704
rect 10836 9664 10842 9676
rect 11330 9664 11336 9676
rect 11388 9664 11394 9716
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 12069 9707 12127 9713
rect 12069 9704 12081 9707
rect 11756 9676 12081 9704
rect 11756 9664 11762 9676
rect 12069 9673 12081 9676
rect 12115 9673 12127 9707
rect 12069 9667 12127 9673
rect 12158 9664 12164 9716
rect 12216 9664 12222 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 12768 9676 14964 9704
rect 12768 9664 12774 9676
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 8110 9636 8116 9648
rect 7055 9608 8116 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 8110 9596 8116 9608
rect 8168 9596 8174 9648
rect 8205 9639 8263 9645
rect 8205 9605 8217 9639
rect 8251 9636 8263 9639
rect 9122 9636 9128 9648
rect 8251 9608 9128 9636
rect 8251 9605 8263 9608
rect 8205 9599 8263 9605
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 10502 9596 10508 9648
rect 10560 9636 10566 9648
rect 12176 9636 12204 9664
rect 10560 9608 12204 9636
rect 10560 9596 10566 9608
rect 12342 9596 12348 9648
rect 12400 9636 12406 9648
rect 12986 9636 12992 9648
rect 12400 9608 12992 9636
rect 12400 9596 12406 9608
rect 12986 9596 12992 9608
rect 13044 9636 13050 9648
rect 13449 9639 13507 9645
rect 13449 9636 13461 9639
rect 13044 9608 13461 9636
rect 13044 9596 13050 9608
rect 13449 9605 13461 9608
rect 13495 9605 13507 9639
rect 13449 9599 13507 9605
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 5316 9540 5457 9568
rect 5316 9528 5322 9540
rect 5445 9537 5457 9540
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9568 7159 9571
rect 7282 9568 7288 9580
rect 7147 9540 7288 9568
rect 7147 9537 7159 9540
rect 7101 9531 7159 9537
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 7668 9540 8953 9568
rect 2774 9500 2780 9512
rect 1688 9472 2780 9500
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9469 3019 9503
rect 2961 9463 3019 9469
rect 2501 9435 2559 9441
rect 2501 9401 2513 9435
rect 2547 9432 2559 9435
rect 2976 9432 3004 9463
rect 3142 9460 3148 9512
rect 3200 9500 3206 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 3200 9472 3525 9500
rect 3200 9460 3206 9472
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 5152 9503 5210 9509
rect 5152 9469 5164 9503
rect 5198 9500 5210 9503
rect 5350 9500 5356 9512
rect 5198 9472 5356 9500
rect 5198 9469 5210 9472
rect 5152 9463 5210 9469
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7668 9509 7696 9540
rect 8941 9537 8953 9540
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 6972 9472 7665 9500
rect 6972 9460 6978 9472
rect 7653 9469 7665 9472
rect 7699 9469 7711 9503
rect 7653 9463 7711 9469
rect 8018 9460 8024 9512
rect 8076 9500 8082 9512
rect 9876 9500 9904 9531
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11480 9540 11989 9568
rect 11480 9528 11486 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 12526 9568 12532 9580
rect 11977 9531 12035 9537
rect 12360 9540 12532 9568
rect 8076 9472 9904 9500
rect 11885 9503 11943 9509
rect 8076 9460 8082 9472
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 12360 9500 12388 9540
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 14093 9571 14151 9577
rect 14093 9568 14105 9571
rect 12676 9540 14105 9568
rect 12676 9528 12682 9540
rect 14093 9537 14105 9540
rect 14139 9537 14151 9571
rect 14093 9531 14151 9537
rect 14303 9571 14361 9577
rect 14303 9537 14315 9571
rect 14349 9568 14361 9571
rect 14826 9568 14832 9580
rect 14349 9540 14832 9568
rect 14349 9537 14361 9540
rect 14303 9531 14361 9537
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 11931 9472 12388 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 12434 9460 12440 9512
rect 12492 9460 12498 9512
rect 14458 9500 14464 9512
rect 13280 9472 14464 9500
rect 2547 9404 3004 9432
rect 2547 9401 2559 9404
rect 2501 9395 2559 9401
rect 6546 9392 6552 9444
rect 6604 9432 6610 9444
rect 8113 9435 8171 9441
rect 8113 9432 8125 9435
rect 6604 9404 8125 9432
rect 6604 9392 6610 9404
rect 8113 9401 8125 9404
rect 8159 9432 8171 9435
rect 10229 9435 10287 9441
rect 10229 9432 10241 9435
rect 8159 9404 10241 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 10229 9401 10241 9404
rect 10275 9401 10287 9435
rect 10229 9395 10287 9401
rect 10686 9392 10692 9444
rect 10744 9432 10750 9444
rect 11054 9432 11060 9444
rect 10744 9404 11060 9432
rect 10744 9392 10750 9404
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 12452 9432 12480 9460
rect 12989 9435 13047 9441
rect 12989 9432 13001 9435
rect 11756 9404 13001 9432
rect 11756 9392 11762 9404
rect 12989 9401 13001 9404
rect 13035 9401 13047 9435
rect 12989 9395 13047 9401
rect 13170 9392 13176 9444
rect 13228 9392 13234 9444
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 3142 9364 3148 9376
rect 2648 9336 3148 9364
rect 2648 9324 2654 9336
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 4706 9324 4712 9376
rect 4764 9324 4770 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 8018 9364 8024 9376
rect 7340 9336 8024 9364
rect 7340 9324 7346 9336
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 12342 9324 12348 9376
rect 12400 9364 12406 9376
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 12400 9336 12449 9364
rect 12400 9324 12406 9336
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12437 9327 12495 9333
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 13280 9364 13308 9472
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 14936 9500 14964 9676
rect 15102 9664 15108 9716
rect 15160 9664 15166 9716
rect 15120 9636 15148 9664
rect 15028 9608 15148 9636
rect 15028 9577 15056 9608
rect 17310 9596 17316 9648
rect 17368 9596 17374 9648
rect 19334 9636 19340 9648
rect 17420 9608 19340 9636
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15933 9571 15991 9577
rect 15933 9568 15945 9571
rect 15105 9531 15163 9537
rect 15764 9540 15945 9568
rect 15120 9500 15148 9531
rect 15764 9512 15792 9540
rect 15933 9537 15945 9540
rect 15979 9537 15991 9571
rect 15933 9531 15991 9537
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9537 16175 9571
rect 16117 9531 16175 9537
rect 14936 9472 15148 9500
rect 15746 9460 15752 9512
rect 15804 9460 15810 9512
rect 15841 9503 15899 9509
rect 15841 9469 15853 9503
rect 15887 9469 15899 9503
rect 15841 9463 15899 9469
rect 13538 9392 13544 9444
rect 13596 9432 13602 9444
rect 13596 9404 14044 9432
rect 13596 9392 13602 9404
rect 14016 9373 14044 9404
rect 14182 9392 14188 9444
rect 14240 9432 14246 9444
rect 15856 9432 15884 9463
rect 14240 9404 15884 9432
rect 15948 9432 15976 9531
rect 16132 9500 16160 9531
rect 16206 9528 16212 9580
rect 16264 9528 16270 9580
rect 16666 9528 16672 9580
rect 16724 9528 16730 9580
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17420 9568 17448 9608
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 17083 9540 17448 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17494 9528 17500 9580
rect 17552 9568 17558 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17552 9540 17877 9568
rect 17552 9528 17558 9540
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 16224 9500 16252 9528
rect 16390 9500 16396 9512
rect 16132 9472 16396 9500
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 16684 9500 16712 9528
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16684 9472 16865 9500
rect 16853 9469 16865 9472
rect 16899 9500 16911 9503
rect 16942 9500 16948 9512
rect 16899 9472 16948 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17405 9503 17463 9509
rect 17405 9469 17417 9503
rect 17451 9500 17463 9503
rect 18064 9500 18092 9531
rect 17451 9472 18092 9500
rect 17451 9469 17463 9472
rect 17405 9463 17463 9469
rect 16666 9432 16672 9444
rect 15948 9404 16672 9432
rect 14240 9392 14246 9404
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 17034 9392 17040 9444
rect 17092 9432 17098 9444
rect 17420 9432 17448 9463
rect 17092 9404 17448 9432
rect 17092 9392 17098 9404
rect 17954 9392 17960 9444
rect 18012 9392 18018 9444
rect 12860 9336 13308 9364
rect 14001 9367 14059 9373
rect 12860 9324 12866 9336
rect 14001 9333 14013 9367
rect 14047 9333 14059 9367
rect 14001 9327 14059 9333
rect 14090 9324 14096 9376
rect 14148 9364 14154 9376
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 14148 9336 15301 9364
rect 14148 9324 14154 9336
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 15289 9327 15347 9333
rect 15746 9324 15752 9376
rect 15804 9364 15810 9376
rect 18046 9364 18052 9376
rect 15804 9336 18052 9364
rect 15804 9324 15810 9336
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 1104 9274 18860 9296
rect 1104 9222 1502 9274
rect 1554 9222 1566 9274
rect 1618 9222 1630 9274
rect 1682 9222 1694 9274
rect 1746 9222 1758 9274
rect 1810 9222 1822 9274
rect 1874 9222 1886 9274
rect 1938 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 2270 9274
rect 2322 9222 2334 9274
rect 2386 9222 2398 9274
rect 2450 9222 2462 9274
rect 2514 9222 2526 9274
rect 2578 9222 2590 9274
rect 2642 9222 2654 9274
rect 2706 9222 9502 9274
rect 9554 9222 9566 9274
rect 9618 9222 9630 9274
rect 9682 9222 9694 9274
rect 9746 9222 9758 9274
rect 9810 9222 9822 9274
rect 9874 9222 9886 9274
rect 9938 9222 9950 9274
rect 10002 9222 10014 9274
rect 10066 9222 10078 9274
rect 10130 9222 10142 9274
rect 10194 9222 10206 9274
rect 10258 9222 10270 9274
rect 10322 9222 10334 9274
rect 10386 9222 10398 9274
rect 10450 9222 10462 9274
rect 10514 9222 10526 9274
rect 10578 9222 10590 9274
rect 10642 9222 10654 9274
rect 10706 9222 17502 9274
rect 17554 9222 17566 9274
rect 17618 9222 17630 9274
rect 17682 9222 17694 9274
rect 17746 9222 17758 9274
rect 17810 9222 17822 9274
rect 17874 9222 17886 9274
rect 17938 9222 17950 9274
rect 18002 9222 18014 9274
rect 18066 9222 18078 9274
rect 18130 9222 18142 9274
rect 18194 9222 18206 9274
rect 18258 9222 18270 9274
rect 18322 9222 18334 9274
rect 18386 9222 18398 9274
rect 18450 9222 18462 9274
rect 18514 9222 18526 9274
rect 18578 9222 18590 9274
rect 18642 9222 18654 9274
rect 18706 9222 18860 9274
rect 1104 9200 18860 9222
rect 5258 9120 5264 9172
rect 5316 9160 5322 9172
rect 9950 9160 9956 9172
rect 5316 9132 9956 9160
rect 5316 9120 5322 9132
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 12526 9160 12532 9172
rect 12400 9132 12532 9160
rect 12400 9120 12406 9132
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 15102 9160 15108 9172
rect 13044 9132 15108 9160
rect 13044 9120 13050 9132
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17497 9163 17555 9169
rect 17497 9160 17509 9163
rect 17184 9132 17509 9160
rect 17184 9120 17190 9132
rect 17497 9129 17509 9132
rect 17543 9129 17555 9163
rect 17497 9123 17555 9129
rect 3050 9052 3056 9104
rect 3108 9092 3114 9104
rect 3108 9064 5580 9092
rect 3108 9052 3114 9064
rect 2866 9024 2872 9036
rect 1596 8996 2872 9024
rect 1596 8965 1624 8996
rect 2866 8984 2872 8996
rect 2924 9024 2930 9036
rect 2924 8996 4108 9024
rect 2924 8984 2930 8996
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 2958 8956 2964 8968
rect 2179 8928 2964 8956
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 4080 8965 4108 8996
rect 5552 8965 5580 9064
rect 7742 9052 7748 9104
rect 7800 9052 7806 9104
rect 13170 9052 13176 9104
rect 13228 9092 13234 9104
rect 13357 9095 13415 9101
rect 13357 9092 13369 9095
rect 13228 9064 13369 9092
rect 13228 9052 13234 9064
rect 13357 9061 13369 9064
rect 13403 9092 13415 9095
rect 13446 9092 13452 9104
rect 13403 9064 13452 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 7760 9024 7788 9052
rect 5644 8996 7788 9024
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3108 8928 3249 8956
rect 3108 8916 3114 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 1673 8891 1731 8897
rect 1673 8857 1685 8891
rect 1719 8888 1731 8891
rect 2222 8888 2228 8900
rect 1719 8860 2228 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 2222 8848 2228 8860
rect 2280 8848 2286 8900
rect 2682 8848 2688 8900
rect 2740 8848 2746 8900
rect 2774 8848 2780 8900
rect 2832 8888 2838 8900
rect 3973 8891 4031 8897
rect 3973 8888 3985 8891
rect 2832 8860 3985 8888
rect 2832 8848 2838 8860
rect 3973 8857 3985 8860
rect 4019 8857 4031 8891
rect 3973 8851 4031 8857
rect 4430 8848 4436 8900
rect 4488 8888 4494 8900
rect 5258 8888 5264 8900
rect 4488 8860 5264 8888
rect 4488 8848 4494 8860
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 5644 8820 5672 8996
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9769 9027 9827 9033
rect 9769 9024 9781 9027
rect 9548 8996 9781 9024
rect 9548 8984 9554 8996
rect 9769 8993 9781 8996
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 9024 9919 9027
rect 10686 9024 10692 9036
rect 9907 8996 10692 9024
rect 9907 8993 9919 8996
rect 9861 8987 9919 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 11609 9027 11667 9033
rect 11609 8993 11621 9027
rect 11655 9024 11667 9027
rect 14277 9027 14335 9033
rect 14277 9024 14289 9027
rect 11655 8996 14289 9024
rect 11655 8993 11667 8996
rect 11609 8987 11667 8993
rect 14277 8993 14289 8996
rect 14323 9024 14335 9027
rect 15194 9024 15200 9036
rect 14323 8996 15200 9024
rect 14323 8993 14335 8996
rect 14277 8987 14335 8993
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 7282 8916 7288 8968
rect 7340 8916 7346 8968
rect 7742 8916 7748 8968
rect 7800 8916 7806 8968
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 8220 8928 9321 8956
rect 6365 8891 6423 8897
rect 6365 8857 6377 8891
rect 6411 8888 6423 8891
rect 7300 8888 7328 8916
rect 6411 8860 7328 8888
rect 6411 8857 6423 8860
rect 6365 8851 6423 8857
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 8220 8897 8248 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 10228 8959 10286 8965
rect 10228 8925 10240 8959
rect 10274 8956 10286 8959
rect 11054 8956 11060 8968
rect 10274 8928 11060 8956
rect 10274 8925 10286 8928
rect 10228 8919 10286 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11624 8956 11652 8987
rect 15194 8984 15200 8996
rect 15252 8984 15258 9036
rect 17678 9024 17684 9036
rect 16684 8996 17684 9024
rect 16684 8968 16712 8996
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 18046 8984 18052 9036
rect 18104 8984 18110 9036
rect 14182 8956 14188 8968
rect 11195 8928 11652 8956
rect 13018 8928 14188 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 15654 8916 15660 8968
rect 15712 8916 15718 8968
rect 16666 8916 16672 8968
rect 16724 8916 16730 8968
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 8205 8891 8263 8897
rect 8205 8888 8217 8891
rect 8168 8860 8217 8888
rect 8168 8848 8174 8860
rect 8205 8857 8217 8860
rect 8251 8857 8263 8891
rect 8205 8851 8263 8857
rect 8297 8891 8355 8897
rect 8297 8857 8309 8891
rect 8343 8857 8355 8891
rect 8297 8851 8355 8857
rect 10413 8891 10471 8897
rect 10413 8857 10425 8891
rect 10459 8888 10471 8891
rect 10459 8860 11100 8888
rect 10459 8857 10471 8860
rect 10413 8851 10471 8857
rect 3384 8792 5672 8820
rect 7101 8823 7159 8829
rect 3384 8780 3390 8792
rect 7101 8789 7113 8823
rect 7147 8820 7159 8823
rect 8312 8820 8340 8851
rect 11072 8832 11100 8860
rect 11882 8848 11888 8900
rect 11940 8848 11946 8900
rect 13170 8848 13176 8900
rect 13228 8888 13234 8900
rect 14090 8888 14096 8900
rect 13228 8860 14096 8888
rect 13228 8848 13234 8860
rect 14090 8848 14096 8860
rect 14148 8848 14154 8900
rect 14553 8891 14611 8897
rect 14553 8857 14565 8891
rect 14599 8888 14611 8891
rect 14642 8888 14648 8900
rect 14599 8860 14648 8888
rect 14599 8857 14611 8860
rect 14553 8851 14611 8857
rect 14642 8848 14648 8860
rect 14700 8848 14706 8900
rect 16390 8848 16396 8900
rect 16448 8888 16454 8900
rect 16868 8888 16896 8919
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 17586 8956 17592 8968
rect 17276 8928 17592 8956
rect 17276 8916 17282 8928
rect 17586 8916 17592 8928
rect 17644 8956 17650 8968
rect 17865 8959 17923 8965
rect 17865 8956 17877 8959
rect 17644 8928 17877 8956
rect 17644 8916 17650 8928
rect 17865 8925 17877 8928
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 18966 8956 18972 8968
rect 18012 8928 18972 8956
rect 18012 8916 18018 8928
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 17034 8888 17040 8900
rect 16448 8860 17040 8888
rect 16448 8848 16454 8860
rect 17034 8848 17040 8860
rect 17092 8848 17098 8900
rect 7147 8792 8340 8820
rect 7147 8789 7159 8792
rect 7101 8783 7159 8789
rect 9214 8780 9220 8832
rect 9272 8780 9278 8832
rect 10962 8780 10968 8832
rect 11020 8780 11026 8832
rect 11054 8780 11060 8832
rect 11112 8780 11118 8832
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 14516 8792 16037 8820
rect 14516 8780 14522 8792
rect 16025 8789 16037 8792
rect 16071 8789 16083 8823
rect 16025 8783 16083 8789
rect 16666 8780 16672 8832
rect 16724 8780 16730 8832
rect 1104 8730 18860 8752
rect 1104 8678 5502 8730
rect 5554 8678 5566 8730
rect 5618 8678 5630 8730
rect 5682 8678 5694 8730
rect 5746 8678 5758 8730
rect 5810 8678 5822 8730
rect 5874 8678 5886 8730
rect 5938 8678 5950 8730
rect 6002 8678 6014 8730
rect 6066 8678 6078 8730
rect 6130 8678 6142 8730
rect 6194 8678 6206 8730
rect 6258 8678 6270 8730
rect 6322 8678 6334 8730
rect 6386 8678 6398 8730
rect 6450 8678 6462 8730
rect 6514 8678 6526 8730
rect 6578 8678 6590 8730
rect 6642 8678 6654 8730
rect 6706 8678 13502 8730
rect 13554 8678 13566 8730
rect 13618 8678 13630 8730
rect 13682 8678 13694 8730
rect 13746 8678 13758 8730
rect 13810 8678 13822 8730
rect 13874 8678 13886 8730
rect 13938 8678 13950 8730
rect 14002 8678 14014 8730
rect 14066 8678 14078 8730
rect 14130 8678 14142 8730
rect 14194 8678 14206 8730
rect 14258 8678 14270 8730
rect 14322 8678 14334 8730
rect 14386 8678 14398 8730
rect 14450 8678 14462 8730
rect 14514 8678 14526 8730
rect 14578 8678 14590 8730
rect 14642 8678 14654 8730
rect 14706 8678 18860 8730
rect 1104 8656 18860 8678
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 2740 8588 4169 8616
rect 2740 8576 2746 8588
rect 4157 8585 4169 8588
rect 4203 8585 4215 8619
rect 4157 8579 4215 8585
rect 4430 8576 4436 8628
rect 4488 8616 4494 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 4488 8588 5273 8616
rect 4488 8576 4494 8588
rect 5261 8585 5273 8588
rect 5307 8616 5319 8619
rect 5442 8616 5448 8628
rect 5307 8588 5448 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 7742 8616 7748 8628
rect 6564 8588 7748 8616
rect 2222 8508 2228 8560
rect 2280 8548 2286 8560
rect 2280 8520 3096 8548
rect 2280 8508 2286 8520
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 1903 8452 2329 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2317 8449 2329 8452
rect 2363 8480 2375 8483
rect 2866 8480 2872 8492
rect 2363 8452 2872 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 1688 8412 1716 8443
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3068 8489 3096 8520
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 4304 8520 5488 8548
rect 4304 8508 4310 8520
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3099 8452 4077 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4522 8440 4528 8492
rect 4580 8480 4586 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4580 8452 4905 8480
rect 4580 8440 4586 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 5074 8440 5080 8492
rect 5132 8489 5138 8492
rect 5132 8483 5181 8489
rect 5132 8449 5135 8483
rect 5169 8449 5181 8483
rect 5132 8443 5181 8449
rect 5132 8440 5138 8443
rect 5258 8440 5264 8492
rect 5316 8480 5322 8492
rect 5460 8489 5488 8520
rect 6564 8489 6592 8588
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 12802 8616 12808 8628
rect 11808 8588 12808 8616
rect 7009 8551 7067 8557
rect 7009 8517 7021 8551
rect 7055 8548 7067 8551
rect 8110 8548 8116 8560
rect 7055 8520 8116 8548
rect 7055 8517 7067 8520
rect 7009 8511 7067 8517
rect 8110 8508 8116 8520
rect 8168 8508 8174 8560
rect 8205 8551 8263 8557
rect 8205 8517 8217 8551
rect 8251 8548 8263 8551
rect 9214 8548 9220 8560
rect 8251 8520 9220 8548
rect 8251 8517 8263 8520
rect 8205 8511 8263 8517
rect 9214 8508 9220 8520
rect 9272 8508 9278 8560
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 5316 8452 5365 8480
rect 5316 8440 5322 8452
rect 5353 8449 5365 8452
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 7282 8480 7288 8492
rect 7147 8452 7288 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 2774 8412 2780 8424
rect 1688 8384 2780 8412
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8381 3019 8415
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 2961 8375 3019 8381
rect 3068 8384 3525 8412
rect 2501 8347 2559 8353
rect 2501 8313 2513 8347
rect 2547 8344 2559 8347
rect 2976 8344 3004 8375
rect 3068 8356 3096 8384
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 5276 8412 5304 8440
rect 3513 8375 3571 8381
rect 5092 8384 5304 8412
rect 5092 8356 5120 8384
rect 2547 8316 3004 8344
rect 2547 8313 2559 8316
rect 2501 8307 2559 8313
rect 3050 8304 3056 8356
rect 3108 8304 3114 8356
rect 3602 8304 3608 8356
rect 3660 8344 3666 8356
rect 4709 8347 4767 8353
rect 4709 8344 4721 8347
rect 3660 8316 4721 8344
rect 3660 8304 3666 8316
rect 4709 8313 4721 8316
rect 4755 8313 4767 8347
rect 4709 8307 4767 8313
rect 5074 8304 5080 8356
rect 5132 8304 5138 8356
rect 5258 8304 5264 8356
rect 5316 8344 5322 8356
rect 6564 8344 6592 8443
rect 7282 8440 7288 8452
rect 7340 8480 7346 8492
rect 7653 8483 7711 8489
rect 7340 8452 7604 8480
rect 7340 8440 7346 8452
rect 7576 8412 7604 8452
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 8941 8483 8999 8489
rect 8941 8480 8953 8483
rect 7699 8452 8953 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 8941 8449 8953 8452
rect 8987 8480 8999 8483
rect 9030 8480 9036 8492
rect 8987 8452 9036 8480
rect 8987 8449 8999 8452
rect 8941 8443 8999 8449
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8480 11759 8483
rect 11808 8480 11836 8588
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 13412 8588 13584 8616
rect 13412 8576 13418 8588
rect 12618 8548 12624 8560
rect 12084 8520 12624 8548
rect 12084 8489 12112 8520
rect 12618 8508 12624 8520
rect 12676 8508 12682 8560
rect 13556 8557 13584 8588
rect 15010 8576 15016 8628
rect 15068 8576 15074 8628
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15712 8588 16037 8616
rect 15712 8576 15718 8588
rect 16025 8585 16037 8588
rect 16071 8616 16083 8619
rect 16390 8616 16396 8628
rect 16071 8588 16396 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17865 8619 17923 8625
rect 17865 8616 17877 8619
rect 17368 8588 17877 8616
rect 17368 8576 17374 8588
rect 17865 8585 17877 8588
rect 17911 8616 17923 8619
rect 17954 8616 17960 8628
rect 17911 8588 17960 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 18138 8576 18144 8628
rect 18196 8576 18202 8628
rect 13541 8551 13599 8557
rect 13541 8517 13553 8551
rect 13587 8517 13599 8551
rect 16666 8548 16672 8560
rect 14766 8520 16672 8548
rect 13541 8511 13599 8517
rect 16666 8508 16672 8520
rect 16724 8508 16730 8560
rect 17586 8508 17592 8560
rect 17644 8508 17650 8560
rect 11747 8452 11836 8480
rect 12069 8483 12127 8489
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 9876 8412 9904 8443
rect 7576 8384 9904 8412
rect 9950 8372 9956 8424
rect 10008 8412 10014 8424
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 10008 8384 11805 8412
rect 10008 8372 10014 8384
rect 11793 8381 11805 8384
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 8113 8347 8171 8353
rect 8113 8344 8125 8347
rect 5316 8316 6592 8344
rect 7208 8316 8125 8344
rect 5316 8304 5322 8316
rect 7208 8288 7236 8316
rect 8113 8313 8125 8316
rect 8159 8344 8171 8347
rect 10229 8347 10287 8353
rect 10229 8344 10241 8347
rect 8159 8316 10241 8344
rect 8159 8313 8171 8316
rect 8113 8307 8171 8313
rect 10229 8313 10241 8316
rect 10275 8313 10287 8347
rect 10229 8307 10287 8313
rect 11698 8304 11704 8356
rect 11756 8344 11762 8356
rect 12176 8344 12204 8443
rect 14826 8440 14832 8492
rect 14884 8480 14890 8492
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 14884 8452 15853 8480
rect 14884 8440 14890 8452
rect 15841 8449 15853 8452
rect 15887 8449 15899 8483
rect 15841 8443 15899 8449
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8412 13323 8415
rect 13538 8412 13544 8424
rect 13311 8384 13544 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 13538 8372 13544 8384
rect 13596 8412 13602 8424
rect 15194 8412 15200 8424
rect 13596 8384 15200 8412
rect 13596 8372 13602 8384
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 16132 8412 16160 8443
rect 17402 8440 17408 8492
rect 17460 8480 17466 8492
rect 17773 8483 17831 8489
rect 17773 8480 17785 8483
rect 17460 8452 17785 8480
rect 17460 8440 17466 8452
rect 17773 8449 17785 8452
rect 17819 8449 17831 8483
rect 17773 8443 17831 8449
rect 17957 8483 18015 8489
rect 17957 8449 17969 8483
rect 18003 8480 18015 8483
rect 18046 8480 18052 8492
rect 18003 8452 18052 8480
rect 18003 8449 18015 8452
rect 17957 8443 18015 8449
rect 18046 8440 18052 8452
rect 18104 8480 18110 8492
rect 18782 8480 18788 8492
rect 18104 8452 18788 8480
rect 18104 8440 18110 8452
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 18966 8412 18972 8424
rect 16132 8384 18972 8412
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 11756 8316 12204 8344
rect 11756 8304 11762 8316
rect 15102 8304 15108 8356
rect 15160 8344 15166 8356
rect 15657 8347 15715 8353
rect 15657 8344 15669 8347
rect 15160 8316 15669 8344
rect 15160 8304 15166 8316
rect 15657 8313 15669 8316
rect 15703 8313 15715 8347
rect 15657 8307 15715 8313
rect 16390 8304 16396 8356
rect 16448 8344 16454 8356
rect 17494 8344 17500 8356
rect 16448 8316 17500 8344
rect 16448 8304 16454 8316
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 7190 8236 7196 8288
rect 7248 8236 7254 8288
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12618 8276 12624 8288
rect 12308 8248 12624 8276
rect 12308 8236 12314 8248
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 13354 8276 13360 8288
rect 13228 8248 13360 8276
rect 13228 8236 13234 8248
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 14826 8236 14832 8288
rect 14884 8276 14890 8288
rect 15378 8276 15384 8288
rect 14884 8248 15384 8276
rect 14884 8236 14890 8248
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 17126 8276 17132 8288
rect 16724 8248 17132 8276
rect 16724 8236 16730 8248
rect 17126 8236 17132 8248
rect 17184 8236 17190 8288
rect 17678 8236 17684 8288
rect 17736 8276 17742 8288
rect 17736 8248 18920 8276
rect 17736 8236 17742 8248
rect 1104 8186 18860 8208
rect 1104 8134 1502 8186
rect 1554 8134 1566 8186
rect 1618 8134 1630 8186
rect 1682 8134 1694 8186
rect 1746 8134 1758 8186
rect 1810 8134 1822 8186
rect 1874 8134 1886 8186
rect 1938 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 2270 8186
rect 2322 8134 2334 8186
rect 2386 8134 2398 8186
rect 2450 8134 2462 8186
rect 2514 8134 2526 8186
rect 2578 8134 2590 8186
rect 2642 8134 2654 8186
rect 2706 8134 9502 8186
rect 9554 8134 9566 8186
rect 9618 8134 9630 8186
rect 9682 8134 9694 8186
rect 9746 8134 9758 8186
rect 9810 8134 9822 8186
rect 9874 8134 9886 8186
rect 9938 8134 9950 8186
rect 10002 8134 10014 8186
rect 10066 8134 10078 8186
rect 10130 8134 10142 8186
rect 10194 8134 10206 8186
rect 10258 8134 10270 8186
rect 10322 8134 10334 8186
rect 10386 8134 10398 8186
rect 10450 8134 10462 8186
rect 10514 8134 10526 8186
rect 10578 8134 10590 8186
rect 10642 8134 10654 8186
rect 10706 8134 17502 8186
rect 17554 8134 17566 8186
rect 17618 8134 17630 8186
rect 17682 8134 17694 8186
rect 17746 8134 17758 8186
rect 17810 8134 17822 8186
rect 17874 8134 17886 8186
rect 17938 8134 17950 8186
rect 18002 8134 18014 8186
rect 18066 8134 18078 8186
rect 18130 8134 18142 8186
rect 18194 8134 18206 8186
rect 18258 8134 18270 8186
rect 18322 8134 18334 8186
rect 18386 8134 18398 8186
rect 18450 8134 18462 8186
rect 18514 8134 18526 8186
rect 18578 8134 18590 8186
rect 18642 8134 18654 8186
rect 18706 8134 18860 8186
rect 1104 8112 18860 8134
rect 382 8032 388 8084
rect 440 8072 446 8084
rect 934 8072 940 8084
rect 440 8044 940 8072
rect 440 8032 446 8044
rect 934 8032 940 8044
rect 992 8032 998 8084
rect 1302 8032 1308 8084
rect 1360 8072 1366 8084
rect 2130 8072 2136 8084
rect 1360 8044 2136 8072
rect 1360 8032 1366 8044
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 11606 8072 11612 8084
rect 10091 8044 11612 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 12526 8072 12532 8084
rect 12360 8044 12532 8072
rect 3694 7964 3700 8016
rect 3752 8004 3758 8016
rect 10689 8007 10747 8013
rect 3752 7976 5580 8004
rect 3752 7964 3758 7976
rect 2866 7936 2872 7948
rect 1596 7908 2872 7936
rect 1596 7877 1624 7908
rect 2866 7896 2872 7908
rect 2924 7936 2930 7948
rect 2924 7908 4108 7936
rect 2924 7896 2930 7908
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7837 1639 7871
rect 1581 7831 1639 7837
rect 2130 7828 2136 7880
rect 2188 7828 2194 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3694 7868 3700 7880
rect 3283 7840 3700 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 3694 7828 3700 7840
rect 3752 7828 3758 7880
rect 4080 7877 4108 7908
rect 5552 7877 5580 7976
rect 10689 7973 10701 8007
rect 10735 8004 10747 8007
rect 10735 7976 10916 8004
rect 10735 7973 10747 7976
rect 10689 7967 10747 7973
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 6880 7908 7757 7936
rect 6880 7896 6886 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 7745 7899 7803 7905
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 10888 7936 10916 7976
rect 11422 7936 11428 7948
rect 7892 7908 10824 7936
rect 10888 7908 11428 7936
rect 7892 7896 7898 7908
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 7190 7868 7196 7880
rect 6595 7840 7196 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 8220 7840 9321 7868
rect 1673 7803 1731 7809
rect 1673 7769 1685 7803
rect 1719 7769 1731 7803
rect 1673 7763 1731 7769
rect 1688 7732 1716 7763
rect 2682 7760 2688 7812
rect 2740 7760 2746 7812
rect 2774 7760 2780 7812
rect 2832 7800 2838 7812
rect 3973 7803 4031 7809
rect 3973 7800 3985 7803
rect 2832 7772 3985 7800
rect 2832 7760 2838 7772
rect 3973 7769 3985 7772
rect 4019 7769 4031 7803
rect 3973 7763 4031 7769
rect 6365 7803 6423 7809
rect 6365 7769 6377 7803
rect 6411 7800 6423 7803
rect 7300 7800 7328 7828
rect 6411 7772 7328 7800
rect 6411 7769 6423 7772
rect 6365 7763 6423 7769
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 8220 7809 8248 7840
rect 9309 7837 9321 7840
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9766 7828 9772 7880
rect 9824 7828 9830 7880
rect 8205 7803 8263 7809
rect 8205 7800 8217 7803
rect 8168 7772 8217 7800
rect 8168 7760 8174 7772
rect 8205 7769 8217 7772
rect 8251 7769 8263 7803
rect 8205 7763 8263 7769
rect 8297 7803 8355 7809
rect 8297 7769 8309 7803
rect 8343 7769 8355 7803
rect 8297 7763 8355 7769
rect 3050 7732 3056 7744
rect 1688 7704 3056 7732
rect 3050 7692 3056 7704
rect 3108 7692 3114 7744
rect 7101 7735 7159 7741
rect 7101 7701 7113 7735
rect 7147 7732 7159 7735
rect 8312 7732 8340 7763
rect 9398 7760 9404 7812
rect 9456 7800 9462 7812
rect 9950 7800 9956 7812
rect 9456 7772 9956 7800
rect 9456 7760 9462 7772
rect 9950 7760 9956 7772
rect 10008 7760 10014 7812
rect 7147 7704 8340 7732
rect 7147 7701 7159 7704
rect 7101 7695 7159 7701
rect 9214 7692 9220 7744
rect 9272 7692 9278 7744
rect 10796 7732 10824 7908
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 12161 7939 12219 7945
rect 12161 7905 12173 7939
rect 12207 7936 12219 7939
rect 12360 7936 12388 8044
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12710 8032 12716 8084
rect 12768 8072 12774 8084
rect 13357 8075 13415 8081
rect 13357 8072 13369 8075
rect 12768 8044 13369 8072
rect 12768 8032 12774 8044
rect 13357 8041 13369 8044
rect 13403 8041 13415 8075
rect 17126 8072 17132 8084
rect 13357 8035 13415 8041
rect 14752 8044 17132 8072
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 14752 8013 14780 8044
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 17310 8032 17316 8084
rect 17368 8032 17374 8084
rect 12989 8007 13047 8013
rect 12989 8004 13001 8007
rect 12676 7976 13001 8004
rect 12676 7964 12682 7976
rect 12989 7973 13001 7976
rect 13035 7973 13047 8007
rect 12989 7967 13047 7973
rect 14737 8007 14795 8013
rect 14737 7973 14749 8007
rect 14783 7973 14795 8007
rect 14737 7967 14795 7973
rect 12207 7908 12388 7936
rect 12437 7939 12495 7945
rect 12207 7905 12219 7908
rect 12161 7899 12219 7905
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 12526 7936 12532 7948
rect 12483 7908 12532 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 12526 7896 12532 7908
rect 12584 7936 12590 7948
rect 13538 7936 13544 7948
rect 12584 7908 13544 7936
rect 12584 7896 12590 7908
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 15838 7896 15844 7948
rect 15896 7896 15902 7948
rect 17034 7896 17040 7948
rect 17092 7936 17098 7948
rect 17092 7908 17908 7936
rect 17092 7896 17098 7908
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12860 7840 12909 7868
rect 12860 7828 12866 7840
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 13078 7828 13084 7880
rect 13136 7868 13142 7880
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 13136 7840 13185 7868
rect 13136 7828 13142 7840
rect 13173 7837 13185 7840
rect 13219 7868 13231 7871
rect 13219 7840 14504 7868
rect 13219 7837 13231 7840
rect 13173 7831 13231 7837
rect 12066 7800 12072 7812
rect 11730 7772 12072 7800
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 14369 7803 14427 7809
rect 14369 7800 14381 7803
rect 12406 7772 14381 7800
rect 12406 7732 12434 7772
rect 14369 7769 14381 7772
rect 14415 7769 14427 7803
rect 14476 7800 14504 7840
rect 14550 7828 14556 7880
rect 14608 7828 14614 7880
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 14844 7800 14872 7831
rect 15286 7828 15292 7880
rect 15344 7868 15350 7880
rect 17880 7877 17908 7908
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 15344 7840 15577 7868
rect 15344 7828 15350 7840
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18892 7868 18920 8248
rect 18187 7840 18920 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 14476 7772 14872 7800
rect 14369 7763 14427 7769
rect 16850 7760 16856 7812
rect 16908 7760 16914 7812
rect 10796 7704 12434 7732
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 14090 7732 14096 7744
rect 12768 7704 14096 7732
rect 12768 7692 12774 7704
rect 14090 7692 14096 7704
rect 14148 7692 14154 7744
rect 17954 7692 17960 7744
rect 18012 7692 18018 7744
rect 1104 7642 18860 7664
rect 1104 7590 5502 7642
rect 5554 7590 5566 7642
rect 5618 7590 5630 7642
rect 5682 7590 5694 7642
rect 5746 7590 5758 7642
rect 5810 7590 5822 7642
rect 5874 7590 5886 7642
rect 5938 7590 5950 7642
rect 6002 7590 6014 7642
rect 6066 7590 6078 7642
rect 6130 7590 6142 7642
rect 6194 7590 6206 7642
rect 6258 7590 6270 7642
rect 6322 7590 6334 7642
rect 6386 7590 6398 7642
rect 6450 7590 6462 7642
rect 6514 7590 6526 7642
rect 6578 7590 6590 7642
rect 6642 7590 6654 7642
rect 6706 7590 13502 7642
rect 13554 7590 13566 7642
rect 13618 7590 13630 7642
rect 13682 7590 13694 7642
rect 13746 7590 13758 7642
rect 13810 7590 13822 7642
rect 13874 7590 13886 7642
rect 13938 7590 13950 7642
rect 14002 7590 14014 7642
rect 14066 7590 14078 7642
rect 14130 7590 14142 7642
rect 14194 7590 14206 7642
rect 14258 7590 14270 7642
rect 14322 7590 14334 7642
rect 14386 7590 14398 7642
rect 14450 7590 14462 7642
rect 14514 7590 14526 7642
rect 14578 7590 14590 7642
rect 14642 7590 14654 7642
rect 14706 7590 18860 7642
rect 19334 7624 19340 7676
rect 19392 7624 19398 7676
rect 1104 7568 18860 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 4157 7531 4215 7537
rect 4157 7528 4169 7531
rect 2740 7500 4169 7528
rect 2740 7488 2746 7500
rect 4157 7497 4169 7500
rect 4203 7497 4215 7531
rect 4157 7491 4215 7497
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5626 7528 5632 7540
rect 4948 7500 5632 7528
rect 4948 7488 4954 7500
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 6914 7528 6920 7540
rect 5951 7500 6920 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7340 7500 9352 7528
rect 7340 7488 7346 7500
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 2958 7460 2964 7472
rect 1719 7432 2964 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 3050 7420 3056 7472
rect 3108 7460 3114 7472
rect 4065 7463 4123 7469
rect 4065 7460 4077 7463
rect 3108 7432 4077 7460
rect 3108 7420 3114 7432
rect 4065 7429 4077 7432
rect 4111 7429 4123 7463
rect 4065 7423 4123 7429
rect 7009 7463 7067 7469
rect 7009 7429 7021 7463
rect 7055 7460 7067 7463
rect 8110 7460 8116 7472
rect 7055 7432 8116 7460
rect 7055 7429 7067 7432
rect 7009 7423 7067 7429
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 8205 7463 8263 7469
rect 8205 7429 8217 7463
rect 8251 7460 8263 7463
rect 9214 7460 9220 7472
rect 8251 7432 9220 7460
rect 8251 7429 8263 7432
rect 8205 7423 8263 7429
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2317 7395 2375 7401
rect 2317 7392 2329 7395
rect 1903 7364 2329 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2317 7361 2329 7364
rect 2363 7392 2375 7395
rect 2866 7392 2872 7404
rect 2363 7364 2872 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7392 5319 7395
rect 6549 7395 6607 7401
rect 5307 7364 6500 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2746 7296 2973 7324
rect 2501 7259 2559 7265
rect 2501 7225 2513 7259
rect 2547 7256 2559 7259
rect 2746 7256 2774 7296
rect 2961 7293 2973 7296
rect 3007 7293 3019 7327
rect 2961 7287 3019 7293
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7293 3571 7327
rect 3513 7287 3571 7293
rect 2547 7228 2774 7256
rect 2547 7225 2559 7228
rect 2501 7219 2559 7225
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 3528 7188 3556 7287
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 5445 7327 5503 7333
rect 5445 7324 5457 7327
rect 3752 7296 5457 7324
rect 3752 7284 3758 7296
rect 5445 7293 5457 7296
rect 5491 7293 5503 7327
rect 5445 7287 5503 7293
rect 5534 7284 5540 7336
rect 5592 7284 5598 7336
rect 5626 7284 5632 7336
rect 5684 7284 5690 7336
rect 5718 7284 5724 7336
rect 5776 7284 5782 7336
rect 2188 7160 3556 7188
rect 6472 7188 6500 7364
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 6822 7392 6828 7404
rect 6595 7364 6828 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7392 7159 7395
rect 7282 7392 7288 7404
rect 7147 7364 7288 7392
rect 7147 7361 7159 7364
rect 7101 7355 7159 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7392 7711 7395
rect 7742 7392 7748 7404
rect 7699 7364 7748 7392
rect 7699 7361 7711 7364
rect 7653 7355 7711 7361
rect 7742 7352 7748 7364
rect 7800 7392 7806 7404
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 7800 7364 8953 7392
rect 7800 7352 7806 7364
rect 8941 7361 8953 7364
rect 8987 7361 8999 7395
rect 9324 7392 9352 7500
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 13078 7528 13084 7540
rect 11296 7500 13084 7528
rect 11296 7488 11302 7500
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 17954 7528 17960 7540
rect 15120 7500 17960 7528
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 11054 7460 11060 7472
rect 9824 7432 11060 7460
rect 9824 7420 9830 7432
rect 11054 7420 11060 7432
rect 11112 7460 11118 7472
rect 12250 7460 12256 7472
rect 11112 7432 12256 7460
rect 11112 7420 11118 7432
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 15120 7460 15148 7500
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 16482 7460 16488 7472
rect 13294 7432 15148 7460
rect 15962 7432 16488 7460
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 17218 7420 17224 7472
rect 17276 7460 17282 7472
rect 17681 7463 17739 7469
rect 17681 7460 17693 7463
rect 17276 7432 17693 7460
rect 17276 7420 17282 7432
rect 17681 7429 17693 7432
rect 17727 7429 17739 7463
rect 17681 7423 17739 7429
rect 19058 7420 19064 7472
rect 19116 7460 19122 7472
rect 19352 7460 19380 7624
rect 19116 7432 19380 7460
rect 19116 7420 19122 7432
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 9324 7364 9873 7392
rect 8941 7355 8999 7361
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9950 7352 9956 7404
rect 10008 7392 10014 7404
rect 11606 7392 11612 7404
rect 10008 7364 11612 7392
rect 10008 7352 10014 7364
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11112 7296 12756 7324
rect 11112 7284 11118 7296
rect 6914 7216 6920 7268
rect 6972 7256 6978 7268
rect 8113 7259 8171 7265
rect 8113 7256 8125 7259
rect 6972 7228 8125 7256
rect 6972 7216 6978 7228
rect 8113 7225 8125 7228
rect 8159 7256 8171 7259
rect 10229 7259 10287 7265
rect 10229 7256 10241 7259
rect 8159 7228 10241 7256
rect 8159 7225 8171 7228
rect 8113 7219 8171 7225
rect 10229 7225 10241 7228
rect 10275 7225 10287 7259
rect 10229 7219 10287 7225
rect 12253 7259 12311 7265
rect 12253 7225 12265 7259
rect 12299 7256 12311 7259
rect 12618 7256 12624 7268
rect 12299 7228 12624 7256
rect 12299 7225 12311 7228
rect 12253 7219 12311 7225
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 11238 7188 11244 7200
rect 6472 7160 11244 7188
rect 2188 7148 2194 7160
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 12728 7188 12756 7296
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 13725 7327 13783 7333
rect 13725 7324 13737 7327
rect 13320 7296 13737 7324
rect 13320 7284 13326 7296
rect 13725 7293 13737 7296
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 13998 7284 14004 7336
rect 14056 7324 14062 7336
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 14056 7296 14473 7324
rect 14056 7284 14062 7296
rect 14461 7293 14473 7296
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 14737 7327 14795 7333
rect 14737 7293 14749 7327
rect 14783 7324 14795 7327
rect 17773 7327 17831 7333
rect 14783 7296 17356 7324
rect 14783 7293 14795 7296
rect 14737 7287 14795 7293
rect 17328 7265 17356 7296
rect 17773 7293 17785 7327
rect 17819 7293 17831 7327
rect 17773 7287 17831 7293
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7324 18015 7327
rect 18003 7296 18920 7324
rect 18003 7293 18015 7296
rect 17957 7287 18015 7293
rect 17313 7259 17371 7265
rect 17313 7225 17325 7259
rect 17359 7225 17371 7259
rect 17313 7219 17371 7225
rect 14734 7188 14740 7200
rect 12728 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 16209 7191 16267 7197
rect 16209 7157 16221 7191
rect 16255 7188 16267 7191
rect 17402 7188 17408 7200
rect 16255 7160 17408 7188
rect 16255 7157 16267 7160
rect 16209 7151 16267 7157
rect 17402 7148 17408 7160
rect 17460 7188 17466 7200
rect 17788 7188 17816 7287
rect 17460 7160 17816 7188
rect 17460 7148 17466 7160
rect 1104 7098 18860 7120
rect 1104 7046 1502 7098
rect 1554 7046 1566 7098
rect 1618 7046 1630 7098
rect 1682 7046 1694 7098
rect 1746 7046 1758 7098
rect 1810 7046 1822 7098
rect 1874 7046 1886 7098
rect 1938 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 2270 7098
rect 2322 7046 2334 7098
rect 2386 7046 2398 7098
rect 2450 7046 2462 7098
rect 2514 7046 2526 7098
rect 2578 7046 2590 7098
rect 2642 7046 2654 7098
rect 2706 7046 9502 7098
rect 9554 7046 9566 7098
rect 9618 7046 9630 7098
rect 9682 7046 9694 7098
rect 9746 7046 9758 7098
rect 9810 7046 9822 7098
rect 9874 7046 9886 7098
rect 9938 7046 9950 7098
rect 10002 7046 10014 7098
rect 10066 7046 10078 7098
rect 10130 7046 10142 7098
rect 10194 7046 10206 7098
rect 10258 7046 10270 7098
rect 10322 7046 10334 7098
rect 10386 7046 10398 7098
rect 10450 7046 10462 7098
rect 10514 7046 10526 7098
rect 10578 7046 10590 7098
rect 10642 7046 10654 7098
rect 10706 7046 17502 7098
rect 17554 7046 17566 7098
rect 17618 7046 17630 7098
rect 17682 7046 17694 7098
rect 17746 7046 17758 7098
rect 17810 7046 17822 7098
rect 17874 7046 17886 7098
rect 17938 7046 17950 7098
rect 18002 7046 18014 7098
rect 18066 7046 18078 7098
rect 18130 7046 18142 7098
rect 18194 7046 18206 7098
rect 18258 7046 18270 7098
rect 18322 7046 18334 7098
rect 18386 7046 18398 7098
rect 18450 7046 18462 7098
rect 18514 7046 18526 7098
rect 18578 7046 18590 7098
rect 18642 7046 18654 7098
rect 18706 7046 18860 7098
rect 1104 7024 18860 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 3326 6984 3332 6996
rect 1452 6956 3332 6984
rect 1452 6944 1458 6956
rect 3326 6944 3332 6956
rect 3384 6944 3390 6996
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 9861 6987 9919 6993
rect 9861 6984 9873 6987
rect 8536 6956 9873 6984
rect 8536 6944 8542 6956
rect 9861 6953 9873 6956
rect 9907 6953 9919 6987
rect 9861 6947 9919 6953
rect 11146 6944 11152 6996
rect 11204 6984 11210 6996
rect 11345 6987 11403 6993
rect 11345 6984 11357 6987
rect 11204 6956 11357 6984
rect 11204 6944 11210 6956
rect 11345 6953 11357 6956
rect 11391 6953 11403 6987
rect 11345 6947 11403 6953
rect 11606 6944 11612 6996
rect 11664 6984 11670 6996
rect 17402 6984 17408 6996
rect 11664 6956 17408 6984
rect 11664 6944 11670 6956
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 12526 6916 12532 6928
rect 12084 6888 12532 6916
rect 2774 6848 2780 6860
rect 1596 6820 2780 6848
rect 1596 6789 1624 6820
rect 2774 6808 2780 6820
rect 2832 6848 2838 6860
rect 2832 6820 4108 6848
rect 2832 6808 2838 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6749 1639 6783
rect 1581 6743 1639 6749
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6780 2191 6783
rect 3142 6780 3148 6792
rect 2179 6752 3148 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3234 6740 3240 6792
rect 3292 6740 3298 6792
rect 4080 6789 4108 6820
rect 12084 6792 12112 6888
rect 12526 6876 12532 6888
rect 12584 6916 12590 6928
rect 13262 6916 13268 6928
rect 12584 6888 13268 6916
rect 12584 6876 12590 6888
rect 13262 6876 13268 6888
rect 13320 6916 13326 6928
rect 13998 6916 14004 6928
rect 13320 6888 14004 6916
rect 13320 6876 13326 6888
rect 13998 6876 14004 6888
rect 14056 6876 14062 6928
rect 15838 6876 15844 6928
rect 15896 6916 15902 6928
rect 16298 6916 16304 6928
rect 15896 6888 16304 6916
rect 15896 6876 15902 6888
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6848 12771 6851
rect 13078 6848 13084 6860
rect 12759 6820 13084 6848
rect 12759 6817 12771 6820
rect 12713 6811 12771 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 14016 6848 14044 6876
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 13280 6820 13584 6848
rect 14016 6820 14289 6848
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 6914 6780 6920 6792
rect 6595 6752 6920 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 2222 6712 2228 6724
rect 1719 6684 2228 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 2682 6672 2688 6724
rect 2740 6672 2746 6724
rect 2777 6715 2835 6721
rect 2777 6681 2789 6715
rect 2823 6712 2835 6715
rect 2958 6712 2964 6724
rect 2823 6684 2964 6712
rect 2823 6681 2835 6684
rect 2777 6675 2835 6681
rect 2958 6672 2964 6684
rect 3016 6712 3022 6724
rect 3973 6715 4031 6721
rect 3973 6712 3985 6715
rect 3016 6684 3985 6712
rect 3016 6672 3022 6684
rect 3973 6681 3985 6684
rect 4019 6681 4031 6715
rect 3973 6675 4031 6681
rect 3234 6604 3240 6656
rect 3292 6644 3298 6656
rect 5552 6644 5580 6743
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7282 6740 7288 6792
rect 7340 6740 7346 6792
rect 7742 6740 7748 6792
rect 7800 6740 7806 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 8220 6752 9321 6780
rect 6365 6715 6423 6721
rect 6365 6681 6377 6715
rect 6411 6712 6423 6715
rect 7300 6712 7328 6740
rect 6411 6684 7328 6712
rect 6411 6681 6423 6684
rect 6365 6675 6423 6681
rect 7466 6672 7472 6724
rect 7524 6712 7530 6724
rect 7926 6712 7932 6724
rect 7524 6684 7932 6712
rect 7524 6672 7530 6684
rect 7926 6672 7932 6684
rect 7984 6672 7990 6724
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 8220 6721 8248 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6780 11667 6783
rect 12066 6780 12072 6792
rect 11655 6752 12072 6780
rect 11655 6749 11667 6752
rect 11609 6743 11667 6749
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 13280 6780 13308 6820
rect 12584 6752 13308 6780
rect 12584 6740 12590 6752
rect 13354 6740 13360 6792
rect 13412 6740 13418 6792
rect 13556 6789 13584 6820
rect 14277 6817 14289 6820
rect 14323 6848 14335 6851
rect 15286 6848 15292 6860
rect 14323 6820 15292 6848
rect 14323 6817 14335 6820
rect 14277 6811 14335 6817
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 18325 6851 18383 6857
rect 18325 6848 18337 6851
rect 16264 6820 18337 6848
rect 16264 6808 16270 6820
rect 18325 6817 18337 6820
rect 18371 6848 18383 6851
rect 18892 6848 18920 7296
rect 18371 6820 18920 6848
rect 18371 6817 18383 6820
rect 18325 6811 18383 6817
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 13541 6743 13599 6749
rect 16040 6752 17509 6780
rect 8205 6715 8263 6721
rect 8205 6712 8217 6715
rect 8168 6684 8217 6712
rect 8168 6672 8174 6684
rect 8205 6681 8217 6684
rect 8251 6681 8263 6715
rect 8205 6675 8263 6681
rect 8297 6715 8355 6721
rect 8297 6681 8309 6715
rect 8343 6681 8355 6715
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 10902 6684 11284 6712
rect 8297 6675 8355 6681
rect 3292 6616 5580 6644
rect 7101 6647 7159 6653
rect 3292 6604 3298 6616
rect 7101 6613 7113 6647
rect 7147 6644 7159 6647
rect 8312 6644 8340 6675
rect 7147 6616 8340 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 9214 6604 9220 6656
rect 9272 6604 9278 6656
rect 11256 6644 11284 6684
rect 11440 6684 13277 6712
rect 11440 6644 11468 6684
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 13265 6675 13323 6681
rect 14553 6715 14611 6721
rect 14553 6681 14565 6715
rect 14599 6712 14611 6715
rect 14826 6712 14832 6724
rect 14599 6684 14832 6712
rect 14599 6681 14611 6684
rect 14553 6675 14611 6681
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 15562 6672 15568 6724
rect 15620 6672 15626 6724
rect 16040 6656 16068 6752
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 17770 6740 17776 6792
rect 17828 6740 17834 6792
rect 11256 6616 11468 6644
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 11848 6616 12081 6644
rect 11848 6604 11854 6616
rect 12069 6613 12081 6616
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 12308 6616 12541 6644
rect 12308 6604 12314 6616
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 12529 6607 12587 6613
rect 16022 6604 16028 6656
rect 16080 6604 16086 6656
rect 1104 6554 18860 6576
rect 1104 6502 5502 6554
rect 5554 6502 5566 6554
rect 5618 6502 5630 6554
rect 5682 6502 5694 6554
rect 5746 6502 5758 6554
rect 5810 6502 5822 6554
rect 5874 6502 5886 6554
rect 5938 6502 5950 6554
rect 6002 6502 6014 6554
rect 6066 6502 6078 6554
rect 6130 6502 6142 6554
rect 6194 6502 6206 6554
rect 6258 6502 6270 6554
rect 6322 6502 6334 6554
rect 6386 6502 6398 6554
rect 6450 6502 6462 6554
rect 6514 6502 6526 6554
rect 6578 6502 6590 6554
rect 6642 6502 6654 6554
rect 6706 6502 13502 6554
rect 13554 6502 13566 6554
rect 13618 6502 13630 6554
rect 13682 6502 13694 6554
rect 13746 6502 13758 6554
rect 13810 6502 13822 6554
rect 13874 6502 13886 6554
rect 13938 6502 13950 6554
rect 14002 6502 14014 6554
rect 14066 6502 14078 6554
rect 14130 6502 14142 6554
rect 14194 6502 14206 6554
rect 14258 6502 14270 6554
rect 14322 6502 14334 6554
rect 14386 6502 14398 6554
rect 14450 6502 14462 6554
rect 14514 6502 14526 6554
rect 14578 6502 14590 6554
rect 14642 6502 14654 6554
rect 14706 6502 18860 6554
rect 1104 6480 18860 6502
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 4157 6443 4215 6449
rect 4157 6440 4169 6443
rect 2740 6412 4169 6440
rect 2740 6400 2746 6412
rect 4157 6409 4169 6412
rect 4203 6409 4215 6443
rect 4157 6403 4215 6409
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 7742 6440 7748 6452
rect 5132 6412 5764 6440
rect 5132 6400 5138 6412
rect 2222 6332 2228 6384
rect 2280 6372 2286 6384
rect 2280 6344 3096 6372
rect 2280 6332 2286 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 1903 6276 2329 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 2317 6273 2329 6276
rect 2363 6304 2375 6307
rect 2774 6304 2780 6316
rect 2363 6276 2780 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 1688 6236 1716 6267
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 3068 6313 3096 6344
rect 5258 6332 5264 6384
rect 5316 6332 5322 6384
rect 5736 6372 5764 6412
rect 6564 6412 7748 6440
rect 5905 6375 5963 6381
rect 5905 6372 5917 6375
rect 5736 6344 5917 6372
rect 5905 6341 5917 6344
rect 5951 6341 5963 6375
rect 5905 6335 5963 6341
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 3099 6276 4077 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 4890 6304 4896 6316
rect 4580 6276 4896 6304
rect 4580 6264 4586 6276
rect 4890 6264 4896 6276
rect 4948 6304 4954 6316
rect 6564 6313 6592 6412
rect 7742 6400 7748 6412
rect 7800 6440 7806 6452
rect 12986 6440 12992 6452
rect 7800 6412 12992 6440
rect 7800 6400 7806 6412
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 15010 6440 15016 6452
rect 13740 6412 15016 6440
rect 7009 6375 7067 6381
rect 7009 6341 7021 6375
rect 7055 6372 7067 6375
rect 8110 6372 8116 6384
rect 7055 6344 8116 6372
rect 7055 6341 7067 6344
rect 7009 6335 7067 6341
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 8205 6375 8263 6381
rect 8205 6341 8217 6375
rect 8251 6372 8263 6375
rect 9214 6372 9220 6384
rect 8251 6344 9220 6372
rect 8251 6341 8263 6344
rect 8205 6335 8263 6341
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 11422 6372 11428 6384
rect 11112 6344 11428 6372
rect 11112 6332 11118 6344
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 13740 6372 13768 6412
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 17218 6440 17224 6452
rect 15436 6412 17224 6440
rect 15436 6400 15442 6412
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 13386 6344 13768 6372
rect 13817 6375 13875 6381
rect 13817 6341 13829 6375
rect 13863 6372 13875 6375
rect 13863 6344 14136 6372
rect 13863 6341 13875 6344
rect 13817 6335 13875 6341
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 4948 6276 5457 6304
rect 4948 6264 4954 6276
rect 5445 6273 5457 6276
rect 5491 6273 5503 6307
rect 5782 6307 5840 6313
rect 5782 6304 5794 6307
rect 5445 6267 5503 6273
rect 5644 6276 5794 6304
rect 2866 6236 2872 6248
rect 1688 6208 2872 6236
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6205 3019 6239
rect 2961 6199 3019 6205
rect 2501 6171 2559 6177
rect 2501 6137 2513 6171
rect 2547 6168 2559 6171
rect 2976 6168 3004 6199
rect 3142 6196 3148 6248
rect 3200 6236 3206 6248
rect 3513 6239 3571 6245
rect 3513 6236 3525 6239
rect 3200 6208 3525 6236
rect 3200 6196 3206 6208
rect 3513 6205 3525 6208
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 4430 6196 4436 6248
rect 4488 6236 4494 6248
rect 5258 6236 5264 6248
rect 4488 6208 5264 6236
rect 4488 6196 4494 6208
rect 5258 6196 5264 6208
rect 5316 6236 5322 6248
rect 5644 6236 5672 6276
rect 5782 6273 5794 6276
rect 5828 6273 5840 6307
rect 5782 6267 5840 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6304 7159 6307
rect 7282 6304 7288 6316
rect 7147 6276 7288 6304
rect 7147 6273 7159 6276
rect 7101 6267 7159 6273
rect 7282 6264 7288 6276
rect 7340 6304 7346 6316
rect 7340 6276 7788 6304
rect 7340 6264 7346 6276
rect 5316 6208 5672 6236
rect 5704 6239 5762 6245
rect 5316 6196 5322 6208
rect 5704 6205 5716 6239
rect 5750 6236 5762 6239
rect 5997 6239 6055 6245
rect 5750 6208 5856 6236
rect 5750 6205 5762 6208
rect 5704 6199 5762 6205
rect 2547 6140 3004 6168
rect 2547 6137 2559 6140
rect 2501 6131 2559 6137
rect 5828 6100 5856 6208
rect 5997 6205 6009 6239
rect 6043 6236 6055 6239
rect 6822 6236 6828 6248
rect 6043 6208 6828 6236
rect 6043 6205 6055 6208
rect 5997 6199 6055 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7653 6239 7711 6245
rect 7653 6236 7665 6239
rect 7524 6208 7665 6236
rect 7524 6196 7530 6208
rect 7653 6205 7665 6208
rect 7699 6205 7711 6239
rect 7760 6236 7788 6276
rect 7926 6264 7932 6316
rect 7984 6304 7990 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 7984 6276 8953 6304
rect 7984 6264 7990 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6273 9919 6307
rect 9861 6267 9919 6273
rect 9876 6236 9904 6267
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 12526 6304 12532 6316
rect 11204 6276 12532 6304
rect 11204 6264 11210 6276
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 14108 6304 14136 6344
rect 14550 6332 14556 6384
rect 14608 6372 14614 6384
rect 14608 6344 14872 6372
rect 14608 6332 14614 6344
rect 14366 6304 14372 6316
rect 14108 6276 14372 6304
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 14844 6313 14872 6344
rect 15102 6332 15108 6384
rect 15160 6372 15166 6384
rect 16206 6372 16212 6384
rect 15160 6344 16212 6372
rect 15160 6332 15166 6344
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 14476 6276 14657 6304
rect 7760 6208 9904 6236
rect 11057 6239 11115 6245
rect 7653 6199 7711 6205
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 11238 6236 11244 6248
rect 11103 6208 11244 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 12250 6236 12256 6248
rect 11480 6208 12256 6236
rect 11480 6196 11486 6208
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 12345 6239 12403 6245
rect 12345 6205 12357 6239
rect 12391 6236 12403 6239
rect 12434 6236 12440 6248
rect 12391 6208 12440 6236
rect 12391 6205 12403 6208
rect 12345 6199 12403 6205
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13320 6208 14105 6236
rect 13320 6196 13326 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 6546 6128 6552 6180
rect 6604 6168 6610 6180
rect 8113 6171 8171 6177
rect 8113 6168 8125 6171
rect 6604 6140 8125 6168
rect 6604 6128 6610 6140
rect 8113 6137 8125 6140
rect 8159 6168 8171 6171
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 8159 6140 10241 6168
rect 8159 6137 8171 6140
rect 8113 6131 8171 6137
rect 10229 6137 10241 6140
rect 10275 6137 10287 6171
rect 10229 6131 10287 6137
rect 6822 6100 6828 6112
rect 5828 6072 6828 6100
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 12618 6100 12624 6112
rect 7156 6072 12624 6100
rect 7156 6060 7162 6072
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 14476 6100 14504 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 14829 6307 14887 6313
rect 14829 6273 14841 6307
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 15378 6264 15384 6316
rect 15436 6264 15442 6316
rect 15654 6310 15660 6316
rect 15580 6282 15660 6310
rect 15580 6245 15608 6282
rect 15654 6264 15660 6282
rect 15712 6264 15718 6316
rect 15764 6313 15792 6344
rect 16206 6332 16212 6344
rect 16264 6332 16270 6384
rect 18325 6375 18383 6381
rect 18325 6341 18337 6375
rect 18371 6372 18383 6375
rect 18782 6372 18788 6384
rect 18371 6344 18788 6372
rect 18371 6341 18383 6344
rect 18325 6335 18383 6341
rect 18782 6332 18788 6344
rect 18840 6332 18846 6384
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6273 15807 6307
rect 15749 6267 15807 6273
rect 15930 6264 15936 6316
rect 15988 6264 15994 6316
rect 16022 6264 16028 6316
rect 16080 6304 16086 6316
rect 17313 6307 17371 6313
rect 17313 6304 17325 6307
rect 16080 6276 17325 6304
rect 16080 6264 16086 6276
rect 17313 6273 17325 6276
rect 17359 6273 17371 6307
rect 17313 6267 17371 6273
rect 17770 6264 17776 6316
rect 17828 6264 17834 6316
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6205 15623 6239
rect 15565 6199 15623 6205
rect 14642 6128 14648 6180
rect 14700 6128 14706 6180
rect 17034 6128 17040 6180
rect 17092 6168 17098 6180
rect 17788 6168 17816 6264
rect 17092 6140 17816 6168
rect 17092 6128 17098 6140
rect 13412 6072 14504 6100
rect 13412 6060 13418 6072
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 16942 6100 16948 6112
rect 15068 6072 16948 6100
rect 15068 6060 15074 6072
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 1104 6010 18860 6032
rect 1104 5958 1502 6010
rect 1554 5958 1566 6010
rect 1618 5958 1630 6010
rect 1682 5958 1694 6010
rect 1746 5958 1758 6010
rect 1810 5958 1822 6010
rect 1874 5958 1886 6010
rect 1938 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 2270 6010
rect 2322 5958 2334 6010
rect 2386 5958 2398 6010
rect 2450 5958 2462 6010
rect 2514 5958 2526 6010
rect 2578 5958 2590 6010
rect 2642 5958 2654 6010
rect 2706 5958 9502 6010
rect 9554 5958 9566 6010
rect 9618 5958 9630 6010
rect 9682 5958 9694 6010
rect 9746 5958 9758 6010
rect 9810 5958 9822 6010
rect 9874 5958 9886 6010
rect 9938 5958 9950 6010
rect 10002 5958 10014 6010
rect 10066 5958 10078 6010
rect 10130 5958 10142 6010
rect 10194 5958 10206 6010
rect 10258 5958 10270 6010
rect 10322 5958 10334 6010
rect 10386 5958 10398 6010
rect 10450 5958 10462 6010
rect 10514 5958 10526 6010
rect 10578 5958 10590 6010
rect 10642 5958 10654 6010
rect 10706 5958 17502 6010
rect 17554 5958 17566 6010
rect 17618 5958 17630 6010
rect 17682 5958 17694 6010
rect 17746 5958 17758 6010
rect 17810 5958 17822 6010
rect 17874 5958 17886 6010
rect 17938 5958 17950 6010
rect 18002 5958 18014 6010
rect 18066 5958 18078 6010
rect 18130 5958 18142 6010
rect 18194 5958 18206 6010
rect 18258 5958 18270 6010
rect 18322 5958 18334 6010
rect 18386 5958 18398 6010
rect 18450 5958 18462 6010
rect 18514 5958 18526 6010
rect 18578 5958 18590 6010
rect 18642 5958 18654 6010
rect 18706 5958 18860 6010
rect 1104 5936 18860 5958
rect 3602 5896 3608 5908
rect 2148 5868 3608 5896
rect 2148 5701 2176 5868
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 4948 5868 8248 5896
rect 4948 5856 4954 5868
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 2866 5828 2872 5840
rect 2823 5800 2872 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 2866 5788 2872 5800
rect 2924 5828 2930 5840
rect 4065 5831 4123 5837
rect 4065 5828 4077 5831
rect 2924 5800 4077 5828
rect 2924 5788 2930 5800
rect 4065 5797 4077 5800
rect 4111 5797 4123 5831
rect 4065 5791 4123 5797
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 4154 5760 4160 5772
rect 2731 5732 4160 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7745 5763 7803 5769
rect 7745 5760 7757 5763
rect 6972 5732 7757 5760
rect 6972 5720 6978 5732
rect 7745 5729 7757 5732
rect 7791 5760 7803 5763
rect 7834 5760 7840 5772
rect 7791 5732 7840 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 8220 5760 8248 5868
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 10321 5899 10379 5905
rect 10321 5896 10333 5899
rect 8352 5868 10333 5896
rect 8352 5856 8358 5868
rect 10321 5865 10333 5868
rect 10367 5896 10379 5899
rect 11422 5896 11428 5908
rect 10367 5868 11428 5896
rect 10367 5865 10379 5868
rect 10321 5859 10379 5865
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12250 5896 12256 5908
rect 12032 5868 12256 5896
rect 12032 5856 12038 5868
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 14366 5856 14372 5908
rect 14424 5856 14430 5908
rect 14476 5868 16620 5896
rect 12342 5788 12348 5840
rect 12400 5828 12406 5840
rect 14476 5828 14504 5868
rect 12400 5800 14504 5828
rect 12400 5788 12406 5800
rect 11146 5760 11152 5772
rect 8220 5732 11152 5760
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 11790 5720 11796 5772
rect 11848 5720 11854 5772
rect 12894 5720 12900 5772
rect 12952 5760 12958 5772
rect 12989 5763 13047 5769
rect 12989 5760 13001 5763
rect 12952 5732 13001 5760
rect 12952 5720 12958 5732
rect 12989 5729 13001 5732
rect 13035 5729 13047 5763
rect 12989 5723 13047 5729
rect 13078 5720 13084 5772
rect 13136 5760 13142 5772
rect 13173 5763 13231 5769
rect 13173 5760 13185 5763
rect 13136 5732 13185 5760
rect 13136 5720 13142 5732
rect 13173 5729 13185 5732
rect 13219 5760 13231 5763
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 13219 5732 14565 5760
rect 13219 5729 13231 5732
rect 13173 5723 13231 5729
rect 14553 5729 14565 5732
rect 14599 5760 14611 5763
rect 15102 5760 15108 5772
rect 14599 5732 15108 5760
rect 14599 5729 14611 5732
rect 14553 5723 14611 5729
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 15286 5720 15292 5772
rect 15344 5720 15350 5772
rect 15565 5763 15623 5769
rect 15565 5729 15577 5763
rect 15611 5760 15623 5763
rect 16022 5760 16028 5772
rect 15611 5732 16028 5760
rect 15611 5729 15623 5732
rect 15565 5723 15623 5729
rect 16022 5720 16028 5732
rect 16080 5720 16086 5772
rect 16592 5760 16620 5868
rect 17034 5856 17040 5908
rect 17092 5856 17098 5908
rect 17218 5856 17224 5908
rect 17276 5896 17282 5908
rect 17276 5868 18184 5896
rect 17276 5856 17282 5868
rect 17402 5788 17408 5840
rect 17460 5828 17466 5840
rect 18156 5837 18184 5868
rect 18141 5831 18199 5837
rect 17460 5800 17724 5828
rect 17460 5788 17466 5800
rect 16592 5732 17632 5760
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 2133 5695 2191 5701
rect 1627 5664 2084 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 1673 5627 1731 5633
rect 1673 5593 1685 5627
rect 1719 5593 1731 5627
rect 2056 5624 2084 5664
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3326 5692 3332 5704
rect 3283 5664 3332 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3436 5664 4077 5692
rect 2314 5624 2320 5636
rect 2056 5596 2320 5624
rect 1673 5587 1731 5593
rect 1688 5556 1716 5587
rect 2314 5584 2320 5596
rect 2372 5624 2378 5636
rect 3436 5624 3464 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 2372 5596 3464 5624
rect 2372 5584 2378 5596
rect 3510 5584 3516 5636
rect 3568 5624 3574 5636
rect 5552 5624 5580 5655
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 7282 5652 7288 5704
rect 7340 5652 7346 5704
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 8220 5664 9321 5692
rect 3568 5596 5580 5624
rect 6365 5627 6423 5633
rect 3568 5584 3574 5596
rect 6365 5593 6377 5627
rect 6411 5624 6423 5627
rect 7300 5624 7328 5652
rect 6411 5596 7328 5624
rect 6411 5593 6423 5596
rect 6365 5587 6423 5593
rect 8110 5584 8116 5636
rect 8168 5624 8174 5636
rect 8220 5633 8248 5664
rect 9309 5661 9321 5664
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 12066 5652 12072 5704
rect 12124 5652 12130 5704
rect 13354 5652 13360 5704
rect 13412 5692 13418 5704
rect 14734 5692 14740 5704
rect 13412 5664 14740 5692
rect 13412 5652 13418 5664
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5692 14887 5695
rect 15194 5692 15200 5704
rect 14875 5664 15200 5692
rect 14875 5661 14887 5664
rect 14829 5655 14887 5661
rect 15194 5652 15200 5664
rect 15252 5652 15258 5704
rect 17604 5701 17632 5732
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5661 17647 5695
rect 17696 5692 17724 5800
rect 18141 5797 18153 5831
rect 18187 5797 18199 5831
rect 18141 5791 18199 5797
rect 17819 5695 17877 5701
rect 17819 5692 17831 5695
rect 17696 5664 17831 5692
rect 17589 5655 17647 5661
rect 17819 5661 17831 5664
rect 17865 5661 17877 5695
rect 17819 5655 17877 5661
rect 8205 5627 8263 5633
rect 8205 5624 8217 5627
rect 8168 5596 8217 5624
rect 8168 5584 8174 5596
rect 8205 5593 8217 5596
rect 8251 5593 8263 5627
rect 8205 5587 8263 5593
rect 8297 5627 8355 5633
rect 8297 5593 8309 5627
rect 8343 5593 8355 5627
rect 8297 5587 8355 5593
rect 3050 5556 3056 5568
rect 1688 5528 3056 5556
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 7101 5559 7159 5565
rect 7101 5525 7113 5559
rect 7147 5556 7159 5559
rect 8312 5556 8340 5587
rect 9122 5584 9128 5636
rect 9180 5584 9186 5636
rect 14642 5624 14648 5636
rect 11362 5596 11560 5624
rect 7147 5528 8340 5556
rect 11532 5556 11560 5596
rect 11900 5596 14648 5624
rect 11900 5556 11928 5596
rect 14642 5584 14648 5596
rect 14700 5584 14706 5636
rect 14752 5624 14780 5652
rect 15470 5624 15476 5636
rect 14752 5596 15476 5624
rect 15470 5584 15476 5596
rect 15528 5584 15534 5636
rect 16114 5584 16120 5636
rect 16172 5584 16178 5636
rect 17957 5627 18015 5633
rect 17957 5624 17969 5627
rect 16868 5596 17969 5624
rect 11532 5528 11928 5556
rect 7147 5525 7159 5528
rect 7101 5519 7159 5525
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12529 5559 12587 5565
rect 12529 5556 12541 5559
rect 12032 5528 12541 5556
rect 12032 5516 12038 5528
rect 12529 5525 12541 5528
rect 12575 5525 12587 5559
rect 12529 5519 12587 5525
rect 12897 5559 12955 5565
rect 12897 5525 12909 5559
rect 12943 5556 12955 5559
rect 14550 5556 14556 5568
rect 12943 5528 14556 5556
rect 12943 5525 12955 5528
rect 12897 5519 12955 5525
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 14734 5516 14740 5568
rect 14792 5556 14798 5568
rect 16868 5556 16896 5596
rect 17957 5593 17969 5596
rect 18003 5593 18015 5627
rect 17957 5587 18015 5593
rect 14792 5528 16896 5556
rect 14792 5516 14798 5528
rect 16942 5516 16948 5568
rect 17000 5556 17006 5568
rect 17773 5559 17831 5565
rect 17773 5556 17785 5559
rect 17000 5528 17785 5556
rect 17000 5516 17006 5528
rect 17773 5525 17785 5528
rect 17819 5525 17831 5559
rect 17773 5519 17831 5525
rect 1104 5466 18860 5488
rect 1104 5414 5502 5466
rect 5554 5414 5566 5466
rect 5618 5414 5630 5466
rect 5682 5414 5694 5466
rect 5746 5414 5758 5466
rect 5810 5414 5822 5466
rect 5874 5414 5886 5466
rect 5938 5414 5950 5466
rect 6002 5414 6014 5466
rect 6066 5414 6078 5466
rect 6130 5414 6142 5466
rect 6194 5414 6206 5466
rect 6258 5414 6270 5466
rect 6322 5414 6334 5466
rect 6386 5414 6398 5466
rect 6450 5414 6462 5466
rect 6514 5414 6526 5466
rect 6578 5414 6590 5466
rect 6642 5414 6654 5466
rect 6706 5414 13502 5466
rect 13554 5414 13566 5466
rect 13618 5414 13630 5466
rect 13682 5414 13694 5466
rect 13746 5414 13758 5466
rect 13810 5414 13822 5466
rect 13874 5414 13886 5466
rect 13938 5414 13950 5466
rect 14002 5414 14014 5466
rect 14066 5414 14078 5466
rect 14130 5414 14142 5466
rect 14194 5414 14206 5466
rect 14258 5414 14270 5466
rect 14322 5414 14334 5466
rect 14386 5414 14398 5466
rect 14450 5414 14462 5466
rect 14514 5414 14526 5466
rect 14578 5414 14590 5466
rect 14642 5414 14654 5466
rect 14706 5414 18860 5466
rect 1104 5392 18860 5414
rect 4154 5312 4160 5364
rect 4212 5312 4218 5364
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 5629 5355 5687 5361
rect 5629 5352 5641 5355
rect 4396 5324 5641 5352
rect 4396 5312 4402 5324
rect 5629 5321 5641 5324
rect 5675 5321 5687 5355
rect 5629 5315 5687 5321
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 7374 5352 7380 5364
rect 5776 5324 7380 5352
rect 5776 5312 5782 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 8018 5352 8024 5364
rect 7616 5324 8024 5352
rect 7616 5312 7622 5324
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 12066 5312 12072 5364
rect 12124 5352 12130 5364
rect 12124 5324 13492 5352
rect 12124 5312 12130 5324
rect 3050 5244 3056 5296
rect 3108 5284 3114 5296
rect 4065 5287 4123 5293
rect 4065 5284 4077 5287
rect 3108 5256 4077 5284
rect 3108 5244 3114 5256
rect 4065 5253 4077 5256
rect 4111 5253 4123 5287
rect 4065 5247 4123 5253
rect 7009 5287 7067 5293
rect 7009 5253 7021 5287
rect 7055 5284 7067 5287
rect 8110 5284 8116 5296
rect 7055 5256 8116 5284
rect 7055 5253 7067 5256
rect 7009 5247 7067 5253
rect 8110 5244 8116 5256
rect 8168 5244 8174 5296
rect 8205 5287 8263 5293
rect 8205 5253 8217 5287
rect 8251 5284 8263 5287
rect 9122 5284 9128 5296
rect 8251 5256 9128 5284
rect 8251 5253 8263 5256
rect 8205 5247 8263 5253
rect 9122 5244 9128 5256
rect 9180 5244 9186 5296
rect 11974 5244 11980 5296
rect 12032 5244 12038 5296
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 12308 5256 12466 5284
rect 12308 5244 12314 5256
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 2314 5216 2320 5228
rect 1903 5188 2320 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 1688 5148 1716 5179
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5216 3571 5219
rect 3602 5216 3608 5228
rect 3559 5188 3608 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4890 5176 4896 5228
rect 4948 5216 4954 5228
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 4948 5188 5273 5216
rect 4948 5176 4954 5188
rect 5261 5185 5273 5188
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 5517 5219 5575 5225
rect 5517 5185 5529 5219
rect 5563 5216 5575 5219
rect 6454 5216 6460 5228
rect 5563 5188 6460 5216
rect 5563 5185 5575 5188
rect 5517 5179 5575 5185
rect 6454 5176 6460 5188
rect 6512 5176 6518 5228
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6914 5216 6920 5228
rect 6595 5188 6920 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7282 5216 7288 5228
rect 7147 5188 7288 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7282 5176 7288 5188
rect 7340 5216 7346 5228
rect 7340 5188 7788 5216
rect 7340 5176 7346 5188
rect 2774 5148 2780 5160
rect 1688 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 2961 5151 3019 5157
rect 2961 5117 2973 5151
rect 3007 5117 3019 5151
rect 2961 5111 3019 5117
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6730 5148 6736 5160
rect 5859 5120 6736 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 2501 5083 2559 5089
rect 2501 5049 2513 5083
rect 2547 5080 2559 5083
rect 2976 5080 3004 5111
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 7558 5108 7564 5160
rect 7616 5148 7622 5160
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 7616 5120 7665 5148
rect 7616 5108 7622 5120
rect 7653 5117 7665 5120
rect 7699 5117 7711 5151
rect 7760 5148 7788 5188
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8076 5188 8953 5216
rect 8076 5176 8082 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5185 9919 5219
rect 13464 5216 13492 5324
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 15749 5355 15807 5361
rect 15749 5352 15761 5355
rect 14608 5324 15761 5352
rect 14608 5312 14614 5324
rect 15749 5321 15761 5324
rect 15795 5352 15807 5355
rect 15838 5352 15844 5364
rect 15795 5324 15844 5352
rect 15795 5321 15807 5324
rect 15749 5315 15807 5321
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 16666 5312 16672 5364
rect 16724 5352 16730 5364
rect 17218 5352 17224 5364
rect 16724 5324 17224 5352
rect 16724 5312 16730 5324
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 19702 5352 19708 5364
rect 17788 5324 19708 5352
rect 17788 5284 17816 5324
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 15502 5256 17816 5284
rect 17862 5244 17868 5296
rect 17920 5244 17926 5296
rect 18049 5287 18107 5293
rect 18049 5253 18061 5287
rect 18095 5253 18107 5287
rect 18049 5247 18107 5253
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13464 5188 14013 5216
rect 9861 5179 9919 5185
rect 14001 5185 14013 5188
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 9876 5148 9904 5179
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16540 5188 16957 5216
rect 16540 5176 16546 5188
rect 16945 5185 16957 5188
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 17034 5176 17040 5228
rect 17092 5216 17098 5228
rect 18064 5216 18092 5247
rect 17092 5188 18092 5216
rect 17092 5176 17098 5188
rect 7760 5120 9904 5148
rect 7653 5111 7711 5117
rect 11606 5108 11612 5160
rect 11664 5148 11670 5160
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 11664 5120 11713 5148
rect 11664 5108 11670 5120
rect 11701 5117 11713 5120
rect 11747 5148 11759 5151
rect 12066 5148 12072 5160
rect 11747 5120 12072 5148
rect 11747 5117 11759 5120
rect 11701 5111 11759 5117
rect 12066 5108 12072 5120
rect 12124 5108 12130 5160
rect 12986 5108 12992 5160
rect 13044 5148 13050 5160
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 13044 5120 13461 5148
rect 13044 5108 13050 5120
rect 13449 5117 13461 5120
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 14274 5108 14280 5160
rect 14332 5108 14338 5160
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 17221 5151 17279 5157
rect 17221 5148 17233 5151
rect 15528 5120 17233 5148
rect 15528 5108 15534 5120
rect 17221 5117 17233 5120
rect 17267 5117 17279 5151
rect 17221 5111 17279 5117
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 18046 5148 18052 5160
rect 17368 5120 18052 5148
rect 17368 5108 17374 5120
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 2547 5052 3004 5080
rect 2547 5049 2559 5052
rect 2501 5043 2559 5049
rect 6546 5040 6552 5092
rect 6604 5080 6610 5092
rect 8113 5083 8171 5089
rect 8113 5080 8125 5083
rect 6604 5052 8125 5080
rect 6604 5040 6610 5052
rect 8113 5049 8125 5052
rect 8159 5080 8171 5083
rect 10229 5083 10287 5089
rect 10229 5080 10241 5083
rect 8159 5052 10241 5080
rect 8159 5049 8171 5052
rect 8113 5043 8171 5049
rect 10229 5049 10241 5052
rect 10275 5049 10287 5083
rect 10229 5043 10287 5049
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 18233 5083 18291 5089
rect 18233 5080 18245 5083
rect 16632 5052 18245 5080
rect 16632 5040 16638 5052
rect 18233 5049 18245 5052
rect 18279 5049 18291 5083
rect 18233 5043 18291 5049
rect 5261 5015 5319 5021
rect 5261 4981 5273 5015
rect 5307 5012 5319 5015
rect 6730 5012 6736 5024
rect 5307 4984 6736 5012
rect 5307 4981 5319 4984
rect 5261 4975 5319 4981
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 14826 5012 14832 5024
rect 8536 4984 14832 5012
rect 8536 4972 8542 4984
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 15286 4972 15292 5024
rect 15344 5012 15350 5024
rect 17037 5015 17095 5021
rect 17037 5012 17049 5015
rect 15344 4984 17049 5012
rect 15344 4972 15350 4984
rect 17037 4981 17049 4984
rect 17083 4981 17095 5015
rect 17037 4975 17095 4981
rect 17218 4972 17224 5024
rect 17276 5012 17282 5024
rect 17862 5012 17868 5024
rect 17276 4984 17868 5012
rect 17276 4972 17282 4984
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18046 4972 18052 5024
rect 18104 4972 18110 5024
rect 1104 4922 18860 4944
rect 1104 4870 1502 4922
rect 1554 4870 1566 4922
rect 1618 4870 1630 4922
rect 1682 4870 1694 4922
rect 1746 4870 1758 4922
rect 1810 4870 1822 4922
rect 1874 4870 1886 4922
rect 1938 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 2270 4922
rect 2322 4870 2334 4922
rect 2386 4870 2398 4922
rect 2450 4870 2462 4922
rect 2514 4870 2526 4922
rect 2578 4870 2590 4922
rect 2642 4870 2654 4922
rect 2706 4870 9502 4922
rect 9554 4870 9566 4922
rect 9618 4870 9630 4922
rect 9682 4870 9694 4922
rect 9746 4870 9758 4922
rect 9810 4870 9822 4922
rect 9874 4870 9886 4922
rect 9938 4870 9950 4922
rect 10002 4870 10014 4922
rect 10066 4870 10078 4922
rect 10130 4870 10142 4922
rect 10194 4870 10206 4922
rect 10258 4870 10270 4922
rect 10322 4870 10334 4922
rect 10386 4870 10398 4922
rect 10450 4870 10462 4922
rect 10514 4870 10526 4922
rect 10578 4870 10590 4922
rect 10642 4870 10654 4922
rect 10706 4870 17502 4922
rect 17554 4870 17566 4922
rect 17618 4870 17630 4922
rect 17682 4870 17694 4922
rect 17746 4870 17758 4922
rect 17810 4870 17822 4922
rect 17874 4870 17886 4922
rect 17938 4870 17950 4922
rect 18002 4870 18014 4922
rect 18066 4870 18078 4922
rect 18130 4870 18142 4922
rect 18194 4870 18206 4922
rect 18258 4870 18270 4922
rect 18322 4870 18334 4922
rect 18386 4870 18398 4922
rect 18450 4870 18462 4922
rect 18514 4870 18526 4922
rect 18578 4870 18590 4922
rect 18642 4870 18654 4922
rect 18706 4870 18860 4922
rect 1104 4848 18860 4870
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 14642 4808 14648 4820
rect 8076 4780 14648 4808
rect 8076 4768 8082 4780
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 16298 4808 16304 4820
rect 14752 4780 16304 4808
rect 5258 4700 5264 4752
rect 5316 4740 5322 4752
rect 6914 4740 6920 4752
rect 5316 4712 6920 4740
rect 5316 4700 5322 4712
rect 6914 4700 6920 4712
rect 6972 4700 6978 4752
rect 12069 4743 12127 4749
rect 12069 4709 12081 4743
rect 12115 4709 12127 4743
rect 12069 4703 12127 4709
rect 1210 4632 1216 4684
rect 1268 4672 1274 4684
rect 1765 4675 1823 4681
rect 1268 4644 1716 4672
rect 1268 4632 1274 4644
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4573 1639 4607
rect 1688 4604 1716 4644
rect 1765 4641 1777 4675
rect 1811 4672 1823 4675
rect 3050 4672 3056 4684
rect 1811 4644 3056 4672
rect 1811 4641 1823 4644
rect 1765 4635 1823 4641
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3970 4672 3976 4684
rect 3283 4644 3976 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 3970 4632 3976 4644
rect 4028 4672 4034 4684
rect 4028 4644 5580 4672
rect 4028 4632 4034 4644
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 1688 4576 2145 4604
rect 1581 4567 1639 4573
rect 2133 4573 2145 4576
rect 2179 4604 2191 4607
rect 3142 4604 3148 4616
rect 2179 4576 3148 4604
rect 2179 4573 2191 4576
rect 2133 4567 2191 4573
rect 1596 4536 1624 4567
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 5552 4613 5580 4644
rect 6730 4632 6736 4684
rect 6788 4672 6794 4684
rect 7745 4675 7803 4681
rect 7745 4672 7757 4675
rect 6788 4644 7757 4672
rect 6788 4632 6794 4644
rect 7745 4641 7757 4644
rect 7791 4641 7803 4675
rect 7745 4635 7803 4641
rect 8202 4632 8208 4684
rect 8260 4672 8266 4684
rect 9217 4675 9275 4681
rect 9217 4672 9229 4675
rect 8260 4644 9229 4672
rect 8260 4632 8266 4644
rect 9217 4641 9229 4644
rect 9263 4641 9275 4675
rect 9217 4635 9275 4641
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 12084 4672 12112 4703
rect 13354 4700 13360 4752
rect 13412 4700 13418 4752
rect 14274 4700 14280 4752
rect 14332 4700 14338 4752
rect 11379 4644 12112 4672
rect 12713 4675 12771 4681
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 12713 4641 12725 4675
rect 12759 4672 12771 4675
rect 13078 4672 13084 4684
rect 12759 4644 13084 4672
rect 12759 4641 12771 4644
rect 12713 4635 12771 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 14752 4672 14780 4780
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 16850 4768 16856 4820
rect 16908 4808 16914 4820
rect 17129 4811 17187 4817
rect 17129 4808 17141 4811
rect 16908 4780 17141 4808
rect 16908 4768 16914 4780
rect 17129 4777 17141 4780
rect 17175 4777 17187 4811
rect 17129 4771 17187 4777
rect 17402 4700 17408 4752
rect 17460 4740 17466 4752
rect 17773 4743 17831 4749
rect 17773 4740 17785 4743
rect 17460 4712 17785 4740
rect 17460 4700 17466 4712
rect 17773 4709 17785 4712
rect 17819 4709 17831 4743
rect 17773 4703 17831 4709
rect 15286 4672 15292 4684
rect 13464 4644 14780 4672
rect 14844 4644 15292 4672
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 1596 4508 2360 4536
rect 2332 4480 2360 4508
rect 2682 4496 2688 4548
rect 2740 4496 2746 4548
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 3973 4539 4031 4545
rect 3973 4536 3985 4539
rect 2832 4508 3985 4536
rect 2832 4496 2838 4508
rect 3973 4505 3985 4508
rect 4019 4505 4031 4539
rect 3973 4499 4031 4505
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 4080 4468 4108 4567
rect 6546 4564 6552 4616
rect 6604 4564 6610 4616
rect 7282 4564 7288 4616
rect 7340 4564 7346 4616
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 8220 4576 9321 4604
rect 6365 4539 6423 4545
rect 6365 4505 6377 4539
rect 6411 4536 6423 4539
rect 7300 4536 7328 4564
rect 6411 4508 7328 4536
rect 6411 4505 6423 4508
rect 6365 4499 6423 4505
rect 8110 4496 8116 4548
rect 8168 4536 8174 4548
rect 8220 4545 8248 4576
rect 9309 4573 9321 4576
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 11606 4564 11612 4616
rect 11664 4564 11670 4616
rect 8205 4539 8263 4545
rect 8205 4536 8217 4539
rect 8168 4508 8217 4536
rect 8168 4496 8174 4508
rect 8205 4505 8217 4508
rect 8251 4505 8263 4539
rect 8205 4499 8263 4505
rect 8297 4539 8355 4545
rect 8297 4505 8309 4539
rect 8343 4505 8355 4539
rect 8297 4499 8355 4505
rect 2372 4440 4108 4468
rect 2372 4428 2378 4440
rect 5074 4428 5080 4480
rect 5132 4468 5138 4480
rect 5718 4468 5724 4480
rect 5132 4440 5724 4468
rect 5132 4428 5138 4440
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 7101 4471 7159 4477
rect 7101 4437 7113 4471
rect 7147 4468 7159 4471
rect 8312 4468 8340 4499
rect 10686 4496 10692 4548
rect 10744 4496 10750 4548
rect 12529 4539 12587 4545
rect 12529 4536 12541 4539
rect 11341 4508 12541 4536
rect 7147 4440 8340 4468
rect 9861 4471 9919 4477
rect 7147 4437 7159 4440
rect 7101 4431 7159 4437
rect 9861 4437 9873 4471
rect 9907 4468 9919 4471
rect 11341 4468 11369 4508
rect 12529 4505 12541 4508
rect 12575 4536 12587 4539
rect 13464 4536 13492 4644
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 14550 4604 14556 4616
rect 13771 4576 14556 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 12575 4508 13492 4536
rect 13556 4536 13584 4567
rect 14550 4564 14556 4576
rect 14608 4564 14614 4616
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4573 14703 4607
rect 14645 4567 14703 4573
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4604 14795 4607
rect 14844 4604 14872 4644
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 15378 4632 15384 4684
rect 15436 4632 15442 4684
rect 15654 4632 15660 4684
rect 15712 4632 15718 4684
rect 16666 4632 16672 4684
rect 16724 4672 16730 4684
rect 18233 4675 18291 4681
rect 18233 4672 18245 4675
rect 16724 4644 18245 4672
rect 16724 4632 16730 4644
rect 18233 4641 18245 4644
rect 18279 4641 18291 4675
rect 18233 4635 18291 4641
rect 14783 4576 14872 4604
rect 14921 4607 14979 4613
rect 14783 4573 14795 4576
rect 14737 4567 14795 4573
rect 14921 4573 14933 4607
rect 14967 4604 14979 4607
rect 15102 4604 15108 4616
rect 14967 4576 15108 4604
rect 14967 4573 14979 4576
rect 14921 4567 14979 4573
rect 14660 4536 14688 4567
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 16758 4564 16764 4616
rect 16816 4564 16822 4616
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4604 17739 4607
rect 18049 4607 18107 4613
rect 17727 4576 18000 4604
rect 17727 4573 17739 4576
rect 17681 4567 17739 4573
rect 15120 4536 15148 4564
rect 15562 4536 15568 4548
rect 13556 4508 14780 4536
rect 15120 4508 15568 4536
rect 12575 4505 12587 4508
rect 12529 4499 12587 4505
rect 9907 4440 11369 4468
rect 9907 4437 9919 4440
rect 9861 4431 9919 4437
rect 11882 4428 11888 4480
rect 11940 4468 11946 4480
rect 12342 4468 12348 4480
rect 11940 4440 12348 4468
rect 11940 4428 11946 4440
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 12434 4428 12440 4480
rect 12492 4428 12498 4480
rect 14752 4468 14780 4508
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 16574 4468 16580 4480
rect 14752 4440 16580 4468
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 17972 4468 18000 4576
rect 18049 4573 18061 4607
rect 18095 4573 18107 4607
rect 18049 4567 18107 4573
rect 18064 4536 18092 4567
rect 18782 4536 18788 4548
rect 18064 4508 18788 4536
rect 18782 4496 18788 4508
rect 18840 4496 18846 4548
rect 19426 4468 19432 4480
rect 17972 4440 19432 4468
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 1104 4378 18860 4400
rect 1104 4326 5502 4378
rect 5554 4326 5566 4378
rect 5618 4326 5630 4378
rect 5682 4326 5694 4378
rect 5746 4326 5758 4378
rect 5810 4326 5822 4378
rect 5874 4326 5886 4378
rect 5938 4326 5950 4378
rect 6002 4326 6014 4378
rect 6066 4326 6078 4378
rect 6130 4326 6142 4378
rect 6194 4326 6206 4378
rect 6258 4326 6270 4378
rect 6322 4326 6334 4378
rect 6386 4326 6398 4378
rect 6450 4326 6462 4378
rect 6514 4326 6526 4378
rect 6578 4326 6590 4378
rect 6642 4326 6654 4378
rect 6706 4326 13502 4378
rect 13554 4326 13566 4378
rect 13618 4326 13630 4378
rect 13682 4326 13694 4378
rect 13746 4326 13758 4378
rect 13810 4326 13822 4378
rect 13874 4326 13886 4378
rect 13938 4326 13950 4378
rect 14002 4326 14014 4378
rect 14066 4326 14078 4378
rect 14130 4326 14142 4378
rect 14194 4326 14206 4378
rect 14258 4326 14270 4378
rect 14322 4326 14334 4378
rect 14386 4326 14398 4378
rect 14450 4326 14462 4378
rect 14514 4326 14526 4378
rect 14578 4326 14590 4378
rect 14642 4326 14654 4378
rect 14706 4326 18860 4378
rect 1104 4304 18860 4326
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 4157 4267 4215 4273
rect 4157 4264 4169 4267
rect 2740 4236 4169 4264
rect 2740 4224 2746 4236
rect 4157 4233 4169 4236
rect 4203 4233 4215 4267
rect 4157 4227 4215 4233
rect 6822 4224 6828 4276
rect 6880 4264 6886 4276
rect 7926 4264 7932 4276
rect 6880 4236 7932 4264
rect 6880 4224 6886 4236
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 11204 4236 12173 4264
rect 11204 4224 11210 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 12161 4227 12219 4233
rect 14734 4224 14740 4276
rect 14792 4264 14798 4276
rect 15289 4267 15347 4273
rect 15289 4264 15301 4267
rect 14792 4236 15301 4264
rect 14792 4224 14798 4236
rect 15289 4233 15301 4236
rect 15335 4233 15347 4267
rect 15289 4227 15347 4233
rect 1673 4199 1731 4205
rect 1673 4165 1685 4199
rect 1719 4196 1731 4199
rect 1719 4168 2774 4196
rect 1719 4165 1731 4168
rect 1673 4159 1731 4165
rect 2746 4140 2774 4168
rect 3050 4156 3056 4208
rect 3108 4196 3114 4208
rect 4065 4199 4123 4205
rect 4065 4196 4077 4199
rect 3108 4168 4077 4196
rect 3108 4156 3114 4168
rect 4065 4165 4077 4168
rect 4111 4165 4123 4199
rect 4065 4159 4123 4165
rect 5169 4199 5227 4205
rect 5169 4165 5181 4199
rect 5215 4196 5227 4199
rect 5718 4196 5724 4208
rect 5215 4168 5724 4196
rect 5215 4165 5227 4168
rect 5169 4159 5227 4165
rect 5718 4156 5724 4168
rect 5776 4156 5782 4208
rect 6638 4196 6644 4208
rect 5828 4168 6644 4196
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 2314 4128 2320 4140
rect 1903 4100 2320 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2746 4100 2780 4140
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3513 4131 3571 4137
rect 3513 4128 3525 4131
rect 3200 4100 3525 4128
rect 3200 4088 3206 4100
rect 3513 4097 3525 4100
rect 3559 4097 3571 4131
rect 5828 4114 5856 4168
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 7009 4199 7067 4205
rect 7009 4165 7021 4199
rect 7055 4196 7067 4199
rect 8110 4196 8116 4208
rect 7055 4168 8116 4196
rect 7055 4165 7067 4168
rect 7009 4159 7067 4165
rect 8110 4156 8116 4168
rect 8168 4156 8174 4208
rect 8202 4156 8208 4208
rect 8260 4156 8266 4208
rect 12434 4156 12440 4208
rect 12492 4196 12498 4208
rect 12492 4168 14780 4196
rect 12492 4156 12498 4168
rect 6549 4131 6607 4137
rect 3513 4091 3571 4097
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6730 4128 6736 4140
rect 6595 4100 6736 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7282 4128 7288 4140
rect 7147 4100 7288 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 7760 4100 8953 4128
rect 2961 4063 3019 4069
rect 2961 4060 2973 4063
rect 2746 4032 2973 4060
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3992 2559 3995
rect 2746 3992 2774 4032
rect 2961 4029 2973 4032
rect 3007 4029 3019 4063
rect 2961 4023 3019 4029
rect 4982 4020 4988 4072
rect 5040 4060 5046 4072
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 5040 4032 5733 4060
rect 5040 4020 5046 4032
rect 5721 4029 5733 4032
rect 5767 4029 5779 4063
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 5721 4023 5779 4029
rect 7024 4032 7665 4060
rect 7024 3992 7052 4032
rect 7653 4029 7665 4032
rect 7699 4060 7711 4063
rect 7760 4060 7788 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 9876 4060 9904 4091
rect 7699 4032 7788 4060
rect 7852 4032 9904 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 2547 3964 2774 3992
rect 5736 3964 7052 3992
rect 2547 3961 2559 3964
rect 2501 3955 2559 3961
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 5736 3924 5764 3964
rect 7282 3952 7288 4004
rect 7340 3992 7346 4004
rect 7852 3992 7880 4032
rect 7340 3964 7880 3992
rect 8113 3995 8171 4001
rect 7340 3952 7346 3964
rect 8113 3961 8125 3995
rect 8159 3992 8171 3995
rect 10229 3995 10287 4001
rect 10229 3992 10241 3995
rect 8159 3964 10241 3992
rect 8159 3961 8171 3964
rect 8113 3955 8171 3961
rect 10229 3961 10241 3964
rect 10275 3961 10287 3995
rect 10229 3955 10287 3961
rect 1452 3896 5764 3924
rect 1452 3884 1458 3896
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 8128 3924 8156 3955
rect 6144 3896 8156 3924
rect 6144 3884 6150 3896
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 10980 3924 11008 4091
rect 11514 4088 11520 4140
rect 11572 4128 11578 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11572 4100 11713 4128
rect 11572 4088 11578 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11848 4100 11897 4128
rect 11848 4088 11854 4100
rect 11885 4097 11897 4100
rect 11931 4128 11943 4131
rect 12066 4128 12072 4140
rect 11931 4100 12072 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12176 4100 12434 4128
rect 12176 4060 12204 4100
rect 11348 4032 12204 4060
rect 11348 3936 11376 4032
rect 12250 4020 12256 4072
rect 12308 4020 12314 4072
rect 12406 4060 12434 4100
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 13541 4131 13599 4137
rect 13541 4128 13553 4131
rect 13412 4100 13553 4128
rect 13412 4088 13418 4100
rect 13541 4097 13553 4100
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 14752 4128 14780 4168
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 15010 4196 15016 4208
rect 14884 4168 15016 4196
rect 14884 4156 14890 4168
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 17034 4196 17040 4208
rect 15304 4168 17040 4196
rect 15304 4128 15332 4168
rect 17034 4156 17040 4168
rect 17092 4196 17098 4208
rect 17218 4196 17224 4208
rect 17092 4168 17224 4196
rect 17092 4156 17098 4168
rect 17218 4156 17224 4168
rect 17276 4156 17282 4208
rect 14752 4100 15332 4128
rect 14001 4091 14059 4097
rect 13170 4060 13176 4072
rect 12406 4032 13176 4060
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13262 4020 13268 4072
rect 13320 4020 13326 4072
rect 14016 4060 14044 4091
rect 16850 4088 16856 4140
rect 16908 4128 16914 4140
rect 17129 4131 17187 4137
rect 17129 4128 17141 4131
rect 16908 4100 17141 4128
rect 16908 4088 16914 4100
rect 17129 4097 17141 4100
rect 17175 4097 17187 4131
rect 17129 4091 17187 4097
rect 17310 4088 17316 4140
rect 17368 4088 17374 4140
rect 18141 4131 18199 4137
rect 18141 4097 18153 4131
rect 18187 4128 18199 4131
rect 18874 4128 18880 4140
rect 18187 4100 18880 4128
rect 18187 4097 18199 4100
rect 18141 4091 18199 4097
rect 18874 4088 18880 4100
rect 18932 4088 18938 4140
rect 15010 4060 15016 4072
rect 14016 4032 15016 4060
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 15194 4020 15200 4072
rect 15252 4060 15258 4072
rect 15381 4063 15439 4069
rect 15381 4060 15393 4063
rect 15252 4032 15393 4060
rect 15252 4020 15258 4032
rect 15381 4029 15393 4032
rect 15427 4029 15439 4063
rect 15381 4023 15439 4029
rect 15562 4020 15568 4072
rect 15620 4020 15626 4072
rect 11882 3952 11888 4004
rect 11940 3992 11946 4004
rect 16942 3992 16948 4004
rect 11940 3964 16948 3992
rect 11940 3952 11946 3964
rect 16942 3952 16948 3964
rect 17000 3952 17006 4004
rect 17126 3952 17132 4004
rect 17184 3992 17190 4004
rect 18874 3992 18880 4004
rect 17184 3964 18880 3992
rect 17184 3952 17190 3964
rect 18874 3952 18880 3964
rect 18932 3952 18938 4004
rect 8904 3896 11008 3924
rect 11057 3927 11115 3933
rect 8904 3884 8910 3896
rect 11057 3893 11069 3927
rect 11103 3924 11115 3927
rect 11330 3924 11336 3936
rect 11103 3896 11336 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 14921 3927 14979 3933
rect 14921 3924 14933 3927
rect 14792 3896 14933 3924
rect 14792 3884 14798 3896
rect 14921 3893 14933 3896
rect 14967 3893 14979 3927
rect 14921 3887 14979 3893
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 17310 3924 17316 3936
rect 15068 3896 17316 3924
rect 15068 3884 15074 3896
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 1104 3834 18860 3856
rect 1104 3782 1502 3834
rect 1554 3782 1566 3834
rect 1618 3782 1630 3834
rect 1682 3782 1694 3834
rect 1746 3782 1758 3834
rect 1810 3782 1822 3834
rect 1874 3782 1886 3834
rect 1938 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 2270 3834
rect 2322 3782 2334 3834
rect 2386 3782 2398 3834
rect 2450 3782 2462 3834
rect 2514 3782 2526 3834
rect 2578 3782 2590 3834
rect 2642 3782 2654 3834
rect 2706 3782 9502 3834
rect 9554 3782 9566 3834
rect 9618 3782 9630 3834
rect 9682 3782 9694 3834
rect 9746 3782 9758 3834
rect 9810 3782 9822 3834
rect 9874 3782 9886 3834
rect 9938 3782 9950 3834
rect 10002 3782 10014 3834
rect 10066 3782 10078 3834
rect 10130 3782 10142 3834
rect 10194 3782 10206 3834
rect 10258 3782 10270 3834
rect 10322 3782 10334 3834
rect 10386 3782 10398 3834
rect 10450 3782 10462 3834
rect 10514 3782 10526 3834
rect 10578 3782 10590 3834
rect 10642 3782 10654 3834
rect 10706 3782 17502 3834
rect 17554 3782 17566 3834
rect 17618 3782 17630 3834
rect 17682 3782 17694 3834
rect 17746 3782 17758 3834
rect 17810 3782 17822 3834
rect 17874 3782 17886 3834
rect 17938 3782 17950 3834
rect 18002 3782 18014 3834
rect 18066 3782 18078 3834
rect 18130 3782 18142 3834
rect 18194 3782 18206 3834
rect 18258 3782 18270 3834
rect 18322 3782 18334 3834
rect 18386 3782 18398 3834
rect 18450 3782 18462 3834
rect 18514 3782 18526 3834
rect 18578 3782 18590 3834
rect 18642 3782 18654 3834
rect 18706 3782 18860 3834
rect 1104 3760 18860 3782
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 6086 3720 6092 3732
rect 4028 3692 6092 3720
rect 4028 3680 4034 3692
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 8297 3723 8355 3729
rect 8297 3720 8309 3723
rect 6880 3692 8309 3720
rect 6880 3680 6886 3692
rect 8297 3689 8309 3692
rect 8343 3689 8355 3723
rect 8297 3683 8355 3689
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 9398 3720 9404 3732
rect 8812 3692 9404 3720
rect 8812 3680 8818 3692
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 11974 3720 11980 3732
rect 10744 3692 11980 3720
rect 10744 3680 10750 3692
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13228 3692 18000 3720
rect 13228 3680 13234 3692
rect 198 3612 204 3664
rect 256 3652 262 3664
rect 934 3652 940 3664
rect 256 3624 940 3652
rect 256 3612 262 3624
rect 934 3612 940 3624
rect 992 3612 998 3664
rect 1394 3612 1400 3664
rect 1452 3652 1458 3664
rect 2774 3652 2780 3664
rect 1452 3624 2780 3652
rect 1452 3612 1458 3624
rect 2774 3612 2780 3624
rect 2832 3652 2838 3664
rect 4249 3655 4307 3661
rect 4249 3652 4261 3655
rect 2832 3624 4261 3652
rect 2832 3612 2838 3624
rect 4249 3621 4261 3624
rect 4295 3652 4307 3655
rect 4798 3652 4804 3664
rect 4295 3624 4804 3652
rect 4295 3621 4307 3624
rect 4249 3615 4307 3621
rect 4798 3612 4804 3624
rect 4856 3612 4862 3664
rect 7745 3655 7803 3661
rect 7745 3621 7757 3655
rect 7791 3652 7803 3655
rect 8478 3652 8484 3664
rect 7791 3624 8484 3652
rect 7791 3621 7803 3624
rect 7745 3615 7803 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 9214 3612 9220 3664
rect 9272 3612 9278 3664
rect 9769 3655 9827 3661
rect 9769 3621 9781 3655
rect 9815 3652 9827 3655
rect 10410 3652 10416 3664
rect 9815 3624 10416 3652
rect 9815 3621 9827 3624
rect 9769 3615 9827 3621
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 10560 3624 12020 3652
rect 10560 3612 10566 3624
rect 290 3544 296 3596
rect 348 3584 354 3596
rect 4706 3584 4712 3596
rect 348 3556 3280 3584
rect 348 3544 354 3556
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 2866 3516 2872 3528
rect 2179 3488 2872 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 1596 3392 1624 3479
rect 2866 3476 2872 3488
rect 2924 3516 2930 3528
rect 3252 3525 3280 3556
rect 3436 3556 4712 3584
rect 3237 3519 3295 3525
rect 2924 3488 3188 3516
rect 2924 3476 2930 3488
rect 1673 3451 1731 3457
rect 1673 3417 1685 3451
rect 1719 3448 1731 3451
rect 2406 3448 2412 3460
rect 1719 3420 2412 3448
rect 1719 3417 1731 3420
rect 1673 3411 1731 3417
rect 2406 3408 2412 3420
rect 2464 3408 2470 3460
rect 2682 3408 2688 3460
rect 2740 3408 2746 3460
rect 3160 3448 3188 3488
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3326 3516 3332 3528
rect 3283 3488 3332 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 3436 3448 3464 3556
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 7006 3584 7012 3596
rect 6012 3556 7012 3584
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 4028 3488 4077 3516
rect 4028 3476 4034 3488
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 6012 3525 6040 3556
rect 7006 3544 7012 3556
rect 7064 3584 7070 3596
rect 11606 3584 11612 3596
rect 7064 3556 11612 3584
rect 7064 3544 7070 3556
rect 11606 3544 11612 3556
rect 11664 3584 11670 3596
rect 11885 3587 11943 3593
rect 11885 3584 11897 3587
rect 11664 3556 11897 3584
rect 11664 3544 11670 3556
rect 11885 3553 11897 3556
rect 11931 3553 11943 3587
rect 11992 3584 12020 3624
rect 13354 3612 13360 3664
rect 13412 3652 13418 3664
rect 13633 3655 13691 3661
rect 13633 3652 13645 3655
rect 13412 3624 13645 3652
rect 13412 3612 13418 3624
rect 13633 3621 13645 3624
rect 13679 3621 13691 3655
rect 13633 3615 13691 3621
rect 14642 3612 14648 3664
rect 14700 3652 14706 3664
rect 15102 3652 15108 3664
rect 14700 3624 15108 3652
rect 14700 3612 14706 3624
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 16684 3624 17908 3652
rect 16684 3584 16712 3624
rect 11992 3556 16712 3584
rect 11885 3547 11943 3553
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 17092 3556 17141 3584
rect 17092 3544 17098 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 17310 3544 17316 3596
rect 17368 3584 17374 3596
rect 17773 3587 17831 3593
rect 17773 3584 17785 3587
rect 17368 3556 17785 3584
rect 17368 3544 17374 3556
rect 17773 3553 17785 3556
rect 17819 3553 17831 3587
rect 17773 3547 17831 3553
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 4212 3488 5549 3516
rect 4212 3476 4218 3488
rect 5537 3485 5549 3488
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3485 6055 3519
rect 5997 3479 6055 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3516 8539 3519
rect 8570 3516 8576 3528
rect 8527 3488 8576 3516
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 3160 3420 3464 3448
rect 1578 3340 1584 3392
rect 1636 3380 1642 3392
rect 3988 3380 4016 3476
rect 5350 3408 5356 3460
rect 5408 3448 5414 3460
rect 6012 3448 6040 3479
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 5408 3420 6040 3448
rect 6273 3451 6331 3457
rect 5408 3408 5414 3420
rect 6273 3417 6285 3451
rect 6319 3417 6331 3451
rect 7742 3448 7748 3460
rect 7498 3420 7748 3448
rect 6273 3411 6331 3417
rect 1636 3352 4016 3380
rect 1636 3340 1642 3352
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 6288 3380 6316 3411
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 7834 3408 7840 3460
rect 7892 3448 7898 3460
rect 9140 3448 9168 3479
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9587 3519 9645 3525
rect 9587 3516 9599 3519
rect 9456 3488 9599 3516
rect 9456 3476 9462 3488
rect 9587 3485 9599 3488
rect 9633 3485 9645 3519
rect 9587 3479 9645 3485
rect 10502 3476 10508 3528
rect 10560 3476 10566 3528
rect 10594 3476 10600 3528
rect 10652 3476 10658 3528
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3516 11207 3519
rect 11238 3516 11244 3528
rect 11195 3488 11244 3516
rect 11195 3485 11207 3488
rect 11149 3479 11207 3485
rect 10520 3448 10548 3476
rect 7892 3420 10548 3448
rect 10888 3448 10916 3479
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3516 11483 3519
rect 11471 3488 11928 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 11900 3448 11928 3488
rect 14458 3476 14464 3528
rect 14516 3476 14522 3528
rect 14568 3488 14964 3516
rect 12066 3448 12072 3460
rect 10888 3420 11468 3448
rect 11900 3420 12072 3448
rect 7892 3408 7898 3420
rect 11440 3392 11468 3420
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 12158 3408 12164 3460
rect 12216 3408 12222 3460
rect 14182 3448 14188 3460
rect 13386 3420 14188 3448
rect 14182 3408 14188 3420
rect 14240 3408 14246 3460
rect 14274 3408 14280 3460
rect 14332 3408 14338 3460
rect 5316 3352 6316 3380
rect 5316 3340 5322 3352
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 9585 3383 9643 3389
rect 9585 3380 9597 3383
rect 9180 3352 9597 3380
rect 9180 3340 9186 3352
rect 9585 3349 9597 3352
rect 9631 3380 9643 3383
rect 10502 3380 10508 3392
rect 9631 3352 10508 3380
rect 9631 3349 9643 3352
rect 9585 3343 9643 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 11422 3340 11428 3392
rect 11480 3340 11486 3392
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 14568 3389 14596 3488
rect 14829 3451 14887 3457
rect 14829 3417 14841 3451
rect 14875 3417 14887 3451
rect 14936 3448 14964 3488
rect 15378 3476 15384 3528
rect 15436 3476 15442 3528
rect 16942 3476 16948 3528
rect 17000 3516 17006 3528
rect 17681 3519 17739 3525
rect 17681 3516 17693 3519
rect 17000 3488 17693 3516
rect 17000 3476 17006 3488
rect 17681 3485 17693 3488
rect 17727 3485 17739 3519
rect 17880 3516 17908 3624
rect 17972 3593 18000 3692
rect 17957 3587 18015 3593
rect 17957 3553 17969 3587
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17880 3488 18153 3516
rect 17681 3479 17739 3485
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 15562 3448 15568 3460
rect 14936 3420 15568 3448
rect 14829 3411 14887 3417
rect 14553 3383 14611 3389
rect 14553 3380 14565 3383
rect 12032 3352 14565 3380
rect 12032 3340 12038 3352
rect 14553 3349 14565 3352
rect 14599 3349 14611 3383
rect 14553 3343 14611 3349
rect 14642 3340 14648 3392
rect 14700 3340 14706 3392
rect 14844 3380 14872 3411
rect 15562 3408 15568 3420
rect 15620 3408 15626 3460
rect 15657 3451 15715 3457
rect 15657 3417 15669 3451
rect 15703 3448 15715 3451
rect 15746 3448 15752 3460
rect 15703 3420 15752 3448
rect 15703 3417 15715 3420
rect 15657 3411 15715 3417
rect 15746 3408 15752 3420
rect 15804 3408 15810 3460
rect 19518 3448 19524 3460
rect 16882 3420 19524 3448
rect 19518 3408 19524 3420
rect 19576 3408 19582 3460
rect 17218 3380 17224 3392
rect 14844 3352 17224 3380
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 1104 3290 18860 3312
rect 1104 3238 5502 3290
rect 5554 3238 5566 3290
rect 5618 3238 5630 3290
rect 5682 3238 5694 3290
rect 5746 3238 5758 3290
rect 5810 3238 5822 3290
rect 5874 3238 5886 3290
rect 5938 3238 5950 3290
rect 6002 3238 6014 3290
rect 6066 3238 6078 3290
rect 6130 3238 6142 3290
rect 6194 3238 6206 3290
rect 6258 3238 6270 3290
rect 6322 3238 6334 3290
rect 6386 3238 6398 3290
rect 6450 3238 6462 3290
rect 6514 3238 6526 3290
rect 6578 3238 6590 3290
rect 6642 3238 6654 3290
rect 6706 3238 13502 3290
rect 13554 3238 13566 3290
rect 13618 3238 13630 3290
rect 13682 3238 13694 3290
rect 13746 3238 13758 3290
rect 13810 3238 13822 3290
rect 13874 3238 13886 3290
rect 13938 3238 13950 3290
rect 14002 3238 14014 3290
rect 14066 3238 14078 3290
rect 14130 3238 14142 3290
rect 14194 3238 14206 3290
rect 14258 3238 14270 3290
rect 14322 3238 14334 3290
rect 14386 3238 14398 3290
rect 14450 3238 14462 3290
rect 14514 3238 14526 3290
rect 14578 3238 14590 3290
rect 14642 3238 14654 3290
rect 14706 3238 18860 3290
rect 1104 3216 18860 3238
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 2740 3148 4077 3176
rect 2740 3136 2746 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 4065 3139 4123 3145
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 6822 3176 6828 3188
rect 5592 3148 6828 3176
rect 5592 3136 5598 3148
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7009 3179 7067 3185
rect 7009 3145 7021 3179
rect 7055 3176 7067 3179
rect 7650 3176 7656 3188
rect 7055 3148 7656 3176
rect 7055 3145 7067 3148
rect 7009 3139 7067 3145
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 8018 3136 8024 3188
rect 8076 3136 8082 3188
rect 8386 3136 8392 3188
rect 8444 3136 8450 3188
rect 8481 3179 8539 3185
rect 8481 3145 8493 3179
rect 8527 3176 8539 3179
rect 9214 3176 9220 3188
rect 8527 3148 9220 3176
rect 8527 3145 8539 3148
rect 8481 3139 8539 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9401 3179 9459 3185
rect 9401 3145 9413 3179
rect 9447 3176 9459 3179
rect 9447 3148 10916 3176
rect 9447 3145 9459 3148
rect 9401 3139 9459 3145
rect 2406 3068 2412 3120
rect 2464 3108 2470 3120
rect 3973 3111 4031 3117
rect 3973 3108 3985 3111
rect 2464 3080 3985 3108
rect 2464 3068 2470 3080
rect 3973 3077 3985 3080
rect 4019 3077 4031 3111
rect 3973 3071 4031 3077
rect 5350 3068 5356 3120
rect 5408 3108 5414 3120
rect 5721 3111 5779 3117
rect 5721 3108 5733 3111
rect 5408 3080 5733 3108
rect 5408 3068 5414 3080
rect 5721 3077 5733 3080
rect 5767 3077 5779 3111
rect 5721 3071 5779 3077
rect 7285 3111 7343 3117
rect 7285 3077 7297 3111
rect 7331 3108 7343 3111
rect 8662 3108 8668 3120
rect 7331 3080 8668 3108
rect 7331 3077 7343 3080
rect 7285 3071 7343 3077
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 9582 3068 9588 3120
rect 9640 3068 9646 3120
rect 10888 3108 10916 3148
rect 12158 3136 12164 3188
rect 12216 3176 12222 3188
rect 13265 3179 13323 3185
rect 13265 3176 13277 3179
rect 12216 3148 13277 3176
rect 12216 3136 12222 3148
rect 13265 3145 13277 3148
rect 13311 3145 13323 3179
rect 13265 3139 13323 3145
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 13725 3179 13783 3185
rect 13725 3176 13737 3179
rect 13412 3148 13737 3176
rect 13412 3136 13418 3148
rect 13725 3145 13737 3148
rect 13771 3145 13783 3179
rect 15378 3176 15384 3188
rect 13725 3139 13783 3145
rect 14476 3148 15384 3176
rect 10888 3080 14412 3108
rect 1578 3000 1584 3052
rect 1636 3000 1642 3052
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 1688 3012 3341 3040
rect 1118 2932 1124 2984
rect 1176 2972 1182 2984
rect 1688 2972 1716 3012
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 5166 3000 5172 3052
rect 5224 3000 5230 3052
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3040 6791 3043
rect 7098 3040 7104 3052
rect 6779 3012 7104 3040
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 7834 3000 7840 3052
rect 7892 3000 7898 3052
rect 8570 3000 8576 3052
rect 8628 3000 8634 3052
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 9364 3012 10057 3040
rect 9364 3000 9370 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 10778 3000 10784 3052
rect 10836 3000 10842 3052
rect 11057 3043 11115 3049
rect 11057 3009 11069 3043
rect 11103 3040 11115 3043
rect 11103 3012 12020 3040
rect 11103 3009 11115 3012
rect 11057 3003 11115 3009
rect 1176 2944 1716 2972
rect 2317 2975 2375 2981
rect 1176 2932 1182 2944
rect 2317 2941 2329 2975
rect 2363 2941 2375 2975
rect 2317 2935 2375 2941
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2904 1823 2907
rect 2332 2904 2360 2935
rect 2866 2932 2872 2984
rect 2924 2932 2930 2984
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 8938 2972 8944 2984
rect 6696 2944 8944 2972
rect 6696 2932 6702 2944
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 11882 2972 11888 2984
rect 9232 2944 11888 2972
rect 1811 2876 2360 2904
rect 1811 2873 1823 2876
rect 1765 2867 1823 2873
rect 4614 2864 4620 2916
rect 4672 2904 4678 2916
rect 6822 2904 6828 2916
rect 4672 2876 6828 2904
rect 4672 2864 4678 2876
rect 6822 2864 6828 2876
rect 6880 2864 6886 2916
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 9232 2913 9260 2944
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 9217 2907 9275 2913
rect 9217 2904 9229 2907
rect 9088 2876 9229 2904
rect 9088 2864 9094 2876
rect 9217 2873 9229 2876
rect 9263 2873 9275 2907
rect 9217 2867 9275 2873
rect 10502 2864 10508 2916
rect 10560 2904 10566 2916
rect 10778 2904 10784 2916
rect 10560 2876 10784 2904
rect 10560 2864 10566 2876
rect 10778 2864 10784 2876
rect 10836 2864 10842 2916
rect 10870 2864 10876 2916
rect 10928 2904 10934 2916
rect 11238 2904 11244 2916
rect 10928 2876 11244 2904
rect 10928 2864 10934 2876
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 11992 2904 12020 3012
rect 12066 3000 12072 3052
rect 12124 3040 12130 3052
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 12124 3012 12173 3040
rect 12124 3000 12130 3012
rect 12161 3009 12173 3012
rect 12207 3040 12219 3043
rect 13262 3040 13268 3052
rect 12207 3012 13268 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 13906 3040 13912 3052
rect 13679 3012 13912 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 12253 2975 12311 2981
rect 12253 2941 12265 2975
rect 12299 2972 12311 2975
rect 12342 2972 12348 2984
rect 12299 2944 12348 2972
rect 12299 2941 12311 2944
rect 12253 2935 12311 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12710 2932 12716 2984
rect 12768 2932 12774 2984
rect 13078 2932 13084 2984
rect 13136 2972 13142 2984
rect 13817 2975 13875 2981
rect 13817 2972 13829 2975
rect 13136 2944 13829 2972
rect 13136 2932 13142 2944
rect 13817 2941 13829 2944
rect 13863 2941 13875 2975
rect 14384 2972 14412 3080
rect 14476 3049 14504 3148
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 16850 3176 16856 3188
rect 15620 3148 16856 3176
rect 15620 3136 15626 3148
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17034 3136 17040 3188
rect 17092 3176 17098 3188
rect 19610 3176 19616 3188
rect 17092 3148 19616 3176
rect 17092 3136 17098 3148
rect 19610 3136 19616 3148
rect 19668 3136 19674 3188
rect 14734 3068 14740 3120
rect 14792 3068 14798 3120
rect 16390 3108 16396 3120
rect 15962 3080 16396 3108
rect 16390 3068 16396 3080
rect 16448 3068 16454 3120
rect 18233 3111 18291 3117
rect 18233 3108 18245 3111
rect 17328 3080 18245 3108
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 16022 3000 16028 3052
rect 16080 3040 16086 3052
rect 16080 3012 17172 3040
rect 16080 3000 16086 3012
rect 14384 2944 16988 2972
rect 13817 2935 13875 2941
rect 12894 2904 12900 2916
rect 11992 2876 12900 2904
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 16960 2913 16988 2944
rect 17034 2932 17040 2984
rect 17092 2932 17098 2984
rect 17144 2972 17172 3012
rect 17218 3000 17224 3052
rect 17276 3040 17282 3052
rect 17328 3049 17356 3080
rect 18233 3077 18245 3080
rect 18279 3077 18291 3111
rect 18233 3071 18291 3077
rect 17313 3043 17371 3049
rect 17313 3040 17325 3043
rect 17276 3012 17325 3040
rect 17276 3000 17282 3012
rect 17313 3009 17325 3012
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 19886 3040 19892 3052
rect 18095 3012 19892 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 17865 2975 17923 2981
rect 17865 2972 17877 2975
rect 17144 2944 17877 2972
rect 17865 2941 17877 2944
rect 17911 2941 17923 2975
rect 17865 2935 17923 2941
rect 16945 2907 17003 2913
rect 16945 2873 16957 2907
rect 16991 2904 17003 2907
rect 17126 2904 17132 2916
rect 16991 2876 17132 2904
rect 16991 2873 17003 2876
rect 16945 2867 17003 2873
rect 17126 2864 17132 2876
rect 17184 2864 17190 2916
rect 3421 2839 3479 2845
rect 3421 2805 3433 2839
rect 3467 2836 3479 2839
rect 9122 2836 9128 2848
rect 3467 2808 9128 2836
rect 3467 2805 3479 2808
rect 3421 2799 3479 2805
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 10686 2836 10692 2848
rect 9447 2808 10692 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 16209 2839 16267 2845
rect 16209 2836 16221 2839
rect 15252 2808 16221 2836
rect 15252 2796 15258 2808
rect 16209 2805 16221 2808
rect 16255 2836 16267 2839
rect 18064 2836 18092 3003
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 16255 2808 18092 2836
rect 16255 2805 16267 2808
rect 16209 2799 16267 2805
rect 1104 2746 18860 2768
rect 1104 2694 1502 2746
rect 1554 2694 1566 2746
rect 1618 2694 1630 2746
rect 1682 2694 1694 2746
rect 1746 2694 1758 2746
rect 1810 2694 1822 2746
rect 1874 2694 1886 2746
rect 1938 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 2270 2746
rect 2322 2694 2334 2746
rect 2386 2694 2398 2746
rect 2450 2694 2462 2746
rect 2514 2694 2526 2746
rect 2578 2694 2590 2746
rect 2642 2694 2654 2746
rect 2706 2694 9502 2746
rect 9554 2694 9566 2746
rect 9618 2694 9630 2746
rect 9682 2694 9694 2746
rect 9746 2694 9758 2746
rect 9810 2694 9822 2746
rect 9874 2694 9886 2746
rect 9938 2694 9950 2746
rect 10002 2694 10014 2746
rect 10066 2694 10078 2746
rect 10130 2694 10142 2746
rect 10194 2694 10206 2746
rect 10258 2694 10270 2746
rect 10322 2694 10334 2746
rect 10386 2694 10398 2746
rect 10450 2694 10462 2746
rect 10514 2694 10526 2746
rect 10578 2694 10590 2746
rect 10642 2694 10654 2746
rect 10706 2694 17502 2746
rect 17554 2694 17566 2746
rect 17618 2694 17630 2746
rect 17682 2694 17694 2746
rect 17746 2694 17758 2746
rect 17810 2694 17822 2746
rect 17874 2694 17886 2746
rect 17938 2694 17950 2746
rect 18002 2694 18014 2746
rect 18066 2694 18078 2746
rect 18130 2694 18142 2746
rect 18194 2694 18206 2746
rect 18258 2694 18270 2746
rect 18322 2694 18334 2746
rect 18386 2694 18398 2746
rect 18450 2694 18462 2746
rect 18514 2694 18526 2746
rect 18578 2694 18590 2746
rect 18642 2694 18654 2746
rect 18706 2694 18860 2746
rect 1104 2672 18860 2694
rect 1394 2592 1400 2644
rect 1452 2632 1458 2644
rect 1581 2635 1639 2641
rect 1581 2632 1593 2635
rect 1452 2604 1593 2632
rect 1452 2592 1458 2604
rect 1581 2601 1593 2604
rect 1627 2601 1639 2635
rect 1581 2595 1639 2601
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 4154 2632 4160 2644
rect 3099 2604 4160 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 6733 2635 6791 2641
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 6822 2632 6828 2644
rect 6779 2604 6828 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 6914 2592 6920 2644
rect 6972 2592 6978 2644
rect 7745 2635 7803 2641
rect 7745 2601 7757 2635
rect 7791 2632 7803 2635
rect 7834 2632 7840 2644
rect 7791 2604 7840 2632
rect 7791 2601 7803 2604
rect 7745 2595 7803 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 8628 2604 10885 2632
rect 8628 2592 8634 2604
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 10873 2595 10931 2601
rect 12894 2592 12900 2644
rect 12952 2592 12958 2644
rect 13906 2592 13912 2644
rect 13964 2632 13970 2644
rect 14553 2635 14611 2641
rect 14553 2632 14565 2635
rect 13964 2604 14565 2632
rect 13964 2592 13970 2604
rect 14553 2601 14565 2604
rect 14599 2632 14611 2635
rect 15010 2632 15016 2644
rect 14599 2604 15016 2632
rect 14599 2601 14611 2604
rect 14553 2595 14611 2601
rect 15010 2592 15016 2604
rect 15068 2592 15074 2644
rect 16043 2635 16101 2641
rect 16043 2601 16055 2635
rect 16089 2632 16101 2635
rect 19242 2632 19248 2644
rect 16089 2604 19248 2632
rect 16089 2601 16101 2604
rect 16043 2595 16101 2601
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 934 2524 940 2576
rect 992 2564 998 2576
rect 5074 2564 5080 2576
rect 992 2536 5080 2564
rect 992 2524 998 2536
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 9416 2536 15056 2564
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2496 1639 2499
rect 4157 2499 4215 2505
rect 4157 2496 4169 2499
rect 1627 2468 4169 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 4157 2465 4169 2468
rect 4203 2465 4215 2499
rect 4157 2459 4215 2465
rect 4430 2456 4436 2508
rect 4488 2496 4494 2508
rect 8205 2499 8263 2505
rect 4488 2468 6592 2496
rect 4488 2456 4494 2468
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 3142 2428 3148 2440
rect 1995 2400 3148 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 3326 2388 3332 2440
rect 3384 2388 3390 2440
rect 5350 2388 5356 2440
rect 5408 2388 5414 2440
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 6564 2369 6592 2468
rect 8205 2465 8217 2499
rect 8251 2496 8263 2499
rect 8386 2496 8392 2508
rect 8251 2468 8392 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 9030 2456 9036 2508
rect 9088 2496 9094 2508
rect 9088 2468 9260 2496
rect 9088 2456 9094 2468
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 4709 2363 4767 2369
rect 4709 2360 4721 2363
rect 4212 2332 4721 2360
rect 4212 2320 4218 2332
rect 4709 2329 4721 2332
rect 4755 2329 4767 2363
rect 4709 2323 4767 2329
rect 6549 2363 6607 2369
rect 6549 2329 6561 2363
rect 6595 2329 6607 2363
rect 6549 2323 6607 2329
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 5224 2264 6745 2292
rect 5224 2252 5230 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 7558 2252 7564 2304
rect 7616 2252 7622 2304
rect 7760 2292 7788 2391
rect 8128 2360 8156 2391
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 9232 2428 9260 2468
rect 9306 2456 9312 2508
rect 9364 2456 9370 2508
rect 9416 2505 9444 2536
rect 15028 2508 15056 2536
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 9766 2456 9772 2508
rect 9824 2496 9830 2508
rect 11054 2496 11060 2508
rect 9824 2468 10364 2496
rect 9824 2456 9830 2468
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 9232 2400 9505 2428
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9674 2428 9680 2440
rect 9631 2400 9680 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10336 2437 10364 2468
rect 10428 2468 11060 2496
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 9214 2360 9220 2372
rect 8128 2332 9220 2360
rect 9214 2320 9220 2332
rect 9272 2360 9278 2372
rect 9769 2363 9827 2369
rect 9769 2360 9781 2363
rect 9272 2332 9781 2360
rect 9272 2320 9278 2332
rect 9769 2329 9781 2332
rect 9815 2329 9827 2363
rect 9769 2323 9827 2329
rect 10428 2292 10456 2468
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11848 2468 11897 2496
rect 11848 2456 11854 2468
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 13078 2456 13084 2508
rect 13136 2456 13142 2508
rect 15010 2456 15016 2508
rect 15068 2456 15074 2508
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 16301 2499 16359 2505
rect 16301 2496 16313 2499
rect 15436 2468 16313 2496
rect 15436 2456 15442 2468
rect 16301 2465 16313 2468
rect 16347 2465 16359 2499
rect 16301 2459 16359 2465
rect 16666 2456 16672 2508
rect 16724 2496 16730 2508
rect 16724 2468 17080 2496
rect 16724 2456 16730 2468
rect 10741 2431 10799 2437
rect 10741 2397 10753 2431
rect 10787 2428 10799 2431
rect 10870 2428 10876 2440
rect 10787 2400 10876 2428
rect 10787 2397 10799 2400
rect 10741 2391 10799 2397
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11572 2400 11989 2428
rect 11572 2388 11578 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12308 2400 12357 2428
rect 12308 2388 12314 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 10505 2363 10563 2369
rect 10505 2329 10517 2363
rect 10551 2329 10563 2363
rect 10505 2323 10563 2329
rect 7760 2264 10456 2292
rect 10520 2292 10548 2323
rect 10594 2320 10600 2372
rect 10652 2360 10658 2372
rect 11238 2360 11244 2372
rect 10652 2332 11244 2360
rect 10652 2320 10658 2332
rect 11238 2320 11244 2332
rect 11296 2320 11302 2372
rect 10778 2292 10784 2304
rect 10520 2264 10784 2292
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 12250 2252 12256 2304
rect 12308 2252 12314 2304
rect 12360 2292 12388 2391
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 12492 2400 13277 2428
rect 12492 2388 12498 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 13354 2388 13360 2440
rect 13412 2388 13418 2440
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 16850 2388 16856 2440
rect 16908 2388 16914 2440
rect 17052 2437 17080 2468
rect 17126 2456 17132 2508
rect 17184 2496 17190 2508
rect 17405 2499 17463 2505
rect 17405 2496 17417 2499
rect 17184 2468 17417 2496
rect 17184 2456 17190 2468
rect 17405 2465 17417 2468
rect 17451 2465 17463 2499
rect 17405 2459 17463 2465
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17862 2388 17868 2440
rect 17920 2388 17926 2440
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2428 18107 2431
rect 19702 2428 19708 2440
rect 18095 2400 19708 2428
rect 18095 2397 18107 2400
rect 18049 2391 18107 2397
rect 19702 2388 19708 2400
rect 19760 2388 19766 2440
rect 18233 2363 18291 2369
rect 18233 2360 18245 2363
rect 14476 2332 14688 2360
rect 14476 2292 14504 2332
rect 12360 2264 14504 2292
rect 14660 2292 14688 2332
rect 16132 2332 18245 2360
rect 16132 2292 16160 2332
rect 18233 2329 18245 2332
rect 18279 2329 18291 2363
rect 18233 2323 18291 2329
rect 14660 2264 16160 2292
rect 17034 2252 17040 2304
rect 17092 2292 17098 2304
rect 17310 2292 17316 2304
rect 17092 2264 17316 2292
rect 17092 2252 17098 2264
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 1104 2202 18860 2224
rect 1104 2150 5502 2202
rect 5554 2150 5566 2202
rect 5618 2150 5630 2202
rect 5682 2150 5694 2202
rect 5746 2150 5758 2202
rect 5810 2150 5822 2202
rect 5874 2150 5886 2202
rect 5938 2150 5950 2202
rect 6002 2150 6014 2202
rect 6066 2150 6078 2202
rect 6130 2150 6142 2202
rect 6194 2150 6206 2202
rect 6258 2150 6270 2202
rect 6322 2150 6334 2202
rect 6386 2150 6398 2202
rect 6450 2150 6462 2202
rect 6514 2150 6526 2202
rect 6578 2150 6590 2202
rect 6642 2150 6654 2202
rect 6706 2150 13502 2202
rect 13554 2150 13566 2202
rect 13618 2150 13630 2202
rect 13682 2150 13694 2202
rect 13746 2150 13758 2202
rect 13810 2150 13822 2202
rect 13874 2150 13886 2202
rect 13938 2150 13950 2202
rect 14002 2150 14014 2202
rect 14066 2150 14078 2202
rect 14130 2150 14142 2202
rect 14194 2150 14206 2202
rect 14258 2150 14270 2202
rect 14322 2150 14334 2202
rect 14386 2150 14398 2202
rect 14450 2150 14462 2202
rect 14514 2150 14526 2202
rect 14578 2150 14590 2202
rect 14642 2150 14654 2202
rect 14706 2150 18860 2202
rect 1104 2128 18860 2150
rect 3510 2048 3516 2100
rect 3568 2088 3574 2100
rect 3568 2060 6914 2088
rect 3568 2048 3574 2060
rect 6886 1952 6914 2060
rect 9674 2048 9680 2100
rect 9732 2088 9738 2100
rect 11146 2088 11152 2100
rect 9732 2060 11152 2088
rect 9732 2048 9738 2060
rect 11146 2048 11152 2060
rect 11204 2048 11210 2100
rect 12250 2048 12256 2100
rect 12308 2088 12314 2100
rect 14826 2088 14832 2100
rect 12308 2060 14832 2088
rect 12308 2048 12314 2060
rect 14826 2048 14832 2060
rect 14884 2048 14890 2100
rect 15010 2048 15016 2100
rect 15068 2088 15074 2100
rect 17034 2088 17040 2100
rect 15068 2060 17040 2088
rect 15068 2048 15074 2060
rect 17034 2048 17040 2060
rect 17092 2048 17098 2100
rect 7926 1980 7932 2032
rect 7984 2020 7990 2032
rect 15838 2020 15844 2032
rect 7984 1992 15844 2020
rect 7984 1980 7990 1992
rect 15838 1980 15844 1992
rect 15896 1980 15902 2032
rect 8110 1952 8116 1964
rect 6886 1924 8116 1952
rect 8110 1912 8116 1924
rect 8168 1952 8174 1964
rect 8168 1924 10916 1952
rect 8168 1912 8174 1924
rect 10888 1884 10916 1924
rect 17862 1884 17868 1896
rect 10888 1856 17868 1884
rect 17862 1844 17868 1856
rect 17920 1844 17926 1896
rect 3418 1776 3424 1828
rect 3476 1816 3482 1828
rect 10594 1816 10600 1828
rect 3476 1788 10600 1816
rect 3476 1776 3482 1788
rect 10594 1776 10600 1788
rect 10652 1776 10658 1828
rect 9122 1708 9128 1760
rect 9180 1748 9186 1760
rect 19334 1748 19340 1760
rect 9180 1720 19340 1748
rect 9180 1708 9186 1720
rect 19334 1708 19340 1720
rect 19392 1708 19398 1760
rect 7558 1640 7564 1692
rect 7616 1680 7622 1692
rect 18782 1680 18788 1692
rect 7616 1652 18788 1680
rect 7616 1640 7622 1652
rect 18782 1640 18788 1652
rect 18840 1640 18846 1692
rect 3418 1300 3424 1352
rect 3476 1340 3482 1352
rect 10962 1340 10968 1352
rect 3476 1312 10968 1340
rect 3476 1300 3482 1312
rect 10962 1300 10968 1312
rect 11020 1300 11026 1352
rect 4062 1232 4068 1284
rect 4120 1272 4126 1284
rect 15378 1272 15384 1284
rect 4120 1244 15384 1272
rect 4120 1232 4126 1244
rect 15378 1232 15384 1244
rect 15436 1232 15442 1284
rect 3326 1164 3332 1216
rect 3384 1204 3390 1216
rect 9582 1204 9588 1216
rect 3384 1176 9588 1204
rect 3384 1164 3390 1176
rect 9582 1164 9588 1176
rect 9640 1164 9646 1216
rect 3510 1028 3516 1080
rect 3568 1068 3574 1080
rect 8846 1068 8852 1080
rect 3568 1040 8852 1068
rect 3568 1028 3574 1040
rect 8846 1028 8852 1040
rect 8904 1028 8910 1080
rect 290 960 296 1012
rect 348 1000 354 1012
rect 5258 1000 5264 1012
rect 348 972 5264 1000
rect 348 960 354 972
rect 5258 960 5264 972
rect 5316 960 5322 1012
<< via1 >>
rect 1584 17484 1636 17536
rect 7932 17484 7984 17536
rect 5502 17382 5554 17434
rect 5566 17382 5618 17434
rect 5630 17382 5682 17434
rect 5694 17382 5746 17434
rect 5758 17382 5810 17434
rect 5822 17382 5874 17434
rect 5886 17382 5938 17434
rect 5950 17382 6002 17434
rect 6014 17382 6066 17434
rect 6078 17382 6130 17434
rect 6142 17382 6194 17434
rect 6206 17382 6258 17434
rect 6270 17382 6322 17434
rect 6334 17382 6386 17434
rect 6398 17382 6450 17434
rect 6462 17382 6514 17434
rect 6526 17382 6578 17434
rect 6590 17382 6642 17434
rect 6654 17382 6706 17434
rect 13502 17382 13554 17434
rect 13566 17382 13618 17434
rect 13630 17382 13682 17434
rect 13694 17382 13746 17434
rect 13758 17382 13810 17434
rect 13822 17382 13874 17434
rect 13886 17382 13938 17434
rect 13950 17382 14002 17434
rect 14014 17382 14066 17434
rect 14078 17382 14130 17434
rect 14142 17382 14194 17434
rect 14206 17382 14258 17434
rect 14270 17382 14322 17434
rect 14334 17382 14386 17434
rect 14398 17382 14450 17434
rect 14462 17382 14514 17434
rect 14526 17382 14578 17434
rect 14590 17382 14642 17434
rect 14654 17382 14706 17434
rect 2320 17280 2372 17332
rect 4436 17280 4488 17332
rect 572 17212 624 17264
rect 20 17144 72 17196
rect 3332 17187 3384 17196
rect 3332 17153 3341 17187
rect 3341 17153 3375 17187
rect 3375 17153 3384 17187
rect 3332 17144 3384 17153
rect 7564 17212 7616 17264
rect 4344 17187 4396 17196
rect 4344 17153 4353 17187
rect 4353 17153 4387 17187
rect 4387 17153 4396 17187
rect 4344 17144 4396 17153
rect 4896 17187 4948 17196
rect 4896 17153 4905 17187
rect 4905 17153 4939 17187
rect 4939 17153 4948 17187
rect 4896 17144 4948 17153
rect 756 17076 808 17128
rect 2044 17076 2096 17128
rect 9036 17144 9088 17196
rect 1216 17008 1268 17060
rect 1952 17008 2004 17060
rect 3240 17008 3292 17060
rect 3884 17008 3936 17060
rect 11152 17008 11204 17060
rect 1308 16940 1360 16992
rect 1768 16940 1820 16992
rect 4528 16940 4580 16992
rect 1502 16838 1554 16890
rect 1566 16838 1618 16890
rect 1630 16838 1682 16890
rect 1694 16838 1746 16890
rect 1758 16838 1810 16890
rect 1822 16838 1874 16890
rect 1886 16838 1938 16890
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 2270 16838 2322 16890
rect 2334 16838 2386 16890
rect 2398 16838 2450 16890
rect 2462 16838 2514 16890
rect 2526 16838 2578 16890
rect 2590 16838 2642 16890
rect 2654 16838 2706 16890
rect 9502 16838 9554 16890
rect 9566 16838 9618 16890
rect 9630 16838 9682 16890
rect 9694 16838 9746 16890
rect 9758 16838 9810 16890
rect 9822 16838 9874 16890
rect 9886 16838 9938 16890
rect 9950 16838 10002 16890
rect 10014 16838 10066 16890
rect 10078 16838 10130 16890
rect 10142 16838 10194 16890
rect 10206 16838 10258 16890
rect 10270 16838 10322 16890
rect 10334 16838 10386 16890
rect 10398 16838 10450 16890
rect 10462 16838 10514 16890
rect 10526 16838 10578 16890
rect 10590 16838 10642 16890
rect 10654 16838 10706 16890
rect 17502 16838 17554 16890
rect 17566 16838 17618 16890
rect 17630 16838 17682 16890
rect 17694 16838 17746 16890
rect 17758 16838 17810 16890
rect 17822 16838 17874 16890
rect 17886 16838 17938 16890
rect 17950 16838 18002 16890
rect 18014 16838 18066 16890
rect 18078 16838 18130 16890
rect 18142 16838 18194 16890
rect 18206 16838 18258 16890
rect 18270 16838 18322 16890
rect 18334 16838 18386 16890
rect 18398 16838 18450 16890
rect 18462 16838 18514 16890
rect 18526 16838 18578 16890
rect 18590 16838 18642 16890
rect 18654 16838 18706 16890
rect 8484 16668 8536 16720
rect 940 16532 992 16584
rect 2780 16532 2832 16584
rect 4804 16532 4856 16584
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 5448 16575 5500 16584
rect 5448 16541 5457 16575
rect 5457 16541 5491 16575
rect 5491 16541 5500 16575
rect 5448 16532 5500 16541
rect 1952 16507 2004 16516
rect 1952 16473 1961 16507
rect 1961 16473 1995 16507
rect 1995 16473 2004 16507
rect 1952 16464 2004 16473
rect 2504 16439 2556 16448
rect 2504 16405 2513 16439
rect 2513 16405 2547 16439
rect 2547 16405 2556 16439
rect 2504 16396 2556 16405
rect 3608 16464 3660 16516
rect 3976 16507 4028 16516
rect 3976 16473 3985 16507
rect 3985 16473 4019 16507
rect 4019 16473 4028 16507
rect 3976 16464 4028 16473
rect 4344 16507 4396 16516
rect 4344 16473 4353 16507
rect 4353 16473 4387 16507
rect 4387 16473 4396 16507
rect 4344 16464 4396 16473
rect 4988 16464 5040 16516
rect 6736 16532 6788 16584
rect 7380 16464 7432 16516
rect 2964 16396 3016 16448
rect 12256 16396 12308 16448
rect 5502 16294 5554 16346
rect 5566 16294 5618 16346
rect 5630 16294 5682 16346
rect 5694 16294 5746 16346
rect 5758 16294 5810 16346
rect 5822 16294 5874 16346
rect 5886 16294 5938 16346
rect 5950 16294 6002 16346
rect 6014 16294 6066 16346
rect 6078 16294 6130 16346
rect 6142 16294 6194 16346
rect 6206 16294 6258 16346
rect 6270 16294 6322 16346
rect 6334 16294 6386 16346
rect 6398 16294 6450 16346
rect 6462 16294 6514 16346
rect 6526 16294 6578 16346
rect 6590 16294 6642 16346
rect 6654 16294 6706 16346
rect 13502 16294 13554 16346
rect 13566 16294 13618 16346
rect 13630 16294 13682 16346
rect 13694 16294 13746 16346
rect 13758 16294 13810 16346
rect 13822 16294 13874 16346
rect 13886 16294 13938 16346
rect 13950 16294 14002 16346
rect 14014 16294 14066 16346
rect 14078 16294 14130 16346
rect 14142 16294 14194 16346
rect 14206 16294 14258 16346
rect 14270 16294 14322 16346
rect 14334 16294 14386 16346
rect 14398 16294 14450 16346
rect 14462 16294 14514 16346
rect 14526 16294 14578 16346
rect 14590 16294 14642 16346
rect 14654 16294 14706 16346
rect 2504 16124 2556 16176
rect 388 16056 440 16108
rect 3056 16056 3108 16108
rect 3424 16099 3476 16108
rect 3424 16065 3433 16099
rect 3433 16065 3467 16099
rect 3467 16065 3476 16099
rect 3424 16056 3476 16065
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 3700 16099 3752 16108
rect 3700 16065 3709 16099
rect 3709 16065 3743 16099
rect 3743 16065 3752 16099
rect 4620 16167 4672 16176
rect 4620 16133 4629 16167
rect 4629 16133 4663 16167
rect 4663 16133 4672 16167
rect 4620 16124 4672 16133
rect 6276 16124 6328 16176
rect 9220 16124 9272 16176
rect 3700 16056 3752 16065
rect 6828 16056 6880 16108
rect 480 15988 532 16040
rect 5264 15988 5316 16040
rect 7472 16099 7524 16108
rect 7472 16065 7481 16099
rect 7481 16065 7515 16099
rect 7515 16065 7524 16099
rect 7472 16056 7524 16065
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 9128 15988 9180 16040
rect 1952 15920 2004 15972
rect 2688 15920 2740 15972
rect 3332 15920 3384 15972
rect 12348 15920 12400 15972
rect 3148 15852 3200 15904
rect 4528 15852 4580 15904
rect 4712 15852 4764 15904
rect 4988 15852 5040 15904
rect 6736 15852 6788 15904
rect 6920 15852 6972 15904
rect 1502 15750 1554 15802
rect 1566 15750 1618 15802
rect 1630 15750 1682 15802
rect 1694 15750 1746 15802
rect 1758 15750 1810 15802
rect 1822 15750 1874 15802
rect 1886 15750 1938 15802
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 2270 15750 2322 15802
rect 2334 15750 2386 15802
rect 2398 15750 2450 15802
rect 2462 15750 2514 15802
rect 2526 15750 2578 15802
rect 2590 15750 2642 15802
rect 2654 15750 2706 15802
rect 9502 15750 9554 15802
rect 9566 15750 9618 15802
rect 9630 15750 9682 15802
rect 9694 15750 9746 15802
rect 9758 15750 9810 15802
rect 9822 15750 9874 15802
rect 9886 15750 9938 15802
rect 9950 15750 10002 15802
rect 10014 15750 10066 15802
rect 10078 15750 10130 15802
rect 10142 15750 10194 15802
rect 10206 15750 10258 15802
rect 10270 15750 10322 15802
rect 10334 15750 10386 15802
rect 10398 15750 10450 15802
rect 10462 15750 10514 15802
rect 10526 15750 10578 15802
rect 10590 15750 10642 15802
rect 10654 15750 10706 15802
rect 17502 15750 17554 15802
rect 17566 15750 17618 15802
rect 17630 15750 17682 15802
rect 17694 15750 17746 15802
rect 17758 15750 17810 15802
rect 17822 15750 17874 15802
rect 17886 15750 17938 15802
rect 17950 15750 18002 15802
rect 18014 15750 18066 15802
rect 18078 15750 18130 15802
rect 18142 15750 18194 15802
rect 18206 15750 18258 15802
rect 18270 15750 18322 15802
rect 18334 15750 18386 15802
rect 18398 15750 18450 15802
rect 18462 15750 18514 15802
rect 18526 15750 18578 15802
rect 18590 15750 18642 15802
rect 18654 15750 18706 15802
rect 2596 15648 2648 15700
rect 2872 15648 2924 15700
rect 1584 15580 1636 15632
rect 3332 15648 3384 15700
rect 5356 15691 5408 15700
rect 5356 15657 5365 15691
rect 5365 15657 5399 15691
rect 5399 15657 5408 15691
rect 5356 15648 5408 15657
rect 6184 15691 6236 15700
rect 6184 15657 6193 15691
rect 6193 15657 6227 15691
rect 6227 15657 6236 15691
rect 6184 15648 6236 15657
rect 6276 15648 6328 15700
rect 8208 15648 8260 15700
rect 3792 15580 3844 15632
rect 296 15512 348 15564
rect 4896 15580 4948 15632
rect 8576 15580 8628 15632
rect 480 15444 532 15496
rect 664 15444 716 15496
rect 1952 15487 2004 15496
rect 1952 15453 1961 15487
rect 1961 15453 1995 15487
rect 1995 15453 2004 15487
rect 1952 15444 2004 15453
rect 2688 15487 2740 15496
rect 2688 15453 2697 15487
rect 2697 15453 2731 15487
rect 2731 15453 2740 15487
rect 2688 15444 2740 15453
rect 2964 15444 3016 15496
rect 7104 15512 7156 15564
rect 8392 15512 8444 15564
rect 204 15376 256 15428
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 4160 15444 4212 15496
rect 7564 15444 7616 15496
rect 19064 15512 19116 15564
rect 664 15308 716 15360
rect 1032 15308 1084 15360
rect 1860 15308 1912 15360
rect 3424 15376 3476 15428
rect 5172 15419 5224 15428
rect 5172 15385 5181 15419
rect 5181 15385 5215 15419
rect 5215 15385 5224 15419
rect 5172 15376 5224 15385
rect 6276 15419 6328 15428
rect 6276 15385 6285 15419
rect 6285 15385 6319 15419
rect 6319 15385 6328 15419
rect 6276 15376 6328 15385
rect 6736 15376 6788 15428
rect 7012 15376 7064 15428
rect 3332 15308 3384 15360
rect 3884 15308 3936 15360
rect 4252 15308 4304 15360
rect 4528 15308 4580 15360
rect 4988 15308 5040 15360
rect 7288 15419 7340 15428
rect 7288 15385 7297 15419
rect 7297 15385 7331 15419
rect 7331 15385 7340 15419
rect 7288 15376 7340 15385
rect 8116 15419 8168 15428
rect 8116 15385 8125 15419
rect 8125 15385 8159 15419
rect 8159 15385 8168 15419
rect 8116 15376 8168 15385
rect 8208 15376 8260 15428
rect 8576 15376 8628 15428
rect 8024 15308 8076 15360
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 12808 15308 12860 15360
rect 296 15240 348 15292
rect 756 15240 808 15292
rect 5502 15206 5554 15258
rect 5566 15206 5618 15258
rect 5630 15206 5682 15258
rect 5694 15206 5746 15258
rect 5758 15206 5810 15258
rect 5822 15206 5874 15258
rect 5886 15206 5938 15258
rect 5950 15206 6002 15258
rect 6014 15206 6066 15258
rect 6078 15206 6130 15258
rect 6142 15206 6194 15258
rect 6206 15206 6258 15258
rect 6270 15206 6322 15258
rect 6334 15206 6386 15258
rect 6398 15206 6450 15258
rect 6462 15206 6514 15258
rect 6526 15206 6578 15258
rect 6590 15206 6642 15258
rect 6654 15206 6706 15258
rect 13502 15206 13554 15258
rect 13566 15206 13618 15258
rect 13630 15206 13682 15258
rect 13694 15206 13746 15258
rect 13758 15206 13810 15258
rect 13822 15206 13874 15258
rect 13886 15206 13938 15258
rect 13950 15206 14002 15258
rect 14014 15206 14066 15258
rect 14078 15206 14130 15258
rect 14142 15206 14194 15258
rect 14206 15206 14258 15258
rect 14270 15206 14322 15258
rect 14334 15206 14386 15258
rect 14398 15206 14450 15258
rect 14462 15206 14514 15258
rect 14526 15206 14578 15258
rect 14590 15206 14642 15258
rect 14654 15206 14706 15258
rect 1860 15147 1912 15156
rect 1860 15113 1869 15147
rect 1869 15113 1903 15147
rect 1903 15113 1912 15147
rect 1860 15104 1912 15113
rect 3424 15104 3476 15156
rect 3700 15104 3752 15156
rect 1308 15036 1360 15088
rect 2872 15036 2924 15088
rect 4068 15036 4120 15088
rect 4344 15036 4396 15088
rect 756 14900 808 14952
rect 1584 14900 1636 14952
rect 2964 14900 3016 14952
rect 1308 14832 1360 14884
rect 1952 14832 2004 14884
rect 1032 14764 1084 14816
rect 4252 14968 4304 15020
rect 4528 15011 4580 15020
rect 4528 14977 4537 15011
rect 4537 14977 4571 15011
rect 4571 14977 4580 15011
rect 4528 14968 4580 14977
rect 4068 14900 4120 14952
rect 5080 14968 5132 15020
rect 5172 14968 5224 15020
rect 6552 15079 6604 15088
rect 6552 15045 6561 15079
rect 6561 15045 6595 15079
rect 6595 15045 6604 15079
rect 6552 15036 6604 15045
rect 7288 15036 7340 15088
rect 8208 15036 8260 15088
rect 8300 15036 8352 15088
rect 7656 14968 7708 15020
rect 4804 14900 4856 14952
rect 6000 14900 6052 14952
rect 8024 14968 8076 15020
rect 14740 15036 14792 15088
rect 7840 14900 7892 14952
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 8852 14900 8904 14952
rect 9128 14900 9180 14952
rect 4252 14832 4304 14884
rect 8760 14832 8812 14884
rect 9404 14875 9456 14884
rect 9404 14841 9413 14875
rect 9413 14841 9447 14875
rect 9447 14841 9456 14875
rect 9404 14832 9456 14841
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 4896 14764 4948 14773
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 6644 14764 6696 14816
rect 7472 14764 7524 14816
rect 8300 14764 8352 14816
rect 8944 14764 8996 14816
rect 1502 14662 1554 14714
rect 1566 14662 1618 14714
rect 1630 14662 1682 14714
rect 1694 14662 1746 14714
rect 1758 14662 1810 14714
rect 1822 14662 1874 14714
rect 1886 14662 1938 14714
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 2270 14662 2322 14714
rect 2334 14662 2386 14714
rect 2398 14662 2450 14714
rect 2462 14662 2514 14714
rect 2526 14662 2578 14714
rect 2590 14662 2642 14714
rect 2654 14662 2706 14714
rect 9502 14662 9554 14714
rect 9566 14662 9618 14714
rect 9630 14662 9682 14714
rect 9694 14662 9746 14714
rect 9758 14662 9810 14714
rect 9822 14662 9874 14714
rect 9886 14662 9938 14714
rect 9950 14662 10002 14714
rect 10014 14662 10066 14714
rect 10078 14662 10130 14714
rect 10142 14662 10194 14714
rect 10206 14662 10258 14714
rect 10270 14662 10322 14714
rect 10334 14662 10386 14714
rect 10398 14662 10450 14714
rect 10462 14662 10514 14714
rect 10526 14662 10578 14714
rect 10590 14662 10642 14714
rect 10654 14662 10706 14714
rect 17502 14662 17554 14714
rect 17566 14662 17618 14714
rect 17630 14662 17682 14714
rect 17694 14662 17746 14714
rect 17758 14662 17810 14714
rect 17822 14662 17874 14714
rect 17886 14662 17938 14714
rect 17950 14662 18002 14714
rect 18014 14662 18066 14714
rect 18078 14662 18130 14714
rect 18142 14662 18194 14714
rect 18206 14662 18258 14714
rect 18270 14662 18322 14714
rect 18334 14662 18386 14714
rect 18398 14662 18450 14714
rect 18462 14662 18514 14714
rect 18526 14662 18578 14714
rect 18590 14662 18642 14714
rect 18654 14662 18706 14714
rect 2136 14560 2188 14612
rect 4344 14603 4396 14612
rect 4344 14569 4353 14603
rect 4353 14569 4387 14603
rect 4387 14569 4396 14603
rect 4344 14560 4396 14569
rect 4528 14560 4580 14612
rect 4160 14492 4212 14544
rect 4804 14492 4856 14544
rect 5080 14560 5132 14612
rect 8024 14560 8076 14612
rect 4988 14492 5040 14544
rect 5816 14492 5868 14544
rect 8668 14492 8720 14544
rect 1216 14356 1268 14408
rect 2228 14356 2280 14408
rect 2964 14356 3016 14408
rect 756 14288 808 14340
rect 3700 14356 3752 14408
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 5448 14424 5500 14476
rect 5080 14356 5132 14408
rect 5724 14399 5776 14408
rect 5724 14365 5733 14399
rect 5733 14365 5767 14399
rect 5767 14365 5776 14399
rect 5724 14356 5776 14365
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 7472 14424 7524 14476
rect 7656 14424 7708 14476
rect 6460 14399 6512 14408
rect 6460 14365 6469 14399
rect 6469 14365 6503 14399
rect 6503 14365 6512 14399
rect 6460 14356 6512 14365
rect 7380 14356 7432 14408
rect 7840 14399 7892 14408
rect 7840 14365 7849 14399
rect 7849 14365 7883 14399
rect 7883 14365 7892 14399
rect 7840 14356 7892 14365
rect 8208 14356 8260 14408
rect 8760 14356 8812 14408
rect 9220 14399 9272 14408
rect 9220 14365 9229 14399
rect 9229 14365 9263 14399
rect 9263 14365 9272 14399
rect 9220 14356 9272 14365
rect 2044 14220 2096 14272
rect 2688 14220 2740 14272
rect 3424 14220 3476 14272
rect 4160 14220 4212 14272
rect 6000 14288 6052 14340
rect 7288 14288 7340 14340
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 13176 14424 13228 14476
rect 11796 14356 11848 14408
rect 15016 14424 15068 14476
rect 12440 14288 12492 14340
rect 15292 14356 15344 14408
rect 13544 14288 13596 14340
rect 19800 14288 19852 14340
rect 5264 14220 5316 14272
rect 6828 14220 6880 14272
rect 8024 14220 8076 14272
rect 8760 14220 8812 14272
rect 9404 14220 9456 14272
rect 10968 14220 11020 14272
rect 18972 14220 19024 14272
rect 5502 14118 5554 14170
rect 5566 14118 5618 14170
rect 5630 14118 5682 14170
rect 5694 14118 5746 14170
rect 5758 14118 5810 14170
rect 5822 14118 5874 14170
rect 5886 14118 5938 14170
rect 5950 14118 6002 14170
rect 6014 14118 6066 14170
rect 6078 14118 6130 14170
rect 6142 14118 6194 14170
rect 6206 14118 6258 14170
rect 6270 14118 6322 14170
rect 6334 14118 6386 14170
rect 6398 14118 6450 14170
rect 6462 14118 6514 14170
rect 6526 14118 6578 14170
rect 6590 14118 6642 14170
rect 6654 14118 6706 14170
rect 13502 14118 13554 14170
rect 13566 14118 13618 14170
rect 13630 14118 13682 14170
rect 13694 14118 13746 14170
rect 13758 14118 13810 14170
rect 13822 14118 13874 14170
rect 13886 14118 13938 14170
rect 13950 14118 14002 14170
rect 14014 14118 14066 14170
rect 14078 14118 14130 14170
rect 14142 14118 14194 14170
rect 14206 14118 14258 14170
rect 14270 14118 14322 14170
rect 14334 14118 14386 14170
rect 14398 14118 14450 14170
rect 14462 14118 14514 14170
rect 14526 14118 14578 14170
rect 14590 14118 14642 14170
rect 14654 14118 14706 14170
rect 1216 14016 1268 14068
rect 3056 14016 3108 14068
rect 572 13948 624 14000
rect 1308 13948 1360 14000
rect 2136 13991 2188 14000
rect 2136 13957 2145 13991
rect 2145 13957 2179 13991
rect 2179 13957 2188 13991
rect 2136 13948 2188 13957
rect 1124 13880 1176 13932
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 2872 13948 2924 14000
rect 3424 14016 3476 14068
rect 4528 14016 4580 14068
rect 4436 13948 4488 14000
rect 5908 13948 5960 14000
rect 572 13812 624 13864
rect 1308 13812 1360 13864
rect 1584 13812 1636 13864
rect 2688 13812 2740 13864
rect 3976 13880 4028 13932
rect 4160 13812 4212 13864
rect 1216 13676 1268 13728
rect 1860 13676 1912 13728
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 4804 13812 4856 13864
rect 6460 13880 6512 13932
rect 7288 13948 7340 14000
rect 9496 14016 9548 14068
rect 7472 13880 7524 13932
rect 7196 13812 7248 13864
rect 3056 13676 3108 13728
rect 4436 13676 4488 13728
rect 6644 13744 6696 13796
rect 8208 13948 8260 14000
rect 8576 13948 8628 14000
rect 9036 13948 9088 14000
rect 7840 13880 7892 13932
rect 5632 13719 5684 13728
rect 5632 13685 5641 13719
rect 5641 13685 5675 13719
rect 5675 13685 5684 13719
rect 5632 13676 5684 13685
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 7932 13676 7984 13728
rect 8300 13812 8352 13864
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 11980 13948 12032 14000
rect 15200 14016 15252 14068
rect 12992 13948 13044 14000
rect 13360 13948 13412 14000
rect 10324 13923 10376 13932
rect 10324 13889 10333 13923
rect 10333 13889 10367 13923
rect 10367 13889 10376 13923
rect 10324 13880 10376 13889
rect 11796 13880 11848 13932
rect 12900 13923 12952 13932
rect 12900 13889 12909 13923
rect 12909 13889 12943 13923
rect 12943 13889 12952 13923
rect 12900 13880 12952 13889
rect 12440 13812 12492 13864
rect 12716 13812 12768 13864
rect 13084 13812 13136 13864
rect 8852 13787 8904 13796
rect 8852 13753 8861 13787
rect 8861 13753 8895 13787
rect 8895 13753 8904 13787
rect 8852 13744 8904 13753
rect 14832 13948 14884 14000
rect 14924 13948 14976 14000
rect 19340 13948 19392 14000
rect 19892 13880 19944 13932
rect 19616 13812 19668 13864
rect 8576 13676 8628 13728
rect 11796 13719 11848 13728
rect 11796 13685 11805 13719
rect 11805 13685 11839 13719
rect 11839 13685 11848 13719
rect 11796 13676 11848 13685
rect 14924 13744 14976 13796
rect 16304 13676 16356 13728
rect 1502 13574 1554 13626
rect 1566 13574 1618 13626
rect 1630 13574 1682 13626
rect 1694 13574 1746 13626
rect 1758 13574 1810 13626
rect 1822 13574 1874 13626
rect 1886 13574 1938 13626
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 2270 13574 2322 13626
rect 2334 13574 2386 13626
rect 2398 13574 2450 13626
rect 2462 13574 2514 13626
rect 2526 13574 2578 13626
rect 2590 13574 2642 13626
rect 2654 13574 2706 13626
rect 9502 13574 9554 13626
rect 9566 13574 9618 13626
rect 9630 13574 9682 13626
rect 9694 13574 9746 13626
rect 9758 13574 9810 13626
rect 9822 13574 9874 13626
rect 9886 13574 9938 13626
rect 9950 13574 10002 13626
rect 10014 13574 10066 13626
rect 10078 13574 10130 13626
rect 10142 13574 10194 13626
rect 10206 13574 10258 13626
rect 10270 13574 10322 13626
rect 10334 13574 10386 13626
rect 10398 13574 10450 13626
rect 10462 13574 10514 13626
rect 10526 13574 10578 13626
rect 10590 13574 10642 13626
rect 10654 13574 10706 13626
rect 17502 13574 17554 13626
rect 17566 13574 17618 13626
rect 17630 13574 17682 13626
rect 17694 13574 17746 13626
rect 17758 13574 17810 13626
rect 17822 13574 17874 13626
rect 17886 13574 17938 13626
rect 17950 13574 18002 13626
rect 18014 13574 18066 13626
rect 18078 13574 18130 13626
rect 18142 13574 18194 13626
rect 18206 13574 18258 13626
rect 18270 13574 18322 13626
rect 18334 13574 18386 13626
rect 18398 13574 18450 13626
rect 18462 13574 18514 13626
rect 18526 13574 18578 13626
rect 18590 13574 18642 13626
rect 18654 13574 18706 13626
rect 664 13472 716 13524
rect 2228 13472 2280 13524
rect 2320 13472 2372 13524
rect 2872 13404 2924 13456
rect 1768 13311 1820 13320
rect 1768 13277 1777 13311
rect 1777 13277 1811 13311
rect 1811 13277 1820 13311
rect 1768 13268 1820 13277
rect 2412 13311 2464 13320
rect 2412 13277 2421 13311
rect 2421 13277 2455 13311
rect 2455 13277 2464 13311
rect 2412 13268 2464 13277
rect 2504 13268 2556 13320
rect 2872 13311 2924 13320
rect 2872 13277 2875 13311
rect 2875 13277 2924 13311
rect 2872 13268 2924 13277
rect 1952 13243 2004 13252
rect 1952 13209 1961 13243
rect 1961 13209 1995 13243
rect 1995 13209 2004 13243
rect 1952 13200 2004 13209
rect 2596 13243 2648 13252
rect 2596 13209 2605 13243
rect 2605 13209 2639 13243
rect 2639 13209 2648 13243
rect 2596 13200 2648 13209
rect 4160 13268 4212 13320
rect 4988 13472 5040 13524
rect 5172 13472 5224 13524
rect 5448 13472 5500 13524
rect 5540 13472 5592 13524
rect 6828 13472 6880 13524
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 4804 13404 4856 13456
rect 5356 13447 5408 13456
rect 5356 13413 5365 13447
rect 5365 13413 5399 13447
rect 5399 13413 5408 13447
rect 5356 13404 5408 13413
rect 5632 13404 5684 13456
rect 4804 13268 4856 13320
rect 8208 13447 8260 13456
rect 8208 13413 8217 13447
rect 8217 13413 8251 13447
rect 8251 13413 8260 13447
rect 8208 13404 8260 13413
rect 7840 13336 7892 13388
rect 8024 13336 8076 13388
rect 5080 13200 5132 13252
rect 6460 13268 6512 13320
rect 6644 13268 6696 13320
rect 8760 13404 8812 13456
rect 9220 13472 9272 13524
rect 12440 13472 12492 13524
rect 12624 13404 12676 13456
rect 11796 13336 11848 13388
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 7840 13200 7892 13252
rect 8760 13268 8812 13320
rect 9588 13311 9640 13320
rect 9588 13277 9597 13311
rect 9597 13277 9631 13311
rect 9631 13277 9640 13311
rect 9588 13268 9640 13277
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10416 13268 10468 13320
rect 11244 13268 11296 13320
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 480 13132 532 13184
rect 2872 13132 2924 13184
rect 4160 13132 4212 13184
rect 5448 13132 5500 13184
rect 7288 13132 7340 13184
rect 9956 13132 10008 13184
rect 10600 13132 10652 13184
rect 10784 13132 10836 13184
rect 11980 13175 12032 13184
rect 11980 13141 11989 13175
rect 11989 13141 12023 13175
rect 12023 13141 12032 13175
rect 11980 13132 12032 13141
rect 12624 13268 12676 13320
rect 15108 13336 15160 13388
rect 15292 13336 15344 13388
rect 16212 13336 16264 13388
rect 14740 13268 14792 13320
rect 14924 13268 14976 13320
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 17132 13268 17184 13320
rect 12716 13200 12768 13252
rect 15936 13200 15988 13252
rect 13360 13132 13412 13184
rect 15384 13132 15436 13184
rect 20 12996 72 13048
rect 480 12996 532 13048
rect 5502 13030 5554 13082
rect 5566 13030 5618 13082
rect 5630 13030 5682 13082
rect 5694 13030 5746 13082
rect 5758 13030 5810 13082
rect 5822 13030 5874 13082
rect 5886 13030 5938 13082
rect 5950 13030 6002 13082
rect 6014 13030 6066 13082
rect 6078 13030 6130 13082
rect 6142 13030 6194 13082
rect 6206 13030 6258 13082
rect 6270 13030 6322 13082
rect 6334 13030 6386 13082
rect 6398 13030 6450 13082
rect 6462 13030 6514 13082
rect 6526 13030 6578 13082
rect 6590 13030 6642 13082
rect 6654 13030 6706 13082
rect 13502 13030 13554 13082
rect 13566 13030 13618 13082
rect 13630 13030 13682 13082
rect 13694 13030 13746 13082
rect 13758 13030 13810 13082
rect 13822 13030 13874 13082
rect 13886 13030 13938 13082
rect 13950 13030 14002 13082
rect 14014 13030 14066 13082
rect 14078 13030 14130 13082
rect 14142 13030 14194 13082
rect 14206 13030 14258 13082
rect 14270 13030 14322 13082
rect 14334 13030 14386 13082
rect 14398 13030 14450 13082
rect 14462 13030 14514 13082
rect 14526 13030 14578 13082
rect 14590 13030 14642 13082
rect 14654 13030 14706 13082
rect 1308 12928 1360 12980
rect 2320 12971 2372 12980
rect 2320 12937 2329 12971
rect 2329 12937 2363 12971
rect 2363 12937 2372 12971
rect 2320 12928 2372 12937
rect 2688 12928 2740 12980
rect 2780 12928 2832 12980
rect 20 12860 72 12912
rect 112 12860 164 12912
rect 2412 12792 2464 12844
rect 3516 12860 3568 12912
rect 3700 12860 3752 12912
rect 4160 12928 4212 12980
rect 6184 12928 6236 12980
rect 4436 12860 4488 12912
rect 4988 12860 5040 12912
rect 2228 12767 2280 12776
rect 2228 12733 2254 12767
rect 2254 12733 2280 12767
rect 2228 12724 2280 12733
rect 2320 12724 2372 12776
rect 4252 12835 4304 12844
rect 2780 12724 2832 12776
rect 2872 12724 2924 12776
rect 3240 12724 3292 12776
rect 4252 12801 4260 12835
rect 4260 12801 4294 12835
rect 4294 12801 4304 12835
rect 4252 12792 4304 12801
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 2596 12656 2648 12708
rect 5448 12801 5500 12810
rect 5448 12767 5457 12801
rect 5457 12767 5491 12801
rect 5491 12767 5500 12801
rect 5448 12758 5500 12767
rect 5540 12835 5592 12844
rect 5540 12801 5549 12835
rect 5549 12801 5583 12835
rect 5583 12801 5592 12835
rect 5540 12792 5592 12801
rect 6736 12792 6788 12844
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 7196 12860 7248 12912
rect 7564 12860 7616 12912
rect 8300 12928 8352 12980
rect 6000 12724 6052 12776
rect 7380 12792 7432 12844
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 8852 12860 8904 12912
rect 9956 12860 10008 12912
rect 12624 12928 12676 12980
rect 13176 12928 13228 12980
rect 19248 12928 19300 12980
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 8208 12724 8260 12776
rect 8668 12792 8720 12844
rect 9496 12792 9548 12844
rect 9588 12792 9640 12844
rect 9036 12724 9088 12776
rect 1492 12588 1544 12640
rect 1860 12588 1912 12640
rect 2964 12588 3016 12640
rect 5172 12656 5224 12708
rect 5264 12656 5316 12708
rect 6552 12656 6604 12708
rect 6644 12656 6696 12708
rect 6920 12656 6972 12708
rect 5908 12588 5960 12640
rect 6368 12588 6420 12640
rect 9220 12656 9272 12708
rect 9772 12724 9824 12776
rect 10508 12724 10560 12776
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 11060 12835 11112 12844
rect 11060 12801 11069 12835
rect 11069 12801 11103 12835
rect 11103 12801 11112 12835
rect 11060 12792 11112 12801
rect 12072 12860 12124 12912
rect 11888 12792 11940 12844
rect 12900 12792 12952 12844
rect 11336 12724 11388 12776
rect 10416 12656 10468 12708
rect 12716 12767 12768 12776
rect 12716 12733 12725 12767
rect 12725 12733 12759 12767
rect 12759 12733 12768 12767
rect 12716 12724 12768 12733
rect 12992 12724 13044 12776
rect 15016 12792 15068 12844
rect 15476 12860 15528 12912
rect 15292 12792 15344 12844
rect 16396 12860 16448 12912
rect 16212 12835 16264 12844
rect 16212 12801 16221 12835
rect 16221 12801 16255 12835
rect 16255 12801 16264 12835
rect 16212 12792 16264 12801
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 16856 12724 16908 12776
rect 13452 12656 13504 12708
rect 7656 12588 7708 12640
rect 10600 12588 10652 12640
rect 10876 12588 10928 12640
rect 13176 12588 13228 12640
rect 14372 12631 14424 12640
rect 14372 12597 14381 12631
rect 14381 12597 14415 12631
rect 14415 12597 14424 12631
rect 14372 12588 14424 12597
rect 19524 12656 19576 12708
rect 19708 12588 19760 12640
rect 1502 12486 1554 12538
rect 1566 12486 1618 12538
rect 1630 12486 1682 12538
rect 1694 12486 1746 12538
rect 1758 12486 1810 12538
rect 1822 12486 1874 12538
rect 1886 12486 1938 12538
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 2270 12486 2322 12538
rect 2334 12486 2386 12538
rect 2398 12486 2450 12538
rect 2462 12486 2514 12538
rect 2526 12486 2578 12538
rect 2590 12486 2642 12538
rect 2654 12486 2706 12538
rect 9502 12486 9554 12538
rect 9566 12486 9618 12538
rect 9630 12486 9682 12538
rect 9694 12486 9746 12538
rect 9758 12486 9810 12538
rect 9822 12486 9874 12538
rect 9886 12486 9938 12538
rect 9950 12486 10002 12538
rect 10014 12486 10066 12538
rect 10078 12486 10130 12538
rect 10142 12486 10194 12538
rect 10206 12486 10258 12538
rect 10270 12486 10322 12538
rect 10334 12486 10386 12538
rect 10398 12486 10450 12538
rect 10462 12486 10514 12538
rect 10526 12486 10578 12538
rect 10590 12486 10642 12538
rect 10654 12486 10706 12538
rect 17502 12486 17554 12538
rect 17566 12486 17618 12538
rect 17630 12486 17682 12538
rect 17694 12486 17746 12538
rect 17758 12486 17810 12538
rect 17822 12486 17874 12538
rect 17886 12486 17938 12538
rect 17950 12486 18002 12538
rect 18014 12486 18066 12538
rect 18078 12486 18130 12538
rect 18142 12486 18194 12538
rect 18206 12486 18258 12538
rect 18270 12486 18322 12538
rect 18334 12486 18386 12538
rect 18398 12486 18450 12538
rect 18462 12486 18514 12538
rect 18526 12486 18578 12538
rect 18590 12486 18642 12538
rect 18654 12486 18706 12538
rect 1768 12384 1820 12436
rect 2872 12384 2924 12436
rect 2504 12316 2556 12368
rect 848 12248 900 12300
rect 2320 12291 2372 12300
rect 2320 12257 2329 12291
rect 2329 12257 2363 12291
rect 2363 12257 2372 12291
rect 2320 12248 2372 12257
rect 1768 12180 1820 12232
rect 4160 12384 4212 12436
rect 4896 12384 4948 12436
rect 5172 12384 5224 12436
rect 6276 12384 6328 12436
rect 8024 12384 8076 12436
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 5540 12316 5592 12368
rect 5632 12316 5684 12368
rect 7196 12316 7248 12368
rect 7932 12316 7984 12368
rect 4160 12248 4212 12300
rect 4252 12248 4304 12300
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 5080 12248 5132 12300
rect 5908 12248 5960 12300
rect 4896 12180 4948 12232
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 5816 12180 5868 12232
rect 7288 12248 7340 12300
rect 7012 12180 7064 12232
rect 5172 12112 5224 12164
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 3884 12044 3936 12096
rect 4252 12044 4304 12096
rect 5356 12112 5408 12164
rect 6276 12112 6328 12164
rect 6736 12044 6788 12096
rect 7288 12146 7340 12198
rect 8208 12316 8260 12368
rect 8668 12384 8720 12436
rect 9220 12384 9272 12436
rect 10416 12384 10468 12436
rect 10600 12427 10652 12436
rect 10600 12393 10609 12427
rect 10609 12393 10643 12427
rect 10643 12393 10652 12427
rect 10600 12384 10652 12393
rect 11336 12384 11388 12436
rect 11428 12384 11480 12436
rect 11704 12384 11756 12436
rect 10048 12316 10100 12368
rect 11244 12316 11296 12368
rect 13452 12384 13504 12436
rect 7748 12112 7800 12164
rect 9404 12248 9456 12300
rect 10232 12248 10284 12300
rect 10600 12248 10652 12300
rect 8944 12180 8996 12232
rect 8852 12112 8904 12164
rect 7288 12044 7340 12096
rect 7564 12044 7616 12096
rect 9680 12180 9732 12232
rect 10416 12180 10468 12232
rect 13360 12316 13412 12368
rect 16028 12316 16080 12368
rect 12532 12248 12584 12300
rect 14372 12248 14424 12300
rect 9864 12112 9916 12164
rect 10508 12112 10560 12164
rect 11888 12180 11940 12232
rect 11980 12180 12032 12232
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12716 12180 12768 12189
rect 12624 12112 12676 12164
rect 14832 12112 14884 12164
rect 15200 12223 15252 12232
rect 15200 12189 15209 12223
rect 15209 12189 15243 12223
rect 15243 12189 15252 12223
rect 15200 12180 15252 12189
rect 17224 12248 17276 12300
rect 16212 12180 16264 12232
rect 16396 12180 16448 12232
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 15660 12112 15712 12164
rect 16580 12112 16632 12164
rect 16764 12112 16816 12164
rect 17316 12112 17368 12164
rect 17868 12155 17920 12164
rect 17868 12121 17877 12155
rect 17877 12121 17911 12155
rect 17911 12121 17920 12155
rect 17868 12112 17920 12121
rect 18788 12112 18840 12164
rect 10876 12044 10928 12096
rect 11520 12044 11572 12096
rect 12440 12044 12492 12096
rect 12992 12044 13044 12096
rect 13360 12044 13412 12096
rect 14924 12044 14976 12096
rect 15384 12044 15436 12096
rect 16120 12087 16172 12096
rect 16120 12053 16129 12087
rect 16129 12053 16163 12087
rect 16163 12053 16172 12087
rect 16120 12044 16172 12053
rect 5502 11942 5554 11994
rect 5566 11942 5618 11994
rect 5630 11942 5682 11994
rect 5694 11942 5746 11994
rect 5758 11942 5810 11994
rect 5822 11942 5874 11994
rect 5886 11942 5938 11994
rect 5950 11942 6002 11994
rect 6014 11942 6066 11994
rect 6078 11942 6130 11994
rect 6142 11942 6194 11994
rect 6206 11942 6258 11994
rect 6270 11942 6322 11994
rect 6334 11942 6386 11994
rect 6398 11942 6450 11994
rect 6462 11942 6514 11994
rect 6526 11942 6578 11994
rect 6590 11942 6642 11994
rect 6654 11942 6706 11994
rect 13502 11942 13554 11994
rect 13566 11942 13618 11994
rect 13630 11942 13682 11994
rect 13694 11942 13746 11994
rect 13758 11942 13810 11994
rect 13822 11942 13874 11994
rect 13886 11942 13938 11994
rect 13950 11942 14002 11994
rect 14014 11942 14066 11994
rect 14078 11942 14130 11994
rect 14142 11942 14194 11994
rect 14206 11942 14258 11994
rect 14270 11942 14322 11994
rect 14334 11942 14386 11994
rect 14398 11942 14450 11994
rect 14462 11942 14514 11994
rect 14526 11942 14578 11994
rect 14590 11942 14642 11994
rect 14654 11942 14706 11994
rect 1400 11840 1452 11892
rect 2412 11772 2464 11824
rect 2596 11815 2648 11824
rect 2596 11781 2605 11815
rect 2605 11781 2639 11815
rect 2639 11781 2648 11815
rect 2596 11772 2648 11781
rect 2872 11815 2924 11824
rect 2872 11781 2881 11815
rect 2881 11781 2915 11815
rect 2915 11781 2924 11815
rect 2872 11772 2924 11781
rect 3148 11840 3200 11892
rect 3884 11840 3936 11892
rect 4620 11840 4672 11892
rect 3424 11772 3476 11824
rect 3792 11704 3844 11756
rect 4252 11704 4304 11756
rect 6368 11772 6420 11824
rect 4436 11636 4488 11688
rect 3516 11568 3568 11620
rect 4804 11704 4856 11756
rect 5172 11704 5224 11756
rect 5264 11704 5316 11756
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 5908 11704 5960 11756
rect 7196 11772 7248 11824
rect 6000 11636 6052 11688
rect 7564 11704 7616 11756
rect 7196 11636 7248 11688
rect 5264 11568 5316 11620
rect 1308 11500 1360 11552
rect 1768 11500 1820 11552
rect 3976 11500 4028 11552
rect 4620 11500 4672 11552
rect 6460 11568 6512 11620
rect 7012 11568 7064 11620
rect 7840 11772 7892 11824
rect 10048 11840 10100 11892
rect 8208 11636 8260 11688
rect 9680 11772 9732 11824
rect 9772 11772 9824 11824
rect 10508 11840 10560 11892
rect 11612 11840 11664 11892
rect 10784 11772 10836 11824
rect 11888 11772 11940 11824
rect 12992 11840 13044 11892
rect 13360 11840 13412 11892
rect 14556 11840 14608 11892
rect 14832 11840 14884 11892
rect 9404 11704 9456 11756
rect 8576 11568 8628 11620
rect 8944 11568 8996 11620
rect 9588 11636 9640 11688
rect 9772 11679 9824 11688
rect 9772 11645 9781 11679
rect 9781 11645 9815 11679
rect 9815 11645 9824 11679
rect 9772 11636 9824 11645
rect 10324 11704 10376 11756
rect 10692 11747 10744 11756
rect 10692 11713 10695 11747
rect 10695 11713 10744 11747
rect 13176 11772 13228 11824
rect 13268 11772 13320 11824
rect 10692 11704 10744 11713
rect 10876 11636 10928 11688
rect 12716 11704 12768 11756
rect 12992 11704 13044 11756
rect 15384 11772 15436 11824
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 18972 11772 19024 11824
rect 16212 11704 16264 11756
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 17132 11747 17184 11756
rect 17132 11713 17141 11747
rect 17141 11713 17175 11747
rect 17175 11713 17184 11747
rect 17132 11704 17184 11713
rect 17408 11704 17460 11756
rect 7656 11500 7708 11552
rect 7748 11500 7800 11552
rect 9404 11500 9456 11552
rect 11152 11500 11204 11552
rect 12532 11568 12584 11620
rect 15200 11636 15252 11688
rect 16488 11636 16540 11688
rect 14280 11568 14332 11620
rect 14832 11568 14884 11620
rect 15568 11568 15620 11620
rect 15844 11568 15896 11620
rect 12716 11500 12768 11552
rect 12808 11543 12860 11552
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 13268 11500 13320 11552
rect 16580 11500 16632 11552
rect 17868 11500 17920 11552
rect 1502 11398 1554 11450
rect 1566 11398 1618 11450
rect 1630 11398 1682 11450
rect 1694 11398 1746 11450
rect 1758 11398 1810 11450
rect 1822 11398 1874 11450
rect 1886 11398 1938 11450
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 2270 11398 2322 11450
rect 2334 11398 2386 11450
rect 2398 11398 2450 11450
rect 2462 11398 2514 11450
rect 2526 11398 2578 11450
rect 2590 11398 2642 11450
rect 2654 11398 2706 11450
rect 9502 11398 9554 11450
rect 9566 11398 9618 11450
rect 9630 11398 9682 11450
rect 9694 11398 9746 11450
rect 9758 11398 9810 11450
rect 9822 11398 9874 11450
rect 9886 11398 9938 11450
rect 9950 11398 10002 11450
rect 10014 11398 10066 11450
rect 10078 11398 10130 11450
rect 10142 11398 10194 11450
rect 10206 11398 10258 11450
rect 10270 11398 10322 11450
rect 10334 11398 10386 11450
rect 10398 11398 10450 11450
rect 10462 11398 10514 11450
rect 10526 11398 10578 11450
rect 10590 11398 10642 11450
rect 10654 11398 10706 11450
rect 17502 11398 17554 11450
rect 17566 11398 17618 11450
rect 17630 11398 17682 11450
rect 17694 11398 17746 11450
rect 17758 11398 17810 11450
rect 17822 11398 17874 11450
rect 17886 11398 17938 11450
rect 17950 11398 18002 11450
rect 18014 11398 18066 11450
rect 18078 11398 18130 11450
rect 18142 11398 18194 11450
rect 18206 11398 18258 11450
rect 18270 11398 18322 11450
rect 18334 11398 18386 11450
rect 18398 11398 18450 11450
rect 18462 11398 18514 11450
rect 18526 11398 18578 11450
rect 18590 11398 18642 11450
rect 18654 11398 18706 11450
rect 1768 11296 1820 11348
rect 3424 11296 3476 11348
rect 7012 11296 7064 11348
rect 7380 11296 7432 11348
rect 8208 11296 8260 11348
rect 9128 11296 9180 11348
rect 9220 11296 9272 11348
rect 9496 11296 9548 11348
rect 1400 11160 1452 11212
rect 4436 11228 4488 11280
rect 4804 11228 4856 11280
rect 5172 11271 5224 11280
rect 5172 11237 5181 11271
rect 5181 11237 5215 11271
rect 5215 11237 5224 11271
rect 5172 11228 5224 11237
rect 5908 11271 5960 11280
rect 5908 11237 5917 11271
rect 5917 11237 5951 11271
rect 5951 11237 5960 11271
rect 5908 11228 5960 11237
rect 6460 11271 6512 11280
rect 4620 11203 4672 11212
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 6460 11237 6469 11271
rect 6469 11237 6503 11271
rect 6503 11237 6512 11271
rect 6460 11228 6512 11237
rect 7196 11228 7248 11280
rect 7932 11228 7984 11280
rect 12072 11296 12124 11348
rect 14280 11339 14332 11348
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 15476 11296 15528 11348
rect 15660 11296 15712 11348
rect 2872 11092 2924 11144
rect 4068 11092 4120 11144
rect 4804 11092 4856 11144
rect 7748 11160 7800 11212
rect 8576 11160 8628 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 10692 11160 10744 11212
rect 1308 11024 1360 11076
rect 2228 11067 2280 11076
rect 2228 11033 2237 11067
rect 2237 11033 2271 11067
rect 2271 11033 2280 11067
rect 2228 11024 2280 11033
rect 3608 10956 3660 11008
rect 3976 10956 4028 11008
rect 4160 10956 4212 11008
rect 4620 11024 4672 11076
rect 6368 11024 6420 11076
rect 7564 11024 7616 11076
rect 8852 11092 8904 11144
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 9864 11092 9916 11144
rect 4712 10956 4764 11008
rect 7380 10956 7432 11008
rect 8024 11024 8076 11076
rect 9496 11024 9548 11076
rect 10692 11024 10744 11076
rect 11060 11160 11112 11212
rect 12348 11228 12400 11280
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 12164 11092 12216 11144
rect 14464 11160 14516 11212
rect 17132 11160 17184 11212
rect 11612 11024 11664 11076
rect 13176 11024 13228 11076
rect 14648 11092 14700 11144
rect 15108 11092 15160 11144
rect 14556 11024 14608 11076
rect 8116 10956 8168 11008
rect 8944 10956 8996 11008
rect 9036 10956 9088 11008
rect 9772 10956 9824 11008
rect 11888 10956 11940 11008
rect 12716 10956 12768 11008
rect 13360 10956 13412 11008
rect 15200 11024 15252 11076
rect 15384 11092 15436 11144
rect 16948 11092 17000 11144
rect 16856 11024 16908 11076
rect 17040 11024 17092 11076
rect 17132 10956 17184 11008
rect 5502 10854 5554 10906
rect 5566 10854 5618 10906
rect 5630 10854 5682 10906
rect 5694 10854 5746 10906
rect 5758 10854 5810 10906
rect 5822 10854 5874 10906
rect 5886 10854 5938 10906
rect 5950 10854 6002 10906
rect 6014 10854 6066 10906
rect 6078 10854 6130 10906
rect 6142 10854 6194 10906
rect 6206 10854 6258 10906
rect 6270 10854 6322 10906
rect 6334 10854 6386 10906
rect 6398 10854 6450 10906
rect 6462 10854 6514 10906
rect 6526 10854 6578 10906
rect 6590 10854 6642 10906
rect 6654 10854 6706 10906
rect 13502 10854 13554 10906
rect 13566 10854 13618 10906
rect 13630 10854 13682 10906
rect 13694 10854 13746 10906
rect 13758 10854 13810 10906
rect 13822 10854 13874 10906
rect 13886 10854 13938 10906
rect 13950 10854 14002 10906
rect 14014 10854 14066 10906
rect 14078 10854 14130 10906
rect 14142 10854 14194 10906
rect 14206 10854 14258 10906
rect 14270 10854 14322 10906
rect 14334 10854 14386 10906
rect 14398 10854 14450 10906
rect 14462 10854 14514 10906
rect 14526 10854 14578 10906
rect 14590 10854 14642 10906
rect 14654 10854 14706 10906
rect 1124 10752 1176 10804
rect 296 10684 348 10736
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 2228 10684 2280 10736
rect 3976 10752 4028 10804
rect 4620 10752 4672 10804
rect 4896 10752 4948 10804
rect 7472 10752 7524 10804
rect 8116 10752 8168 10804
rect 1860 10523 1912 10532
rect 1860 10489 1869 10523
rect 1869 10489 1903 10523
rect 1903 10489 1912 10523
rect 1860 10480 1912 10489
rect 1400 10412 1452 10464
rect 3608 10684 3660 10736
rect 4528 10684 4580 10736
rect 9220 10752 9272 10804
rect 9680 10752 9732 10804
rect 9588 10684 9640 10736
rect 3424 10616 3476 10668
rect 3792 10616 3844 10668
rect 4712 10616 4764 10668
rect 5448 10616 5500 10668
rect 19248 10752 19300 10804
rect 11336 10684 11388 10736
rect 11520 10684 11572 10736
rect 12072 10684 12124 10736
rect 12348 10659 12400 10668
rect 3884 10548 3936 10600
rect 4344 10548 4396 10600
rect 4988 10548 5040 10600
rect 5540 10591 5592 10600
rect 5540 10557 5565 10591
rect 5565 10557 5592 10591
rect 5540 10548 5592 10557
rect 7104 10591 7156 10600
rect 7104 10557 7120 10591
rect 7120 10557 7154 10591
rect 7154 10557 7156 10591
rect 7104 10548 7156 10557
rect 8668 10548 8720 10600
rect 8852 10548 8904 10600
rect 9312 10548 9364 10600
rect 12348 10625 12357 10659
rect 12357 10625 12400 10659
rect 12348 10616 12400 10625
rect 12532 10616 12584 10668
rect 12808 10616 12860 10668
rect 15200 10684 15252 10736
rect 6552 10480 6604 10532
rect 9956 10480 10008 10532
rect 10876 10548 10928 10600
rect 12164 10548 12216 10600
rect 12624 10591 12676 10600
rect 12624 10557 12633 10591
rect 12633 10557 12667 10591
rect 12667 10557 12676 10591
rect 12624 10548 12676 10557
rect 13360 10591 13412 10600
rect 13360 10557 13369 10591
rect 13369 10557 13403 10591
rect 13403 10557 13412 10591
rect 13360 10548 13412 10557
rect 14280 10591 14332 10600
rect 14280 10557 14289 10591
rect 14289 10557 14323 10591
rect 14323 10557 14332 10591
rect 14280 10548 14332 10557
rect 14464 10548 14516 10600
rect 15384 10616 15436 10668
rect 16212 10616 16264 10668
rect 16396 10616 16448 10668
rect 16948 10548 17000 10600
rect 17224 10548 17276 10600
rect 17408 10548 17460 10600
rect 18880 10548 18932 10600
rect 11428 10480 11480 10532
rect 11888 10480 11940 10532
rect 15660 10523 15712 10532
rect 15660 10489 15669 10523
rect 15669 10489 15703 10523
rect 15703 10489 15712 10523
rect 15660 10480 15712 10489
rect 3148 10412 3200 10464
rect 3976 10412 4028 10464
rect 5264 10412 5316 10464
rect 6828 10412 6880 10464
rect 7380 10455 7432 10464
rect 7380 10421 7410 10455
rect 7410 10421 7432 10455
rect 7380 10412 7432 10421
rect 7932 10412 7984 10464
rect 8484 10412 8536 10464
rect 8668 10412 8720 10464
rect 9772 10412 9824 10464
rect 10140 10412 10192 10464
rect 12624 10412 12676 10464
rect 13360 10412 13412 10464
rect 15016 10412 15068 10464
rect 16028 10412 16080 10464
rect 16304 10412 16356 10464
rect 17224 10412 17276 10464
rect 1502 10310 1554 10362
rect 1566 10310 1618 10362
rect 1630 10310 1682 10362
rect 1694 10310 1746 10362
rect 1758 10310 1810 10362
rect 1822 10310 1874 10362
rect 1886 10310 1938 10362
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 2270 10310 2322 10362
rect 2334 10310 2386 10362
rect 2398 10310 2450 10362
rect 2462 10310 2514 10362
rect 2526 10310 2578 10362
rect 2590 10310 2642 10362
rect 2654 10310 2706 10362
rect 9502 10310 9554 10362
rect 9566 10310 9618 10362
rect 9630 10310 9682 10362
rect 9694 10310 9746 10362
rect 9758 10310 9810 10362
rect 9822 10310 9874 10362
rect 9886 10310 9938 10362
rect 9950 10310 10002 10362
rect 10014 10310 10066 10362
rect 10078 10310 10130 10362
rect 10142 10310 10194 10362
rect 10206 10310 10258 10362
rect 10270 10310 10322 10362
rect 10334 10310 10386 10362
rect 10398 10310 10450 10362
rect 10462 10310 10514 10362
rect 10526 10310 10578 10362
rect 10590 10310 10642 10362
rect 10654 10310 10706 10362
rect 17502 10310 17554 10362
rect 17566 10310 17618 10362
rect 17630 10310 17682 10362
rect 17694 10310 17746 10362
rect 17758 10310 17810 10362
rect 17822 10310 17874 10362
rect 17886 10310 17938 10362
rect 17950 10310 18002 10362
rect 18014 10310 18066 10362
rect 18078 10310 18130 10362
rect 18142 10310 18194 10362
rect 18206 10310 18258 10362
rect 18270 10310 18322 10362
rect 18334 10310 18386 10362
rect 18398 10310 18450 10362
rect 18462 10310 18514 10362
rect 18526 10310 18578 10362
rect 18590 10310 18642 10362
rect 18654 10310 18706 10362
rect 2596 10208 2648 10260
rect 2872 10208 2924 10260
rect 3148 10208 3200 10260
rect 4896 10208 4948 10260
rect 4988 10208 5040 10260
rect 10508 10208 10560 10260
rect 3332 10140 3384 10192
rect 2320 10072 2372 10124
rect 2872 10004 2924 10056
rect 3148 10004 3200 10056
rect 3332 10004 3384 10056
rect 4712 10004 4764 10056
rect 5448 10004 5500 10056
rect 12164 10208 12216 10260
rect 14648 10208 14700 10260
rect 16304 10208 16356 10260
rect 17132 10208 17184 10260
rect 17500 10208 17552 10260
rect 6920 10072 6972 10124
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 1032 9936 1084 9988
rect 2412 9936 2464 9988
rect 2688 9979 2740 9988
rect 2688 9945 2697 9979
rect 2697 9945 2731 9979
rect 2731 9945 2740 9979
rect 2688 9936 2740 9945
rect 8576 10072 8628 10124
rect 9128 10072 9180 10124
rect 17224 10140 17276 10192
rect 18696 10140 18748 10192
rect 8116 9936 8168 9988
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 11336 10004 11388 10056
rect 12532 10004 12584 10056
rect 15016 10072 15068 10124
rect 1216 9868 1268 9920
rect 4988 9868 5040 9920
rect 6644 9868 6696 9920
rect 9128 9979 9180 9988
rect 9128 9945 9137 9979
rect 9137 9945 9171 9979
rect 9171 9945 9180 9979
rect 9128 9936 9180 9945
rect 10876 9936 10928 9988
rect 11244 9936 11296 9988
rect 11704 9979 11756 9988
rect 11704 9945 11713 9979
rect 11713 9945 11747 9979
rect 11747 9945 11756 9979
rect 11704 9936 11756 9945
rect 12072 9936 12124 9988
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 15384 10072 15436 10124
rect 17132 10072 17184 10124
rect 18788 10072 18840 10124
rect 15200 10004 15252 10056
rect 17040 9936 17092 9988
rect 11060 9868 11112 9920
rect 13268 9868 13320 9920
rect 14832 9868 14884 9920
rect 15292 9868 15344 9920
rect 15936 9868 15988 9920
rect 16396 9868 16448 9920
rect 17408 9936 17460 9988
rect 18788 9936 18840 9988
rect 17224 9911 17276 9920
rect 17224 9877 17233 9911
rect 17233 9877 17267 9911
rect 17267 9877 17276 9911
rect 17224 9868 17276 9877
rect 18052 9868 18104 9920
rect 296 9800 348 9852
rect 848 9800 900 9852
rect 5502 9766 5554 9818
rect 5566 9766 5618 9818
rect 5630 9766 5682 9818
rect 5694 9766 5746 9818
rect 5758 9766 5810 9818
rect 5822 9766 5874 9818
rect 5886 9766 5938 9818
rect 5950 9766 6002 9818
rect 6014 9766 6066 9818
rect 6078 9766 6130 9818
rect 6142 9766 6194 9818
rect 6206 9766 6258 9818
rect 6270 9766 6322 9818
rect 6334 9766 6386 9818
rect 6398 9766 6450 9818
rect 6462 9766 6514 9818
rect 6526 9766 6578 9818
rect 6590 9766 6642 9818
rect 6654 9766 6706 9818
rect 13502 9766 13554 9818
rect 13566 9766 13618 9818
rect 13630 9766 13682 9818
rect 13694 9766 13746 9818
rect 13758 9766 13810 9818
rect 13822 9766 13874 9818
rect 13886 9766 13938 9818
rect 13950 9766 14002 9818
rect 14014 9766 14066 9818
rect 14078 9766 14130 9818
rect 14142 9766 14194 9818
rect 14206 9766 14258 9818
rect 14270 9766 14322 9818
rect 14334 9766 14386 9818
rect 14398 9766 14450 9818
rect 14462 9766 14514 9818
rect 14526 9766 14578 9818
rect 14590 9766 14642 9818
rect 14654 9766 14706 9818
rect 112 9664 164 9716
rect 3976 9664 4028 9716
rect 5080 9664 5132 9716
rect 5356 9707 5408 9716
rect 5356 9673 5365 9707
rect 5365 9673 5399 9707
rect 5399 9673 5408 9707
rect 5356 9664 5408 9673
rect 2688 9596 2740 9648
rect 4528 9596 4580 9648
rect 4712 9596 4764 9648
rect 2320 9571 2372 9580
rect 572 9460 624 9512
rect 1032 9460 1084 9512
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 2412 9528 2464 9580
rect 5264 9528 5316 9580
rect 6920 9664 6972 9716
rect 10784 9664 10836 9716
rect 11336 9664 11388 9716
rect 11704 9664 11756 9716
rect 12164 9664 12216 9716
rect 12716 9664 12768 9716
rect 8116 9596 8168 9648
rect 9128 9596 9180 9648
rect 10508 9596 10560 9648
rect 12348 9596 12400 9648
rect 12992 9596 13044 9648
rect 7288 9528 7340 9580
rect 2780 9460 2832 9512
rect 3148 9460 3200 9512
rect 5356 9460 5408 9512
rect 6920 9460 6972 9512
rect 8024 9460 8076 9512
rect 11428 9528 11480 9580
rect 12532 9528 12584 9580
rect 12624 9528 12676 9580
rect 14832 9528 14884 9580
rect 12440 9460 12492 9512
rect 14464 9503 14516 9512
rect 6552 9392 6604 9444
rect 10692 9392 10744 9444
rect 11060 9392 11112 9444
rect 11704 9392 11756 9444
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 2596 9324 2648 9376
rect 3148 9324 3200 9376
rect 4712 9367 4764 9376
rect 4712 9333 4721 9367
rect 4721 9333 4755 9367
rect 4755 9333 4764 9367
rect 4712 9324 4764 9333
rect 7288 9324 7340 9376
rect 8024 9324 8076 9376
rect 12348 9324 12400 9376
rect 12808 9324 12860 9376
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 15108 9664 15160 9716
rect 17316 9639 17368 9648
rect 17316 9605 17325 9639
rect 17325 9605 17359 9639
rect 17359 9605 17368 9639
rect 17316 9596 17368 9605
rect 15752 9460 15804 9512
rect 13544 9392 13596 9444
rect 14188 9392 14240 9444
rect 16212 9528 16264 9580
rect 16672 9528 16724 9580
rect 19340 9596 19392 9648
rect 17500 9528 17552 9580
rect 16396 9460 16448 9512
rect 16948 9460 17000 9512
rect 16672 9392 16724 9444
rect 17040 9392 17092 9444
rect 17960 9435 18012 9444
rect 17960 9401 17969 9435
rect 17969 9401 18003 9435
rect 18003 9401 18012 9435
rect 17960 9392 18012 9401
rect 14096 9324 14148 9376
rect 15752 9324 15804 9376
rect 18052 9324 18104 9376
rect 1502 9222 1554 9274
rect 1566 9222 1618 9274
rect 1630 9222 1682 9274
rect 1694 9222 1746 9274
rect 1758 9222 1810 9274
rect 1822 9222 1874 9274
rect 1886 9222 1938 9274
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 2270 9222 2322 9274
rect 2334 9222 2386 9274
rect 2398 9222 2450 9274
rect 2462 9222 2514 9274
rect 2526 9222 2578 9274
rect 2590 9222 2642 9274
rect 2654 9222 2706 9274
rect 9502 9222 9554 9274
rect 9566 9222 9618 9274
rect 9630 9222 9682 9274
rect 9694 9222 9746 9274
rect 9758 9222 9810 9274
rect 9822 9222 9874 9274
rect 9886 9222 9938 9274
rect 9950 9222 10002 9274
rect 10014 9222 10066 9274
rect 10078 9222 10130 9274
rect 10142 9222 10194 9274
rect 10206 9222 10258 9274
rect 10270 9222 10322 9274
rect 10334 9222 10386 9274
rect 10398 9222 10450 9274
rect 10462 9222 10514 9274
rect 10526 9222 10578 9274
rect 10590 9222 10642 9274
rect 10654 9222 10706 9274
rect 17502 9222 17554 9274
rect 17566 9222 17618 9274
rect 17630 9222 17682 9274
rect 17694 9222 17746 9274
rect 17758 9222 17810 9274
rect 17822 9222 17874 9274
rect 17886 9222 17938 9274
rect 17950 9222 18002 9274
rect 18014 9222 18066 9274
rect 18078 9222 18130 9274
rect 18142 9222 18194 9274
rect 18206 9222 18258 9274
rect 18270 9222 18322 9274
rect 18334 9222 18386 9274
rect 18398 9222 18450 9274
rect 18462 9222 18514 9274
rect 18526 9222 18578 9274
rect 18590 9222 18642 9274
rect 18654 9222 18706 9274
rect 5264 9120 5316 9172
rect 9956 9120 10008 9172
rect 12348 9120 12400 9172
rect 12532 9120 12584 9172
rect 12992 9120 13044 9172
rect 15108 9120 15160 9172
rect 17132 9120 17184 9172
rect 3056 9052 3108 9104
rect 2872 8984 2924 9036
rect 2964 8916 3016 8968
rect 3056 8916 3108 8968
rect 7748 9052 7800 9104
rect 13176 9052 13228 9104
rect 13452 9052 13504 9104
rect 2228 8848 2280 8900
rect 2688 8891 2740 8900
rect 2688 8857 2697 8891
rect 2697 8857 2731 8891
rect 2731 8857 2740 8891
rect 2688 8848 2740 8857
rect 2780 8891 2832 8900
rect 2780 8857 2789 8891
rect 2789 8857 2823 8891
rect 2823 8857 2832 8891
rect 2780 8848 2832 8857
rect 4436 8848 4488 8900
rect 5264 8848 5316 8900
rect 3332 8780 3384 8832
rect 9496 8984 9548 9036
rect 10692 8984 10744 9036
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 8116 8848 8168 8900
rect 11060 8916 11112 8968
rect 15200 8984 15252 9036
rect 17684 8984 17736 9036
rect 18052 9027 18104 9036
rect 18052 8993 18061 9027
rect 18061 8993 18095 9027
rect 18095 8993 18104 9027
rect 18052 8984 18104 8993
rect 14188 8916 14240 8968
rect 15660 8916 15712 8968
rect 16672 8959 16724 8968
rect 16672 8925 16681 8959
rect 16681 8925 16715 8959
rect 16715 8925 16724 8959
rect 16672 8916 16724 8925
rect 11888 8891 11940 8900
rect 11888 8857 11897 8891
rect 11897 8857 11931 8891
rect 11931 8857 11940 8891
rect 11888 8848 11940 8857
rect 13176 8848 13228 8900
rect 14096 8848 14148 8900
rect 14648 8848 14700 8900
rect 16396 8848 16448 8900
rect 17224 8916 17276 8968
rect 17592 8916 17644 8968
rect 17960 8959 18012 8968
rect 17960 8925 17969 8959
rect 17969 8925 18003 8959
rect 18003 8925 18012 8959
rect 17960 8916 18012 8925
rect 18972 8916 19024 8968
rect 17040 8848 17092 8900
rect 9220 8823 9272 8832
rect 9220 8789 9229 8823
rect 9229 8789 9263 8823
rect 9263 8789 9272 8823
rect 9220 8780 9272 8789
rect 10968 8823 11020 8832
rect 10968 8789 10977 8823
rect 10977 8789 11011 8823
rect 11011 8789 11020 8823
rect 10968 8780 11020 8789
rect 11060 8780 11112 8832
rect 14464 8780 14516 8832
rect 16672 8823 16724 8832
rect 16672 8789 16681 8823
rect 16681 8789 16715 8823
rect 16715 8789 16724 8823
rect 16672 8780 16724 8789
rect 5502 8678 5554 8730
rect 5566 8678 5618 8730
rect 5630 8678 5682 8730
rect 5694 8678 5746 8730
rect 5758 8678 5810 8730
rect 5822 8678 5874 8730
rect 5886 8678 5938 8730
rect 5950 8678 6002 8730
rect 6014 8678 6066 8730
rect 6078 8678 6130 8730
rect 6142 8678 6194 8730
rect 6206 8678 6258 8730
rect 6270 8678 6322 8730
rect 6334 8678 6386 8730
rect 6398 8678 6450 8730
rect 6462 8678 6514 8730
rect 6526 8678 6578 8730
rect 6590 8678 6642 8730
rect 6654 8678 6706 8730
rect 13502 8678 13554 8730
rect 13566 8678 13618 8730
rect 13630 8678 13682 8730
rect 13694 8678 13746 8730
rect 13758 8678 13810 8730
rect 13822 8678 13874 8730
rect 13886 8678 13938 8730
rect 13950 8678 14002 8730
rect 14014 8678 14066 8730
rect 14078 8678 14130 8730
rect 14142 8678 14194 8730
rect 14206 8678 14258 8730
rect 14270 8678 14322 8730
rect 14334 8678 14386 8730
rect 14398 8678 14450 8730
rect 14462 8678 14514 8730
rect 14526 8678 14578 8730
rect 14590 8678 14642 8730
rect 14654 8678 14706 8730
rect 2688 8576 2740 8628
rect 4436 8576 4488 8628
rect 5448 8576 5500 8628
rect 2228 8508 2280 8560
rect 2872 8440 2924 8492
rect 4252 8508 4304 8560
rect 4528 8440 4580 8492
rect 5080 8440 5132 8492
rect 5264 8440 5316 8492
rect 7748 8576 7800 8628
rect 8116 8508 8168 8560
rect 9220 8508 9272 8560
rect 2780 8372 2832 8424
rect 3056 8304 3108 8356
rect 3608 8304 3660 8356
rect 5080 8304 5132 8356
rect 5264 8304 5316 8356
rect 7288 8440 7340 8492
rect 9036 8440 9088 8492
rect 12808 8576 12860 8628
rect 13360 8576 13412 8628
rect 12624 8508 12676 8560
rect 15016 8619 15068 8628
rect 15016 8585 15025 8619
rect 15025 8585 15059 8619
rect 15059 8585 15068 8619
rect 15016 8576 15068 8585
rect 15660 8576 15712 8628
rect 16396 8576 16448 8628
rect 17316 8576 17368 8628
rect 17960 8576 18012 8628
rect 18144 8619 18196 8628
rect 18144 8585 18153 8619
rect 18153 8585 18187 8619
rect 18187 8585 18196 8619
rect 18144 8576 18196 8585
rect 16672 8508 16724 8560
rect 17592 8551 17644 8560
rect 17592 8517 17601 8551
rect 17601 8517 17635 8551
rect 17635 8517 17644 8551
rect 17592 8508 17644 8517
rect 9956 8372 10008 8424
rect 11704 8304 11756 8356
rect 14832 8440 14884 8492
rect 13544 8372 13596 8424
rect 15200 8372 15252 8424
rect 17408 8440 17460 8492
rect 18052 8440 18104 8492
rect 18788 8440 18840 8492
rect 18972 8372 19024 8424
rect 15108 8304 15160 8356
rect 16396 8304 16448 8356
rect 17500 8304 17552 8356
rect 7196 8236 7248 8288
rect 12256 8236 12308 8288
rect 12624 8236 12676 8288
rect 13176 8236 13228 8288
rect 13360 8236 13412 8288
rect 14832 8236 14884 8288
rect 15384 8236 15436 8288
rect 16672 8236 16724 8288
rect 17132 8236 17184 8288
rect 17684 8236 17736 8288
rect 1502 8134 1554 8186
rect 1566 8134 1618 8186
rect 1630 8134 1682 8186
rect 1694 8134 1746 8186
rect 1758 8134 1810 8186
rect 1822 8134 1874 8186
rect 1886 8134 1938 8186
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 2270 8134 2322 8186
rect 2334 8134 2386 8186
rect 2398 8134 2450 8186
rect 2462 8134 2514 8186
rect 2526 8134 2578 8186
rect 2590 8134 2642 8186
rect 2654 8134 2706 8186
rect 9502 8134 9554 8186
rect 9566 8134 9618 8186
rect 9630 8134 9682 8186
rect 9694 8134 9746 8186
rect 9758 8134 9810 8186
rect 9822 8134 9874 8186
rect 9886 8134 9938 8186
rect 9950 8134 10002 8186
rect 10014 8134 10066 8186
rect 10078 8134 10130 8186
rect 10142 8134 10194 8186
rect 10206 8134 10258 8186
rect 10270 8134 10322 8186
rect 10334 8134 10386 8186
rect 10398 8134 10450 8186
rect 10462 8134 10514 8186
rect 10526 8134 10578 8186
rect 10590 8134 10642 8186
rect 10654 8134 10706 8186
rect 17502 8134 17554 8186
rect 17566 8134 17618 8186
rect 17630 8134 17682 8186
rect 17694 8134 17746 8186
rect 17758 8134 17810 8186
rect 17822 8134 17874 8186
rect 17886 8134 17938 8186
rect 17950 8134 18002 8186
rect 18014 8134 18066 8186
rect 18078 8134 18130 8186
rect 18142 8134 18194 8186
rect 18206 8134 18258 8186
rect 18270 8134 18322 8186
rect 18334 8134 18386 8186
rect 18398 8134 18450 8186
rect 18462 8134 18514 8186
rect 18526 8134 18578 8186
rect 18590 8134 18642 8186
rect 18654 8134 18706 8186
rect 388 8032 440 8084
rect 940 8032 992 8084
rect 1308 8032 1360 8084
rect 2136 8032 2188 8084
rect 11612 8032 11664 8084
rect 3700 7964 3752 8016
rect 2872 7896 2924 7948
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 3700 7828 3752 7880
rect 6828 7896 6880 7948
rect 7840 7896 7892 7948
rect 7196 7828 7248 7880
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 2688 7803 2740 7812
rect 2688 7769 2697 7803
rect 2697 7769 2731 7803
rect 2731 7769 2740 7803
rect 2688 7760 2740 7769
rect 2780 7803 2832 7812
rect 2780 7769 2789 7803
rect 2789 7769 2823 7803
rect 2823 7769 2832 7803
rect 2780 7760 2832 7769
rect 8116 7760 8168 7812
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 3056 7692 3108 7744
rect 9404 7760 9456 7812
rect 9956 7803 10008 7812
rect 9956 7769 9965 7803
rect 9965 7769 9999 7803
rect 9999 7769 10008 7803
rect 9956 7760 10008 7769
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 11428 7896 11480 7948
rect 12532 8032 12584 8084
rect 12716 8032 12768 8084
rect 12624 7964 12676 8016
rect 17132 8032 17184 8084
rect 17316 8075 17368 8084
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 12532 7896 12584 7948
rect 13544 7896 13596 7948
rect 15844 7939 15896 7948
rect 15844 7905 15853 7939
rect 15853 7905 15887 7939
rect 15887 7905 15896 7939
rect 15844 7896 15896 7905
rect 17040 7896 17092 7948
rect 12808 7828 12860 7880
rect 13084 7828 13136 7880
rect 12072 7760 12124 7812
rect 14556 7871 14608 7880
rect 14556 7837 14565 7871
rect 14565 7837 14599 7871
rect 14599 7837 14608 7871
rect 14556 7828 14608 7837
rect 15292 7828 15344 7880
rect 16856 7760 16908 7812
rect 12716 7692 12768 7744
rect 14096 7692 14148 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 5502 7590 5554 7642
rect 5566 7590 5618 7642
rect 5630 7590 5682 7642
rect 5694 7590 5746 7642
rect 5758 7590 5810 7642
rect 5822 7590 5874 7642
rect 5886 7590 5938 7642
rect 5950 7590 6002 7642
rect 6014 7590 6066 7642
rect 6078 7590 6130 7642
rect 6142 7590 6194 7642
rect 6206 7590 6258 7642
rect 6270 7590 6322 7642
rect 6334 7590 6386 7642
rect 6398 7590 6450 7642
rect 6462 7590 6514 7642
rect 6526 7590 6578 7642
rect 6590 7590 6642 7642
rect 6654 7590 6706 7642
rect 13502 7590 13554 7642
rect 13566 7590 13618 7642
rect 13630 7590 13682 7642
rect 13694 7590 13746 7642
rect 13758 7590 13810 7642
rect 13822 7590 13874 7642
rect 13886 7590 13938 7642
rect 13950 7590 14002 7642
rect 14014 7590 14066 7642
rect 14078 7590 14130 7642
rect 14142 7590 14194 7642
rect 14206 7590 14258 7642
rect 14270 7590 14322 7642
rect 14334 7590 14386 7642
rect 14398 7590 14450 7642
rect 14462 7590 14514 7642
rect 14526 7590 14578 7642
rect 14590 7590 14642 7642
rect 14654 7590 14706 7642
rect 19340 7624 19392 7676
rect 2688 7488 2740 7540
rect 4896 7488 4948 7540
rect 5632 7488 5684 7540
rect 6920 7488 6972 7540
rect 7288 7488 7340 7540
rect 2964 7420 3016 7472
rect 3056 7463 3108 7472
rect 3056 7429 3065 7463
rect 3065 7429 3099 7463
rect 3099 7429 3108 7463
rect 3056 7420 3108 7429
rect 8116 7420 8168 7472
rect 9220 7420 9272 7472
rect 2872 7352 2924 7404
rect 2136 7148 2188 7200
rect 3700 7284 3752 7336
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 6828 7352 6880 7404
rect 7288 7352 7340 7404
rect 7748 7352 7800 7404
rect 11244 7488 11296 7540
rect 13084 7488 13136 7540
rect 9772 7420 9824 7472
rect 11060 7420 11112 7472
rect 12256 7420 12308 7472
rect 17960 7488 18012 7540
rect 16488 7420 16540 7472
rect 17224 7420 17276 7472
rect 19064 7420 19116 7472
rect 9956 7352 10008 7404
rect 11612 7352 11664 7404
rect 11060 7284 11112 7336
rect 6920 7216 6972 7268
rect 12624 7216 12676 7268
rect 11244 7148 11296 7200
rect 13268 7284 13320 7336
rect 14004 7327 14056 7336
rect 14004 7293 14013 7327
rect 14013 7293 14047 7327
rect 14047 7293 14056 7327
rect 14004 7284 14056 7293
rect 14740 7148 14792 7200
rect 17408 7148 17460 7200
rect 1502 7046 1554 7098
rect 1566 7046 1618 7098
rect 1630 7046 1682 7098
rect 1694 7046 1746 7098
rect 1758 7046 1810 7098
rect 1822 7046 1874 7098
rect 1886 7046 1938 7098
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 2270 7046 2322 7098
rect 2334 7046 2386 7098
rect 2398 7046 2450 7098
rect 2462 7046 2514 7098
rect 2526 7046 2578 7098
rect 2590 7046 2642 7098
rect 2654 7046 2706 7098
rect 9502 7046 9554 7098
rect 9566 7046 9618 7098
rect 9630 7046 9682 7098
rect 9694 7046 9746 7098
rect 9758 7046 9810 7098
rect 9822 7046 9874 7098
rect 9886 7046 9938 7098
rect 9950 7046 10002 7098
rect 10014 7046 10066 7098
rect 10078 7046 10130 7098
rect 10142 7046 10194 7098
rect 10206 7046 10258 7098
rect 10270 7046 10322 7098
rect 10334 7046 10386 7098
rect 10398 7046 10450 7098
rect 10462 7046 10514 7098
rect 10526 7046 10578 7098
rect 10590 7046 10642 7098
rect 10654 7046 10706 7098
rect 17502 7046 17554 7098
rect 17566 7046 17618 7098
rect 17630 7046 17682 7098
rect 17694 7046 17746 7098
rect 17758 7046 17810 7098
rect 17822 7046 17874 7098
rect 17886 7046 17938 7098
rect 17950 7046 18002 7098
rect 18014 7046 18066 7098
rect 18078 7046 18130 7098
rect 18142 7046 18194 7098
rect 18206 7046 18258 7098
rect 18270 7046 18322 7098
rect 18334 7046 18386 7098
rect 18398 7046 18450 7098
rect 18462 7046 18514 7098
rect 18526 7046 18578 7098
rect 18590 7046 18642 7098
rect 18654 7046 18706 7098
rect 1400 6944 1452 6996
rect 3332 6944 3384 6996
rect 8484 6944 8536 6996
rect 11152 6944 11204 6996
rect 11612 6944 11664 6996
rect 17408 6944 17460 6996
rect 2780 6808 2832 6860
rect 3148 6740 3200 6792
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 12532 6876 12584 6928
rect 13268 6876 13320 6928
rect 14004 6876 14056 6928
rect 15844 6876 15896 6928
rect 16304 6876 16356 6928
rect 13084 6808 13136 6860
rect 2228 6672 2280 6724
rect 2688 6715 2740 6724
rect 2688 6681 2697 6715
rect 2697 6681 2731 6715
rect 2731 6681 2740 6715
rect 2688 6672 2740 6681
rect 2964 6672 3016 6724
rect 3240 6604 3292 6656
rect 6920 6740 6972 6792
rect 7288 6783 7340 6792
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 7472 6672 7524 6724
rect 7932 6672 7984 6724
rect 8116 6672 8168 6724
rect 12072 6740 12124 6792
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 12532 6740 12584 6792
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 15292 6808 15344 6860
rect 16212 6808 16264 6860
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 14832 6672 14884 6724
rect 15568 6672 15620 6724
rect 17776 6783 17828 6792
rect 17776 6749 17785 6783
rect 17785 6749 17819 6783
rect 17819 6749 17828 6783
rect 17776 6740 17828 6749
rect 11796 6604 11848 6656
rect 12256 6604 12308 6656
rect 16028 6647 16080 6656
rect 16028 6613 16037 6647
rect 16037 6613 16071 6647
rect 16071 6613 16080 6647
rect 16028 6604 16080 6613
rect 5502 6502 5554 6554
rect 5566 6502 5618 6554
rect 5630 6502 5682 6554
rect 5694 6502 5746 6554
rect 5758 6502 5810 6554
rect 5822 6502 5874 6554
rect 5886 6502 5938 6554
rect 5950 6502 6002 6554
rect 6014 6502 6066 6554
rect 6078 6502 6130 6554
rect 6142 6502 6194 6554
rect 6206 6502 6258 6554
rect 6270 6502 6322 6554
rect 6334 6502 6386 6554
rect 6398 6502 6450 6554
rect 6462 6502 6514 6554
rect 6526 6502 6578 6554
rect 6590 6502 6642 6554
rect 6654 6502 6706 6554
rect 13502 6502 13554 6554
rect 13566 6502 13618 6554
rect 13630 6502 13682 6554
rect 13694 6502 13746 6554
rect 13758 6502 13810 6554
rect 13822 6502 13874 6554
rect 13886 6502 13938 6554
rect 13950 6502 14002 6554
rect 14014 6502 14066 6554
rect 14078 6502 14130 6554
rect 14142 6502 14194 6554
rect 14206 6502 14258 6554
rect 14270 6502 14322 6554
rect 14334 6502 14386 6554
rect 14398 6502 14450 6554
rect 14462 6502 14514 6554
rect 14526 6502 14578 6554
rect 14590 6502 14642 6554
rect 14654 6502 14706 6554
rect 2688 6400 2740 6452
rect 5080 6400 5132 6452
rect 2228 6332 2280 6384
rect 2780 6264 2832 6316
rect 5264 6375 5316 6384
rect 5264 6341 5273 6375
rect 5273 6341 5307 6375
rect 5307 6341 5316 6375
rect 5264 6332 5316 6341
rect 4528 6264 4580 6316
rect 4896 6264 4948 6316
rect 7748 6400 7800 6452
rect 12992 6400 13044 6452
rect 8116 6332 8168 6384
rect 9220 6332 9272 6384
rect 11060 6332 11112 6384
rect 11428 6332 11480 6384
rect 15016 6400 15068 6452
rect 15384 6400 15436 6452
rect 17224 6400 17276 6452
rect 2872 6196 2924 6248
rect 3148 6196 3200 6248
rect 4436 6196 4488 6248
rect 5264 6196 5316 6248
rect 7288 6264 7340 6316
rect 6828 6196 6880 6248
rect 7472 6196 7524 6248
rect 7932 6264 7984 6316
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 12532 6264 12584 6316
rect 14556 6332 14608 6384
rect 14372 6264 14424 6316
rect 15108 6332 15160 6384
rect 11244 6196 11296 6248
rect 11428 6196 11480 6248
rect 12256 6196 12308 6248
rect 12440 6196 12492 6248
rect 13268 6196 13320 6248
rect 6552 6128 6604 6180
rect 6828 6060 6880 6112
rect 7104 6060 7156 6112
rect 12624 6060 12676 6112
rect 13360 6060 13412 6112
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 15660 6264 15712 6316
rect 16212 6332 16264 6384
rect 18788 6332 18840 6384
rect 15936 6307 15988 6316
rect 15936 6273 15945 6307
rect 15945 6273 15979 6307
rect 15979 6273 15988 6307
rect 15936 6264 15988 6273
rect 16028 6264 16080 6316
rect 17776 6264 17828 6316
rect 14648 6171 14700 6180
rect 14648 6137 14657 6171
rect 14657 6137 14691 6171
rect 14691 6137 14700 6171
rect 14648 6128 14700 6137
rect 17040 6128 17092 6180
rect 15016 6060 15068 6112
rect 16948 6060 17000 6112
rect 1502 5958 1554 6010
rect 1566 5958 1618 6010
rect 1630 5958 1682 6010
rect 1694 5958 1746 6010
rect 1758 5958 1810 6010
rect 1822 5958 1874 6010
rect 1886 5958 1938 6010
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 2270 5958 2322 6010
rect 2334 5958 2386 6010
rect 2398 5958 2450 6010
rect 2462 5958 2514 6010
rect 2526 5958 2578 6010
rect 2590 5958 2642 6010
rect 2654 5958 2706 6010
rect 9502 5958 9554 6010
rect 9566 5958 9618 6010
rect 9630 5958 9682 6010
rect 9694 5958 9746 6010
rect 9758 5958 9810 6010
rect 9822 5958 9874 6010
rect 9886 5958 9938 6010
rect 9950 5958 10002 6010
rect 10014 5958 10066 6010
rect 10078 5958 10130 6010
rect 10142 5958 10194 6010
rect 10206 5958 10258 6010
rect 10270 5958 10322 6010
rect 10334 5958 10386 6010
rect 10398 5958 10450 6010
rect 10462 5958 10514 6010
rect 10526 5958 10578 6010
rect 10590 5958 10642 6010
rect 10654 5958 10706 6010
rect 17502 5958 17554 6010
rect 17566 5958 17618 6010
rect 17630 5958 17682 6010
rect 17694 5958 17746 6010
rect 17758 5958 17810 6010
rect 17822 5958 17874 6010
rect 17886 5958 17938 6010
rect 17950 5958 18002 6010
rect 18014 5958 18066 6010
rect 18078 5958 18130 6010
rect 18142 5958 18194 6010
rect 18206 5958 18258 6010
rect 18270 5958 18322 6010
rect 18334 5958 18386 6010
rect 18398 5958 18450 6010
rect 18462 5958 18514 6010
rect 18526 5958 18578 6010
rect 18590 5958 18642 6010
rect 18654 5958 18706 6010
rect 3608 5856 3660 5908
rect 4896 5856 4948 5908
rect 2872 5788 2924 5840
rect 4160 5720 4212 5772
rect 6920 5720 6972 5772
rect 7840 5720 7892 5772
rect 8300 5856 8352 5908
rect 11428 5856 11480 5908
rect 11980 5856 12032 5908
rect 12256 5856 12308 5908
rect 14372 5899 14424 5908
rect 14372 5865 14381 5899
rect 14381 5865 14415 5899
rect 14415 5865 14424 5899
rect 14372 5856 14424 5865
rect 12348 5788 12400 5840
rect 11152 5720 11204 5772
rect 11796 5763 11848 5772
rect 11796 5729 11805 5763
rect 11805 5729 11839 5763
rect 11839 5729 11848 5763
rect 11796 5720 11848 5729
rect 12900 5720 12952 5772
rect 13084 5720 13136 5772
rect 15108 5720 15160 5772
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 16028 5720 16080 5772
rect 17040 5899 17092 5908
rect 17040 5865 17049 5899
rect 17049 5865 17083 5899
rect 17083 5865 17092 5899
rect 17040 5856 17092 5865
rect 17224 5856 17276 5908
rect 17408 5788 17460 5840
rect 3332 5652 3384 5704
rect 2320 5584 2372 5636
rect 3516 5584 3568 5636
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 8116 5584 8168 5636
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 13360 5652 13412 5704
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 15200 5652 15252 5704
rect 3056 5516 3108 5568
rect 9128 5627 9180 5636
rect 9128 5593 9137 5627
rect 9137 5593 9171 5627
rect 9171 5593 9180 5627
rect 9128 5584 9180 5593
rect 14648 5584 14700 5636
rect 15476 5584 15528 5636
rect 16120 5584 16172 5636
rect 11980 5516 12032 5568
rect 14556 5516 14608 5568
rect 14740 5516 14792 5568
rect 16948 5516 17000 5568
rect 5502 5414 5554 5466
rect 5566 5414 5618 5466
rect 5630 5414 5682 5466
rect 5694 5414 5746 5466
rect 5758 5414 5810 5466
rect 5822 5414 5874 5466
rect 5886 5414 5938 5466
rect 5950 5414 6002 5466
rect 6014 5414 6066 5466
rect 6078 5414 6130 5466
rect 6142 5414 6194 5466
rect 6206 5414 6258 5466
rect 6270 5414 6322 5466
rect 6334 5414 6386 5466
rect 6398 5414 6450 5466
rect 6462 5414 6514 5466
rect 6526 5414 6578 5466
rect 6590 5414 6642 5466
rect 6654 5414 6706 5466
rect 13502 5414 13554 5466
rect 13566 5414 13618 5466
rect 13630 5414 13682 5466
rect 13694 5414 13746 5466
rect 13758 5414 13810 5466
rect 13822 5414 13874 5466
rect 13886 5414 13938 5466
rect 13950 5414 14002 5466
rect 14014 5414 14066 5466
rect 14078 5414 14130 5466
rect 14142 5414 14194 5466
rect 14206 5414 14258 5466
rect 14270 5414 14322 5466
rect 14334 5414 14386 5466
rect 14398 5414 14450 5466
rect 14462 5414 14514 5466
rect 14526 5414 14578 5466
rect 14590 5414 14642 5466
rect 14654 5414 14706 5466
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 4344 5312 4396 5364
rect 5724 5355 5776 5364
rect 5724 5321 5733 5355
rect 5733 5321 5767 5355
rect 5767 5321 5776 5355
rect 5724 5312 5776 5321
rect 7380 5312 7432 5364
rect 7564 5312 7616 5364
rect 8024 5312 8076 5364
rect 12072 5312 12124 5364
rect 3056 5287 3108 5296
rect 3056 5253 3065 5287
rect 3065 5253 3099 5287
rect 3099 5253 3108 5287
rect 3056 5244 3108 5253
rect 8116 5244 8168 5296
rect 9128 5244 9180 5296
rect 11980 5287 12032 5296
rect 11980 5253 11989 5287
rect 11989 5253 12023 5287
rect 12023 5253 12032 5287
rect 11980 5244 12032 5253
rect 12256 5244 12308 5296
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 3608 5176 3660 5228
rect 4896 5176 4948 5228
rect 6460 5176 6512 5228
rect 6920 5176 6972 5228
rect 7288 5176 7340 5228
rect 2780 5108 2832 5160
rect 6736 5108 6788 5160
rect 7564 5108 7616 5160
rect 8024 5176 8076 5228
rect 14556 5312 14608 5364
rect 15844 5312 15896 5364
rect 16672 5312 16724 5364
rect 17224 5312 17276 5364
rect 19708 5312 19760 5364
rect 17868 5287 17920 5296
rect 17868 5253 17877 5287
rect 17877 5253 17911 5287
rect 17911 5253 17920 5287
rect 17868 5244 17920 5253
rect 16488 5176 16540 5228
rect 17040 5176 17092 5228
rect 11612 5108 11664 5160
rect 12072 5108 12124 5160
rect 12992 5108 13044 5160
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 15476 5108 15528 5160
rect 17316 5108 17368 5160
rect 18052 5108 18104 5160
rect 6552 5040 6604 5092
rect 16580 5040 16632 5092
rect 6736 4972 6788 5024
rect 8484 4972 8536 5024
rect 14832 4972 14884 5024
rect 15292 4972 15344 5024
rect 17224 4972 17276 5024
rect 17868 4972 17920 5024
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 1502 4870 1554 4922
rect 1566 4870 1618 4922
rect 1630 4870 1682 4922
rect 1694 4870 1746 4922
rect 1758 4870 1810 4922
rect 1822 4870 1874 4922
rect 1886 4870 1938 4922
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 2270 4870 2322 4922
rect 2334 4870 2386 4922
rect 2398 4870 2450 4922
rect 2462 4870 2514 4922
rect 2526 4870 2578 4922
rect 2590 4870 2642 4922
rect 2654 4870 2706 4922
rect 9502 4870 9554 4922
rect 9566 4870 9618 4922
rect 9630 4870 9682 4922
rect 9694 4870 9746 4922
rect 9758 4870 9810 4922
rect 9822 4870 9874 4922
rect 9886 4870 9938 4922
rect 9950 4870 10002 4922
rect 10014 4870 10066 4922
rect 10078 4870 10130 4922
rect 10142 4870 10194 4922
rect 10206 4870 10258 4922
rect 10270 4870 10322 4922
rect 10334 4870 10386 4922
rect 10398 4870 10450 4922
rect 10462 4870 10514 4922
rect 10526 4870 10578 4922
rect 10590 4870 10642 4922
rect 10654 4870 10706 4922
rect 17502 4870 17554 4922
rect 17566 4870 17618 4922
rect 17630 4870 17682 4922
rect 17694 4870 17746 4922
rect 17758 4870 17810 4922
rect 17822 4870 17874 4922
rect 17886 4870 17938 4922
rect 17950 4870 18002 4922
rect 18014 4870 18066 4922
rect 18078 4870 18130 4922
rect 18142 4870 18194 4922
rect 18206 4870 18258 4922
rect 18270 4870 18322 4922
rect 18334 4870 18386 4922
rect 18398 4870 18450 4922
rect 18462 4870 18514 4922
rect 18526 4870 18578 4922
rect 18590 4870 18642 4922
rect 18654 4870 18706 4922
rect 8024 4768 8076 4820
rect 14648 4768 14700 4820
rect 5264 4700 5316 4752
rect 6920 4700 6972 4752
rect 1216 4632 1268 4684
rect 3056 4632 3108 4684
rect 3976 4632 4028 4684
rect 3148 4564 3200 4616
rect 6736 4632 6788 4684
rect 8208 4632 8260 4684
rect 13360 4743 13412 4752
rect 13360 4709 13369 4743
rect 13369 4709 13403 4743
rect 13403 4709 13412 4743
rect 13360 4700 13412 4709
rect 14280 4743 14332 4752
rect 14280 4709 14289 4743
rect 14289 4709 14323 4743
rect 14323 4709 14332 4743
rect 14280 4700 14332 4709
rect 13084 4632 13136 4684
rect 16304 4768 16356 4820
rect 16856 4768 16908 4820
rect 17408 4700 17460 4752
rect 2688 4539 2740 4548
rect 2688 4505 2697 4539
rect 2697 4505 2731 4539
rect 2731 4505 2740 4539
rect 2688 4496 2740 4505
rect 2780 4539 2832 4548
rect 2780 4505 2789 4539
rect 2789 4505 2823 4539
rect 2823 4505 2832 4539
rect 2780 4496 2832 4505
rect 2320 4428 2372 4480
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 8116 4496 8168 4548
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 5080 4428 5132 4480
rect 5724 4428 5776 4480
rect 10692 4496 10744 4548
rect 14556 4607 14608 4616
rect 14556 4573 14564 4607
rect 14564 4573 14598 4607
rect 14598 4573 14608 4607
rect 14556 4564 14608 4573
rect 15292 4632 15344 4684
rect 15384 4675 15436 4684
rect 15384 4641 15393 4675
rect 15393 4641 15427 4675
rect 15427 4641 15436 4675
rect 15384 4632 15436 4641
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 16672 4632 16724 4684
rect 15108 4564 15160 4616
rect 16764 4564 16816 4616
rect 11888 4428 11940 4480
rect 12348 4428 12400 4480
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 15568 4496 15620 4548
rect 16580 4428 16632 4480
rect 18788 4496 18840 4548
rect 19432 4428 19484 4480
rect 5502 4326 5554 4378
rect 5566 4326 5618 4378
rect 5630 4326 5682 4378
rect 5694 4326 5746 4378
rect 5758 4326 5810 4378
rect 5822 4326 5874 4378
rect 5886 4326 5938 4378
rect 5950 4326 6002 4378
rect 6014 4326 6066 4378
rect 6078 4326 6130 4378
rect 6142 4326 6194 4378
rect 6206 4326 6258 4378
rect 6270 4326 6322 4378
rect 6334 4326 6386 4378
rect 6398 4326 6450 4378
rect 6462 4326 6514 4378
rect 6526 4326 6578 4378
rect 6590 4326 6642 4378
rect 6654 4326 6706 4378
rect 13502 4326 13554 4378
rect 13566 4326 13618 4378
rect 13630 4326 13682 4378
rect 13694 4326 13746 4378
rect 13758 4326 13810 4378
rect 13822 4326 13874 4378
rect 13886 4326 13938 4378
rect 13950 4326 14002 4378
rect 14014 4326 14066 4378
rect 14078 4326 14130 4378
rect 14142 4326 14194 4378
rect 14206 4326 14258 4378
rect 14270 4326 14322 4378
rect 14334 4326 14386 4378
rect 14398 4326 14450 4378
rect 14462 4326 14514 4378
rect 14526 4326 14578 4378
rect 14590 4326 14642 4378
rect 14654 4326 14706 4378
rect 2688 4224 2740 4276
rect 6828 4224 6880 4276
rect 7932 4224 7984 4276
rect 11152 4224 11204 4276
rect 14740 4224 14792 4276
rect 3056 4199 3108 4208
rect 3056 4165 3065 4199
rect 3065 4165 3099 4199
rect 3099 4165 3108 4199
rect 3056 4156 3108 4165
rect 5724 4156 5776 4208
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2780 4088 2832 4140
rect 3148 4088 3200 4140
rect 6644 4156 6696 4208
rect 8116 4156 8168 4208
rect 8208 4199 8260 4208
rect 8208 4165 8217 4199
rect 8217 4165 8251 4199
rect 8251 4165 8260 4199
rect 8208 4156 8260 4165
rect 12440 4156 12492 4208
rect 6736 4088 6788 4140
rect 7288 4088 7340 4140
rect 4988 4020 5040 4072
rect 1400 3884 1452 3936
rect 7288 3952 7340 4004
rect 6092 3884 6144 3936
rect 8852 3884 8904 3936
rect 11520 4088 11572 4140
rect 11796 4088 11848 4140
rect 12072 4088 12124 4140
rect 12256 4063 12308 4072
rect 12256 4029 12265 4063
rect 12265 4029 12299 4063
rect 12299 4029 12308 4063
rect 12256 4020 12308 4029
rect 13360 4088 13412 4140
rect 14832 4156 14884 4208
rect 15016 4156 15068 4208
rect 17040 4156 17092 4208
rect 17224 4156 17276 4208
rect 13176 4020 13228 4072
rect 13268 4063 13320 4072
rect 13268 4029 13277 4063
rect 13277 4029 13311 4063
rect 13311 4029 13320 4063
rect 13268 4020 13320 4029
rect 16856 4088 16908 4140
rect 17316 4131 17368 4140
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 18880 4088 18932 4140
rect 15016 4020 15068 4072
rect 15200 4020 15252 4072
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 11888 3952 11940 4004
rect 16948 3952 17000 4004
rect 17132 3952 17184 4004
rect 18880 3952 18932 4004
rect 11336 3884 11388 3936
rect 14740 3884 14792 3936
rect 15016 3884 15068 3936
rect 17316 3884 17368 3936
rect 1502 3782 1554 3834
rect 1566 3782 1618 3834
rect 1630 3782 1682 3834
rect 1694 3782 1746 3834
rect 1758 3782 1810 3834
rect 1822 3782 1874 3834
rect 1886 3782 1938 3834
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 2270 3782 2322 3834
rect 2334 3782 2386 3834
rect 2398 3782 2450 3834
rect 2462 3782 2514 3834
rect 2526 3782 2578 3834
rect 2590 3782 2642 3834
rect 2654 3782 2706 3834
rect 9502 3782 9554 3834
rect 9566 3782 9618 3834
rect 9630 3782 9682 3834
rect 9694 3782 9746 3834
rect 9758 3782 9810 3834
rect 9822 3782 9874 3834
rect 9886 3782 9938 3834
rect 9950 3782 10002 3834
rect 10014 3782 10066 3834
rect 10078 3782 10130 3834
rect 10142 3782 10194 3834
rect 10206 3782 10258 3834
rect 10270 3782 10322 3834
rect 10334 3782 10386 3834
rect 10398 3782 10450 3834
rect 10462 3782 10514 3834
rect 10526 3782 10578 3834
rect 10590 3782 10642 3834
rect 10654 3782 10706 3834
rect 17502 3782 17554 3834
rect 17566 3782 17618 3834
rect 17630 3782 17682 3834
rect 17694 3782 17746 3834
rect 17758 3782 17810 3834
rect 17822 3782 17874 3834
rect 17886 3782 17938 3834
rect 17950 3782 18002 3834
rect 18014 3782 18066 3834
rect 18078 3782 18130 3834
rect 18142 3782 18194 3834
rect 18206 3782 18258 3834
rect 18270 3782 18322 3834
rect 18334 3782 18386 3834
rect 18398 3782 18450 3834
rect 18462 3782 18514 3834
rect 18526 3782 18578 3834
rect 18590 3782 18642 3834
rect 18654 3782 18706 3834
rect 3976 3680 4028 3732
rect 6092 3680 6144 3732
rect 6828 3680 6880 3732
rect 8760 3680 8812 3732
rect 9404 3680 9456 3732
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 11980 3680 12032 3732
rect 13176 3680 13228 3732
rect 204 3612 256 3664
rect 940 3612 992 3664
rect 1400 3612 1452 3664
rect 2780 3655 2832 3664
rect 2780 3621 2789 3655
rect 2789 3621 2823 3655
rect 2823 3621 2832 3655
rect 2780 3612 2832 3621
rect 4804 3612 4856 3664
rect 8484 3612 8536 3664
rect 9220 3655 9272 3664
rect 9220 3621 9229 3655
rect 9229 3621 9263 3655
rect 9263 3621 9272 3655
rect 9220 3612 9272 3621
rect 10416 3612 10468 3664
rect 10508 3612 10560 3664
rect 296 3544 348 3596
rect 2872 3476 2924 3528
rect 2412 3408 2464 3460
rect 2688 3451 2740 3460
rect 2688 3417 2697 3451
rect 2697 3417 2731 3451
rect 2731 3417 2740 3451
rect 2688 3408 2740 3417
rect 3332 3476 3384 3528
rect 4712 3544 4764 3596
rect 3976 3476 4028 3528
rect 4160 3476 4212 3528
rect 7012 3544 7064 3596
rect 11612 3544 11664 3596
rect 13360 3612 13412 3664
rect 14648 3612 14700 3664
rect 15108 3612 15160 3664
rect 17040 3544 17092 3596
rect 17316 3544 17368 3596
rect 1584 3340 1636 3392
rect 5356 3408 5408 3460
rect 8576 3476 8628 3528
rect 5264 3340 5316 3392
rect 7748 3408 7800 3460
rect 7840 3408 7892 3460
rect 9404 3476 9456 3528
rect 10508 3476 10560 3528
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 11244 3476 11296 3528
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 12072 3408 12124 3460
rect 12164 3451 12216 3460
rect 12164 3417 12173 3451
rect 12173 3417 12207 3451
rect 12207 3417 12216 3451
rect 12164 3408 12216 3417
rect 14188 3408 14240 3460
rect 14280 3451 14332 3460
rect 14280 3417 14289 3451
rect 14289 3417 14323 3451
rect 14323 3417 14332 3451
rect 14280 3408 14332 3417
rect 9128 3340 9180 3392
rect 10508 3340 10560 3392
rect 11428 3340 11480 3392
rect 11980 3340 12032 3392
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 16948 3476 17000 3528
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 15568 3408 15620 3460
rect 15752 3408 15804 3460
rect 19524 3408 19576 3460
rect 17224 3340 17276 3392
rect 5502 3238 5554 3290
rect 5566 3238 5618 3290
rect 5630 3238 5682 3290
rect 5694 3238 5746 3290
rect 5758 3238 5810 3290
rect 5822 3238 5874 3290
rect 5886 3238 5938 3290
rect 5950 3238 6002 3290
rect 6014 3238 6066 3290
rect 6078 3238 6130 3290
rect 6142 3238 6194 3290
rect 6206 3238 6258 3290
rect 6270 3238 6322 3290
rect 6334 3238 6386 3290
rect 6398 3238 6450 3290
rect 6462 3238 6514 3290
rect 6526 3238 6578 3290
rect 6590 3238 6642 3290
rect 6654 3238 6706 3290
rect 13502 3238 13554 3290
rect 13566 3238 13618 3290
rect 13630 3238 13682 3290
rect 13694 3238 13746 3290
rect 13758 3238 13810 3290
rect 13822 3238 13874 3290
rect 13886 3238 13938 3290
rect 13950 3238 14002 3290
rect 14014 3238 14066 3290
rect 14078 3238 14130 3290
rect 14142 3238 14194 3290
rect 14206 3238 14258 3290
rect 14270 3238 14322 3290
rect 14334 3238 14386 3290
rect 14398 3238 14450 3290
rect 14462 3238 14514 3290
rect 14526 3238 14578 3290
rect 14590 3238 14642 3290
rect 14654 3238 14706 3290
rect 2688 3136 2740 3188
rect 5540 3136 5592 3188
rect 6828 3136 6880 3188
rect 7656 3136 7708 3188
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 8392 3179 8444 3188
rect 8392 3145 8401 3179
rect 8401 3145 8435 3179
rect 8435 3145 8444 3179
rect 8392 3136 8444 3145
rect 9220 3136 9272 3188
rect 2412 3111 2464 3120
rect 2412 3077 2421 3111
rect 2421 3077 2455 3111
rect 2455 3077 2464 3111
rect 2412 3068 2464 3077
rect 5356 3068 5408 3120
rect 8668 3068 8720 3120
rect 9588 3111 9640 3120
rect 9588 3077 9597 3111
rect 9597 3077 9631 3111
rect 9631 3077 9640 3111
rect 9588 3068 9640 3077
rect 12164 3136 12216 3188
rect 13360 3136 13412 3188
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 1124 2932 1176 2984
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 7104 3000 7156 3052
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 9312 3000 9364 3052
rect 10784 3000 10836 3052
rect 2872 2975 2924 2984
rect 2872 2941 2881 2975
rect 2881 2941 2915 2975
rect 2915 2941 2924 2975
rect 2872 2932 2924 2941
rect 6644 2975 6696 2984
rect 6644 2941 6653 2975
rect 6653 2941 6687 2975
rect 6687 2941 6696 2975
rect 6644 2932 6696 2941
rect 8944 2932 8996 2984
rect 4620 2864 4672 2916
rect 6828 2864 6880 2916
rect 9036 2864 9088 2916
rect 11888 2932 11940 2984
rect 10508 2864 10560 2916
rect 10784 2864 10836 2916
rect 10876 2864 10928 2916
rect 11244 2864 11296 2916
rect 12072 3000 12124 3052
rect 13268 3000 13320 3052
rect 13912 3000 13964 3052
rect 12348 2932 12400 2984
rect 12716 2975 12768 2984
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 12716 2932 12768 2941
rect 13084 2932 13136 2984
rect 15384 3136 15436 3188
rect 15568 3136 15620 3188
rect 16856 3136 16908 3188
rect 17040 3136 17092 3188
rect 19616 3136 19668 3188
rect 14740 3111 14792 3120
rect 14740 3077 14749 3111
rect 14749 3077 14783 3111
rect 14783 3077 14792 3111
rect 14740 3068 14792 3077
rect 16396 3068 16448 3120
rect 16028 3000 16080 3052
rect 12900 2864 12952 2916
rect 17040 2975 17092 2984
rect 17040 2941 17049 2975
rect 17049 2941 17083 2975
rect 17083 2941 17092 2975
rect 17040 2932 17092 2941
rect 17224 3000 17276 3052
rect 17132 2864 17184 2916
rect 9128 2796 9180 2848
rect 10692 2796 10744 2848
rect 15200 2796 15252 2848
rect 19892 3000 19944 3052
rect 1502 2694 1554 2746
rect 1566 2694 1618 2746
rect 1630 2694 1682 2746
rect 1694 2694 1746 2746
rect 1758 2694 1810 2746
rect 1822 2694 1874 2746
rect 1886 2694 1938 2746
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 2270 2694 2322 2746
rect 2334 2694 2386 2746
rect 2398 2694 2450 2746
rect 2462 2694 2514 2746
rect 2526 2694 2578 2746
rect 2590 2694 2642 2746
rect 2654 2694 2706 2746
rect 9502 2694 9554 2746
rect 9566 2694 9618 2746
rect 9630 2694 9682 2746
rect 9694 2694 9746 2746
rect 9758 2694 9810 2746
rect 9822 2694 9874 2746
rect 9886 2694 9938 2746
rect 9950 2694 10002 2746
rect 10014 2694 10066 2746
rect 10078 2694 10130 2746
rect 10142 2694 10194 2746
rect 10206 2694 10258 2746
rect 10270 2694 10322 2746
rect 10334 2694 10386 2746
rect 10398 2694 10450 2746
rect 10462 2694 10514 2746
rect 10526 2694 10578 2746
rect 10590 2694 10642 2746
rect 10654 2694 10706 2746
rect 17502 2694 17554 2746
rect 17566 2694 17618 2746
rect 17630 2694 17682 2746
rect 17694 2694 17746 2746
rect 17758 2694 17810 2746
rect 17822 2694 17874 2746
rect 17886 2694 17938 2746
rect 17950 2694 18002 2746
rect 18014 2694 18066 2746
rect 18078 2694 18130 2746
rect 18142 2694 18194 2746
rect 18206 2694 18258 2746
rect 18270 2694 18322 2746
rect 18334 2694 18386 2746
rect 18398 2694 18450 2746
rect 18462 2694 18514 2746
rect 18526 2694 18578 2746
rect 18590 2694 18642 2746
rect 18654 2694 18706 2746
rect 1400 2592 1452 2644
rect 4160 2592 4212 2644
rect 6828 2592 6880 2644
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 7840 2592 7892 2644
rect 8576 2592 8628 2644
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 13912 2592 13964 2644
rect 15016 2592 15068 2644
rect 19248 2592 19300 2644
rect 940 2524 992 2576
rect 5080 2524 5132 2576
rect 4436 2456 4488 2508
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 4160 2320 4212 2372
rect 8392 2456 8444 2508
rect 9036 2456 9088 2508
rect 5172 2252 5224 2304
rect 7564 2295 7616 2304
rect 7564 2261 7573 2295
rect 7573 2261 7607 2295
rect 7607 2261 7616 2295
rect 7564 2252 7616 2261
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9312 2499 9364 2508
rect 9312 2465 9321 2499
rect 9321 2465 9355 2499
rect 9355 2465 9364 2499
rect 9312 2456 9364 2465
rect 9772 2456 9824 2508
rect 9680 2388 9732 2440
rect 9220 2320 9272 2372
rect 11060 2456 11112 2508
rect 11796 2456 11848 2508
rect 13084 2499 13136 2508
rect 13084 2465 13093 2499
rect 13093 2465 13127 2499
rect 13127 2465 13136 2499
rect 13084 2456 13136 2465
rect 15016 2456 15068 2508
rect 15384 2456 15436 2508
rect 16672 2456 16724 2508
rect 10876 2388 10928 2440
rect 11520 2388 11572 2440
rect 12256 2388 12308 2440
rect 10600 2363 10652 2372
rect 10600 2329 10609 2363
rect 10609 2329 10643 2363
rect 10643 2329 10652 2363
rect 10600 2320 10652 2329
rect 11244 2320 11296 2372
rect 10784 2252 10836 2304
rect 12256 2295 12308 2304
rect 12256 2261 12265 2295
rect 12265 2261 12299 2295
rect 12299 2261 12308 2295
rect 12256 2252 12308 2261
rect 12440 2388 12492 2440
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 14924 2388 14976 2440
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 17132 2456 17184 2508
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 19708 2388 19760 2440
rect 17040 2295 17092 2304
rect 17040 2261 17049 2295
rect 17049 2261 17083 2295
rect 17083 2261 17092 2295
rect 17040 2252 17092 2261
rect 17316 2252 17368 2304
rect 5502 2150 5554 2202
rect 5566 2150 5618 2202
rect 5630 2150 5682 2202
rect 5694 2150 5746 2202
rect 5758 2150 5810 2202
rect 5822 2150 5874 2202
rect 5886 2150 5938 2202
rect 5950 2150 6002 2202
rect 6014 2150 6066 2202
rect 6078 2150 6130 2202
rect 6142 2150 6194 2202
rect 6206 2150 6258 2202
rect 6270 2150 6322 2202
rect 6334 2150 6386 2202
rect 6398 2150 6450 2202
rect 6462 2150 6514 2202
rect 6526 2150 6578 2202
rect 6590 2150 6642 2202
rect 6654 2150 6706 2202
rect 13502 2150 13554 2202
rect 13566 2150 13618 2202
rect 13630 2150 13682 2202
rect 13694 2150 13746 2202
rect 13758 2150 13810 2202
rect 13822 2150 13874 2202
rect 13886 2150 13938 2202
rect 13950 2150 14002 2202
rect 14014 2150 14066 2202
rect 14078 2150 14130 2202
rect 14142 2150 14194 2202
rect 14206 2150 14258 2202
rect 14270 2150 14322 2202
rect 14334 2150 14386 2202
rect 14398 2150 14450 2202
rect 14462 2150 14514 2202
rect 14526 2150 14578 2202
rect 14590 2150 14642 2202
rect 14654 2150 14706 2202
rect 3516 2048 3568 2100
rect 9680 2048 9732 2100
rect 11152 2048 11204 2100
rect 12256 2048 12308 2100
rect 14832 2048 14884 2100
rect 15016 2048 15068 2100
rect 17040 2048 17092 2100
rect 7932 1980 7984 2032
rect 15844 1980 15896 2032
rect 8116 1912 8168 1964
rect 17868 1844 17920 1896
rect 3424 1776 3476 1828
rect 10600 1776 10652 1828
rect 9128 1708 9180 1760
rect 19340 1708 19392 1760
rect 7564 1640 7616 1692
rect 18788 1640 18840 1692
rect 3424 1300 3476 1352
rect 10968 1300 11020 1352
rect 4068 1232 4120 1284
rect 15384 1232 15436 1284
rect 3332 1164 3384 1216
rect 9588 1164 9640 1216
rect 3516 1028 3568 1080
rect 8852 1028 8904 1080
rect 296 960 348 1012
rect 5264 960 5316 1012
<< metal2 >>
rect 110 19200 166 20000
rect 294 19200 350 20000
rect 478 19200 534 20000
rect 662 19200 718 20000
rect 846 19200 902 20000
rect 1030 19200 1086 20000
rect 1214 19200 1270 20000
rect 1398 19200 1454 20000
rect 1582 19200 1638 20000
rect 1766 19200 1822 20000
rect 1950 19200 2006 20000
rect 2134 19200 2190 20000
rect 2318 19200 2374 20000
rect 20 17196 72 17202
rect 20 17138 72 17144
rect 32 13054 60 17138
rect 20 13048 72 13054
rect 20 12990 72 12996
rect 124 12918 152 19200
rect 308 15570 336 19200
rect 388 16108 440 16114
rect 388 16050 440 16056
rect 296 15564 348 15570
rect 296 15506 348 15512
rect 204 15428 256 15434
rect 204 15370 256 15376
rect 20 12912 72 12918
rect 20 12854 72 12860
rect 112 12912 164 12918
rect 112 12854 164 12860
rect 32 10169 60 12854
rect 110 12744 166 12753
rect 110 12679 166 12688
rect 18 10160 74 10169
rect 18 10095 74 10104
rect 124 9722 152 12679
rect 112 9716 164 9722
rect 112 9658 164 9664
rect 216 3670 244 15370
rect 296 15292 348 15298
rect 296 15234 348 15240
rect 308 10742 336 15234
rect 296 10736 348 10742
rect 296 10678 348 10684
rect 296 9852 348 9858
rect 296 9794 348 9800
rect 204 3664 256 3670
rect 204 3606 256 3612
rect 308 3602 336 9794
rect 400 8090 428 16050
rect 492 16046 520 19200
rect 572 17264 624 17270
rect 572 17206 624 17212
rect 480 16040 532 16046
rect 480 15982 532 15988
rect 480 15496 532 15502
rect 480 15438 532 15444
rect 492 13190 520 15438
rect 584 14385 612 17206
rect 676 15502 704 19200
rect 756 17128 808 17134
rect 756 17070 808 17076
rect 664 15496 716 15502
rect 664 15438 716 15444
rect 664 15360 716 15366
rect 664 15302 716 15308
rect 570 14376 626 14385
rect 570 14311 626 14320
rect 584 14006 612 14311
rect 572 14000 624 14006
rect 572 13942 624 13948
rect 572 13864 624 13870
rect 572 13806 624 13812
rect 480 13184 532 13190
rect 480 13126 532 13132
rect 480 13048 532 13054
rect 480 12990 532 12996
rect 388 8084 440 8090
rect 388 8026 440 8032
rect 296 3596 348 3602
rect 296 3538 348 3544
rect 492 2774 520 12990
rect 584 9518 612 13806
rect 676 13530 704 15302
rect 768 15298 796 17070
rect 756 15292 808 15298
rect 756 15234 808 15240
rect 756 14952 808 14958
rect 756 14894 808 14900
rect 768 14521 796 14894
rect 754 14512 810 14521
rect 754 14447 810 14456
rect 756 14340 808 14346
rect 756 14282 808 14288
rect 664 13524 716 13530
rect 664 13466 716 13472
rect 662 13152 718 13161
rect 662 13087 718 13096
rect 572 9512 624 9518
rect 572 9454 624 9460
rect 676 4593 704 13087
rect 768 11234 796 14282
rect 860 12306 888 19200
rect 940 16584 992 16590
rect 940 16526 992 16532
rect 848 12300 900 12306
rect 848 12242 900 12248
rect 768 11206 888 11234
rect 754 11112 810 11121
rect 754 11047 810 11056
rect 662 4584 718 4593
rect 662 4519 718 4528
rect 124 2746 520 2774
rect 768 2774 796 11047
rect 860 9858 888 11206
rect 848 9852 900 9858
rect 848 9794 900 9800
rect 952 9602 980 16526
rect 1044 15366 1072 19200
rect 1228 17218 1256 19200
rect 1136 17190 1256 17218
rect 1032 15360 1084 15366
rect 1032 15302 1084 15308
rect 1032 14816 1084 14822
rect 1032 14758 1084 14764
rect 1044 9994 1072 14758
rect 1136 13938 1164 17190
rect 1216 17060 1268 17066
rect 1216 17002 1268 17008
rect 1228 14414 1256 17002
rect 1308 16992 1360 16998
rect 1308 16934 1360 16940
rect 1320 15094 1348 16934
rect 1308 15088 1360 15094
rect 1308 15030 1360 15036
rect 1308 14884 1360 14890
rect 1308 14826 1360 14832
rect 1216 14408 1268 14414
rect 1216 14350 1268 14356
rect 1216 14068 1268 14074
rect 1216 14010 1268 14016
rect 1124 13932 1176 13938
rect 1124 13874 1176 13880
rect 1228 13818 1256 14010
rect 1320 14006 1348 14826
rect 1308 14000 1360 14006
rect 1308 13942 1360 13948
rect 1136 13790 1256 13818
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 1136 10810 1164 13790
rect 1216 13728 1268 13734
rect 1216 13670 1268 13676
rect 1124 10804 1176 10810
rect 1124 10746 1176 10752
rect 1228 10146 1256 13670
rect 1320 12986 1348 13806
rect 1308 12980 1360 12986
rect 1308 12922 1360 12928
rect 1412 12730 1440 19200
rect 1596 17542 1624 19200
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1780 16998 1808 19200
rect 1964 17066 1992 19200
rect 2148 17218 2176 19200
rect 2332 17338 2360 19200
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 5502 17436 6706 17445
rect 5502 17434 5516 17436
rect 5572 17434 5596 17436
rect 5652 17434 5676 17436
rect 5732 17434 5756 17436
rect 5812 17434 5836 17436
rect 5892 17434 5916 17436
rect 5972 17434 5996 17436
rect 6052 17434 6076 17436
rect 6132 17434 6156 17436
rect 6212 17434 6236 17436
rect 6292 17434 6316 17436
rect 6372 17434 6396 17436
rect 6452 17434 6476 17436
rect 6532 17434 6556 17436
rect 6612 17434 6636 17436
rect 6692 17434 6706 17436
rect 5746 17382 5756 17434
rect 5812 17382 5822 17434
rect 6066 17382 6076 17434
rect 6132 17382 6142 17434
rect 6386 17382 6396 17434
rect 6452 17382 6462 17434
rect 5502 17380 5516 17382
rect 5572 17380 5596 17382
rect 5652 17380 5676 17382
rect 5732 17380 5756 17382
rect 5812 17380 5836 17382
rect 5892 17380 5916 17382
rect 5972 17380 5996 17382
rect 6052 17380 6076 17382
rect 6132 17380 6156 17382
rect 6212 17380 6236 17382
rect 6292 17380 6316 17382
rect 6372 17380 6396 17382
rect 6452 17380 6476 17382
rect 6532 17380 6556 17382
rect 6612 17380 6636 17382
rect 6692 17380 6706 17382
rect 5502 17371 6706 17380
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 2056 17190 2176 17218
rect 3330 17232 3386 17241
rect 2056 17134 2084 17190
rect 3330 17167 3332 17176
rect 3384 17167 3386 17176
rect 4344 17196 4396 17202
rect 3332 17138 3384 17144
rect 4344 17138 4396 17144
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3884 17060 3936 17066
rect 3884 17002 3936 17008
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1502 16892 2706 16901
rect 1502 16890 1516 16892
rect 1572 16890 1596 16892
rect 1652 16890 1676 16892
rect 1732 16890 1756 16892
rect 1812 16890 1836 16892
rect 1892 16890 1916 16892
rect 1972 16890 1996 16892
rect 2052 16890 2076 16892
rect 2132 16890 2156 16892
rect 2212 16890 2236 16892
rect 2292 16890 2316 16892
rect 2372 16890 2396 16892
rect 2452 16890 2476 16892
rect 2532 16890 2556 16892
rect 2612 16890 2636 16892
rect 2692 16890 2706 16892
rect 1746 16838 1756 16890
rect 1812 16838 1822 16890
rect 2066 16838 2076 16890
rect 2132 16838 2142 16890
rect 2386 16838 2396 16890
rect 2452 16838 2462 16890
rect 1502 16836 1516 16838
rect 1572 16836 1596 16838
rect 1652 16836 1676 16838
rect 1732 16836 1756 16838
rect 1812 16836 1836 16838
rect 1892 16836 1916 16838
rect 1972 16836 1996 16838
rect 2052 16836 2076 16838
rect 2132 16836 2156 16838
rect 2212 16836 2236 16838
rect 2292 16836 2316 16838
rect 2372 16836 2396 16838
rect 2452 16836 2476 16838
rect 2532 16836 2556 16838
rect 2612 16836 2636 16838
rect 2692 16836 2706 16838
rect 1502 16827 2706 16836
rect 2780 16584 2832 16590
rect 2832 16544 2912 16572
rect 2780 16526 2832 16532
rect 1952 16516 2004 16522
rect 1952 16458 2004 16464
rect 1964 15978 1992 16458
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 16182 2544 16390
rect 2504 16176 2556 16182
rect 2504 16118 2556 16124
rect 2700 15978 2820 15994
rect 1952 15972 2004 15978
rect 1952 15914 2004 15920
rect 2688 15972 2820 15978
rect 2740 15966 2820 15972
rect 2688 15914 2740 15920
rect 1502 15804 2706 15813
rect 1502 15802 1516 15804
rect 1572 15802 1596 15804
rect 1652 15802 1676 15804
rect 1732 15802 1756 15804
rect 1812 15802 1836 15804
rect 1892 15802 1916 15804
rect 1972 15802 1996 15804
rect 2052 15802 2076 15804
rect 2132 15802 2156 15804
rect 2212 15802 2236 15804
rect 2292 15802 2316 15804
rect 2372 15802 2396 15804
rect 2452 15802 2476 15804
rect 2532 15802 2556 15804
rect 2612 15802 2636 15804
rect 2692 15802 2706 15804
rect 1746 15750 1756 15802
rect 1812 15750 1822 15802
rect 2066 15750 2076 15802
rect 2132 15750 2142 15802
rect 2386 15750 2396 15802
rect 2452 15750 2462 15802
rect 1502 15748 1516 15750
rect 1572 15748 1596 15750
rect 1652 15748 1676 15750
rect 1732 15748 1756 15750
rect 1812 15748 1836 15750
rect 1892 15748 1916 15750
rect 1972 15748 1996 15750
rect 2052 15748 2076 15750
rect 2132 15748 2156 15750
rect 2212 15748 2236 15750
rect 2292 15748 2316 15750
rect 2372 15748 2396 15750
rect 2452 15748 2476 15750
rect 2532 15748 2556 15750
rect 2612 15748 2636 15750
rect 2692 15748 2706 15750
rect 1502 15739 2706 15748
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 1584 15632 1636 15638
rect 1584 15574 1636 15580
rect 1596 14958 1624 15574
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1872 15162 1900 15302
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1964 14890 1992 15438
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 2608 14804 2636 15642
rect 2792 15586 2820 15966
rect 2884 15706 2912 16544
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2976 15586 3004 16390
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 2700 15558 2820 15586
rect 2884 15558 3004 15586
rect 2700 15502 2728 15558
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2884 15178 2912 15558
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2792 15150 2912 15178
rect 2792 14929 2820 15150
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 2778 14920 2834 14929
rect 2778 14855 2834 14864
rect 2608 14776 2820 14804
rect 1502 14716 2706 14725
rect 1502 14714 1516 14716
rect 1572 14714 1596 14716
rect 1652 14714 1676 14716
rect 1732 14714 1756 14716
rect 1812 14714 1836 14716
rect 1892 14714 1916 14716
rect 1972 14714 1996 14716
rect 2052 14714 2076 14716
rect 2132 14714 2156 14716
rect 2212 14714 2236 14716
rect 2292 14714 2316 14716
rect 2372 14714 2396 14716
rect 2452 14714 2476 14716
rect 2532 14714 2556 14716
rect 2612 14714 2636 14716
rect 2692 14714 2706 14716
rect 1746 14662 1756 14714
rect 1812 14662 1822 14714
rect 2066 14662 2076 14714
rect 2132 14662 2142 14714
rect 2386 14662 2396 14714
rect 2452 14662 2462 14714
rect 1502 14660 1516 14662
rect 1572 14660 1596 14662
rect 1652 14660 1676 14662
rect 1732 14660 1756 14662
rect 1812 14660 1836 14662
rect 1892 14660 1916 14662
rect 1972 14660 1996 14662
rect 2052 14660 2076 14662
rect 2132 14660 2156 14662
rect 2212 14660 2236 14662
rect 2292 14660 2316 14662
rect 2372 14660 2396 14662
rect 2452 14660 2476 14662
rect 2532 14660 2556 14662
rect 2612 14660 2636 14662
rect 2692 14660 2706 14662
rect 1502 14651 2706 14660
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 1582 14512 1638 14521
rect 1582 14447 1638 14456
rect 1596 13870 1624 14447
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 2056 13938 2084 14214
rect 2148 14006 2176 14554
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1584 13864 1636 13870
rect 2240 13841 2268 14350
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 13870 2728 14214
rect 2688 13864 2740 13870
rect 1584 13806 1636 13812
rect 1858 13832 1914 13841
rect 1858 13767 1914 13776
rect 2226 13832 2282 13841
rect 2688 13806 2740 13812
rect 2226 13767 2282 13776
rect 1872 13734 1900 13767
rect 1860 13728 1912 13734
rect 1860 13670 1912 13676
rect 1502 13628 2706 13637
rect 1502 13626 1516 13628
rect 1572 13626 1596 13628
rect 1652 13626 1676 13628
rect 1732 13626 1756 13628
rect 1812 13626 1836 13628
rect 1892 13626 1916 13628
rect 1972 13626 1996 13628
rect 2052 13626 2076 13628
rect 2132 13626 2156 13628
rect 2212 13626 2236 13628
rect 2292 13626 2316 13628
rect 2372 13626 2396 13628
rect 2452 13626 2476 13628
rect 2532 13626 2556 13628
rect 2612 13626 2636 13628
rect 2692 13626 2706 13628
rect 1746 13574 1756 13626
rect 1812 13574 1822 13626
rect 2066 13574 2076 13626
rect 2132 13574 2142 13626
rect 2386 13574 2396 13626
rect 2452 13574 2462 13626
rect 1502 13572 1516 13574
rect 1572 13572 1596 13574
rect 1652 13572 1676 13574
rect 1732 13572 1756 13574
rect 1812 13572 1836 13574
rect 1892 13572 1916 13574
rect 1972 13572 1996 13574
rect 2052 13572 2076 13574
rect 2132 13572 2156 13574
rect 2212 13572 2236 13574
rect 2292 13572 2316 13574
rect 2372 13572 2396 13574
rect 2452 13572 2476 13574
rect 2532 13572 2556 13574
rect 2612 13572 2636 13574
rect 2692 13572 2706 13574
rect 1502 13563 2706 13572
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 1766 13424 1822 13433
rect 1766 13359 1822 13368
rect 1780 13326 1808 13359
rect 1768 13320 1820 13326
rect 1768 13262 1820 13268
rect 1950 13288 2006 13297
rect 1950 13223 1952 13232
rect 2004 13223 2006 13232
rect 1952 13194 2004 13200
rect 2240 12782 2268 13466
rect 2332 13433 2360 13466
rect 2318 13424 2374 13433
rect 2318 13359 2374 13368
rect 2332 12986 2360 13359
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2332 12889 2360 12922
rect 2318 12880 2374 12889
rect 2424 12850 2452 13262
rect 2318 12815 2374 12824
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 1320 12702 1440 12730
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 1320 11778 1348 12702
rect 1492 12640 1544 12646
rect 1412 12600 1492 12628
rect 1412 11898 1440 12600
rect 1492 12582 1544 12588
rect 1860 12640 1912 12646
rect 2332 12628 2360 12718
rect 2516 12696 2544 13262
rect 2596 13252 2648 13258
rect 2792 13240 2820 14776
rect 2884 14006 2912 15030
rect 2976 14958 3004 15438
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2976 13852 3004 14350
rect 3068 14074 3096 16050
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 2884 13824 3004 13852
rect 2884 13462 2912 13824
rect 3056 13728 3108 13734
rect 2962 13696 3018 13705
rect 3056 13670 3108 13676
rect 2962 13631 3018 13640
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2648 13212 2820 13240
rect 2596 13194 2648 13200
rect 2792 12986 2820 13212
rect 2884 13190 2912 13262
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2700 12753 2728 12922
rect 2870 12880 2926 12889
rect 2976 12866 3004 13631
rect 2926 12838 3004 12866
rect 2870 12815 2926 12824
rect 2780 12776 2832 12782
rect 2686 12744 2742 12753
rect 2596 12708 2648 12714
rect 2516 12668 2596 12696
rect 2780 12718 2832 12724
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2686 12679 2742 12688
rect 2596 12650 2648 12656
rect 1912 12600 2360 12628
rect 1860 12582 1912 12588
rect 1502 12540 2706 12549
rect 1502 12538 1516 12540
rect 1572 12538 1596 12540
rect 1652 12538 1676 12540
rect 1732 12538 1756 12540
rect 1812 12538 1836 12540
rect 1892 12538 1916 12540
rect 1972 12538 1996 12540
rect 2052 12538 2076 12540
rect 2132 12538 2156 12540
rect 2212 12538 2236 12540
rect 2292 12538 2316 12540
rect 2372 12538 2396 12540
rect 2452 12538 2476 12540
rect 2532 12538 2556 12540
rect 2612 12538 2636 12540
rect 2692 12538 2706 12540
rect 1746 12486 1756 12538
rect 1812 12486 1822 12538
rect 2066 12486 2076 12538
rect 2132 12486 2142 12538
rect 2386 12486 2396 12538
rect 2452 12486 2462 12538
rect 1502 12484 1516 12486
rect 1572 12484 1596 12486
rect 1652 12484 1676 12486
rect 1732 12484 1756 12486
rect 1812 12484 1836 12486
rect 1892 12484 1916 12486
rect 1972 12484 1996 12486
rect 2052 12484 2076 12486
rect 2132 12484 2156 12486
rect 2212 12484 2236 12486
rect 2292 12484 2316 12486
rect 2372 12484 2396 12486
rect 2452 12484 2476 12486
rect 2532 12484 2556 12486
rect 2612 12484 2636 12486
rect 2692 12484 2706 12486
rect 1502 12475 2706 12484
rect 1768 12436 1820 12442
rect 2792 12424 2820 12718
rect 2884 12442 2912 12718
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 1768 12378 1820 12384
rect 2608 12396 2820 12424
rect 2872 12436 2924 12442
rect 1780 12238 1808 12378
rect 2504 12368 2556 12374
rect 2318 12336 2374 12345
rect 2504 12310 2556 12316
rect 2318 12271 2320 12280
rect 2372 12271 2374 12280
rect 2320 12242 2372 12248
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 2226 12200 2282 12209
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1320 11750 1440 11778
rect 1308 11552 1360 11558
rect 1308 11494 1360 11500
rect 1320 11082 1348 11494
rect 1412 11218 1440 11750
rect 1780 11558 1808 12174
rect 2226 12135 2282 12144
rect 2240 12102 2268 12135
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2424 11665 2452 11766
rect 2410 11656 2466 11665
rect 2516 11642 2544 12310
rect 2608 11830 2636 12396
rect 2872 12378 2924 12384
rect 2870 12336 2926 12345
rect 2870 12271 2926 12280
rect 2884 11830 2912 12271
rect 2596 11824 2648 11830
rect 2594 11792 2596 11801
rect 2872 11824 2924 11830
rect 2648 11792 2650 11801
rect 2872 11766 2924 11772
rect 2594 11727 2650 11736
rect 2516 11614 2820 11642
rect 2410 11591 2466 11600
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1502 11452 2706 11461
rect 1502 11450 1516 11452
rect 1572 11450 1596 11452
rect 1652 11450 1676 11452
rect 1732 11450 1756 11452
rect 1812 11450 1836 11452
rect 1892 11450 1916 11452
rect 1972 11450 1996 11452
rect 2052 11450 2076 11452
rect 2132 11450 2156 11452
rect 2212 11450 2236 11452
rect 2292 11450 2316 11452
rect 2372 11450 2396 11452
rect 2452 11450 2476 11452
rect 2532 11450 2556 11452
rect 2612 11450 2636 11452
rect 2692 11450 2706 11452
rect 1746 11398 1756 11450
rect 1812 11398 1822 11450
rect 2066 11398 2076 11450
rect 2132 11398 2142 11450
rect 2386 11398 2396 11450
rect 2452 11398 2462 11450
rect 1502 11396 1516 11398
rect 1572 11396 1596 11398
rect 1652 11396 1676 11398
rect 1732 11396 1756 11398
rect 1812 11396 1836 11398
rect 1892 11396 1916 11398
rect 1972 11396 1996 11398
rect 2052 11396 2076 11398
rect 2132 11396 2156 11398
rect 2212 11396 2236 11398
rect 2292 11396 2316 11398
rect 2372 11396 2396 11398
rect 2452 11396 2476 11398
rect 2532 11396 2556 11398
rect 2612 11396 2636 11398
rect 2692 11396 2706 11398
rect 1502 11387 2706 11396
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1308 11076 1360 11082
rect 1308 11018 1360 11024
rect 1780 10674 1808 11290
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1872 10538 1900 10911
rect 2240 10742 2268 11018
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 1860 10532 1912 10538
rect 1860 10474 1912 10480
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1228 10118 1348 10146
rect 1032 9988 1084 9994
rect 1032 9930 1084 9936
rect 1216 9920 1268 9926
rect 1216 9862 1268 9868
rect 952 9574 1164 9602
rect 1032 9512 1084 9518
rect 1032 9454 1084 9460
rect 940 8084 992 8090
rect 940 8026 992 8032
rect 952 3777 980 8026
rect 938 3768 994 3777
rect 938 3703 994 3712
rect 940 3664 992 3670
rect 940 3606 992 3612
rect 952 2961 980 3606
rect 1044 3233 1072 9454
rect 1136 3505 1164 9574
rect 1228 4690 1256 9862
rect 1320 8090 1348 10118
rect 1308 8084 1360 8090
rect 1308 8026 1360 8032
rect 1412 7154 1440 10406
rect 1502 10364 2706 10373
rect 1502 10362 1516 10364
rect 1572 10362 1596 10364
rect 1652 10362 1676 10364
rect 1732 10362 1756 10364
rect 1812 10362 1836 10364
rect 1892 10362 1916 10364
rect 1972 10362 1996 10364
rect 2052 10362 2076 10364
rect 2132 10362 2156 10364
rect 2212 10362 2236 10364
rect 2292 10362 2316 10364
rect 2372 10362 2396 10364
rect 2452 10362 2476 10364
rect 2532 10362 2556 10364
rect 2612 10362 2636 10364
rect 2692 10362 2706 10364
rect 1746 10310 1756 10362
rect 1812 10310 1822 10362
rect 2066 10310 2076 10362
rect 2132 10310 2142 10362
rect 2386 10310 2396 10362
rect 2452 10310 2462 10362
rect 1502 10308 1516 10310
rect 1572 10308 1596 10310
rect 1652 10308 1676 10310
rect 1732 10308 1756 10310
rect 1812 10308 1836 10310
rect 1892 10308 1916 10310
rect 1972 10308 1996 10310
rect 2052 10308 2076 10310
rect 2132 10308 2156 10310
rect 2212 10308 2236 10310
rect 2292 10308 2316 10310
rect 2372 10308 2396 10310
rect 2452 10308 2476 10310
rect 2532 10308 2556 10310
rect 2612 10308 2636 10310
rect 2692 10308 2706 10310
rect 1502 10299 2706 10308
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2332 9586 2360 10066
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2424 9586 2452 9930
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2608 9382 2636 10202
rect 2792 10044 2820 11614
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2884 10266 2912 11086
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2872 10056 2924 10062
rect 2792 10016 2872 10044
rect 2872 9998 2924 10004
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2700 9654 2728 9930
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 1502 9276 2706 9285
rect 1502 9274 1516 9276
rect 1572 9274 1596 9276
rect 1652 9274 1676 9276
rect 1732 9274 1756 9276
rect 1812 9274 1836 9276
rect 1892 9274 1916 9276
rect 1972 9274 1996 9276
rect 2052 9274 2076 9276
rect 2132 9274 2156 9276
rect 2212 9274 2236 9276
rect 2292 9274 2316 9276
rect 2372 9274 2396 9276
rect 2452 9274 2476 9276
rect 2532 9274 2556 9276
rect 2612 9274 2636 9276
rect 2692 9274 2706 9276
rect 1746 9222 1756 9274
rect 1812 9222 1822 9274
rect 2066 9222 2076 9274
rect 2132 9222 2142 9274
rect 2386 9222 2396 9274
rect 2452 9222 2462 9274
rect 1502 9220 1516 9222
rect 1572 9220 1596 9222
rect 1652 9220 1676 9222
rect 1732 9220 1756 9222
rect 1812 9220 1836 9222
rect 1892 9220 1916 9222
rect 1972 9220 1996 9222
rect 2052 9220 2076 9222
rect 2132 9220 2156 9222
rect 2212 9220 2236 9222
rect 2292 9220 2316 9222
rect 2372 9220 2396 9222
rect 2452 9220 2476 9222
rect 2532 9220 2556 9222
rect 2612 9220 2636 9222
rect 2692 9220 2706 9222
rect 1502 9211 2706 9220
rect 2792 8906 2820 9454
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2228 8900 2280 8906
rect 2228 8842 2280 8848
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2240 8566 2268 8842
rect 2700 8634 2728 8842
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2884 8498 2912 8978
rect 2976 8974 3004 12582
rect 3068 9110 3096 13670
rect 3160 12628 3188 15846
rect 3252 12782 3280 17002
rect 3608 16516 3660 16522
rect 3608 16458 3660 16464
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3344 15706 3372 15914
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3436 15434 3464 16050
rect 3424 15428 3476 15434
rect 3424 15370 3476 15376
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3160 12600 3280 12628
rect 3146 12472 3202 12481
rect 3146 12407 3202 12416
rect 3160 12238 3188 12407
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3146 12064 3202 12073
rect 3146 11999 3202 12008
rect 3160 11898 3188 11999
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3146 11656 3202 11665
rect 3146 11591 3202 11600
rect 3160 10470 3188 11591
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3160 10266 3188 10406
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3160 9518 3188 9998
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 3068 8974 3096 9046
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 1502 8188 2706 8197
rect 1502 8186 1516 8188
rect 1572 8186 1596 8188
rect 1652 8186 1676 8188
rect 1732 8186 1756 8188
rect 1812 8186 1836 8188
rect 1892 8186 1916 8188
rect 1972 8186 1996 8188
rect 2052 8186 2076 8188
rect 2132 8186 2156 8188
rect 2212 8186 2236 8188
rect 2292 8186 2316 8188
rect 2372 8186 2396 8188
rect 2452 8186 2476 8188
rect 2532 8186 2556 8188
rect 2612 8186 2636 8188
rect 2692 8186 2706 8188
rect 1746 8134 1756 8186
rect 1812 8134 1822 8186
rect 2066 8134 2076 8186
rect 2132 8134 2142 8186
rect 2386 8134 2396 8186
rect 2452 8134 2462 8186
rect 1502 8132 1516 8134
rect 1572 8132 1596 8134
rect 1652 8132 1676 8134
rect 1732 8132 1756 8134
rect 1812 8132 1836 8134
rect 1892 8132 1916 8134
rect 1972 8132 1996 8134
rect 2052 8132 2076 8134
rect 2132 8132 2156 8134
rect 2212 8132 2236 8134
rect 2292 8132 2316 8134
rect 2372 8132 2396 8134
rect 2452 8132 2476 8134
rect 2532 8132 2556 8134
rect 2612 8132 2636 8134
rect 2692 8132 2706 8134
rect 1502 8123 2706 8132
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2148 7886 2176 8026
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2148 7206 2176 7822
rect 2792 7818 2820 8366
rect 2976 8344 3004 8910
rect 3056 8356 3108 8362
rect 2976 8316 3056 8344
rect 3056 8298 3108 8304
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2700 7546 2728 7754
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2884 7410 2912 7890
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7478 3096 7686
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 1320 7126 1440 7154
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 1216 4684 1268 4690
rect 1216 4626 1268 4632
rect 1320 3890 1348 7126
rect 1502 7100 2706 7109
rect 1502 7098 1516 7100
rect 1572 7098 1596 7100
rect 1652 7098 1676 7100
rect 1732 7098 1756 7100
rect 1812 7098 1836 7100
rect 1892 7098 1916 7100
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 2292 7098 2316 7100
rect 2372 7098 2396 7100
rect 2452 7098 2476 7100
rect 2532 7098 2556 7100
rect 2612 7098 2636 7100
rect 2692 7098 2706 7100
rect 1746 7046 1756 7098
rect 1812 7046 1822 7098
rect 2066 7046 2076 7098
rect 2132 7046 2142 7098
rect 2386 7046 2396 7098
rect 2452 7046 2462 7098
rect 1502 7044 1516 7046
rect 1572 7044 1596 7046
rect 1652 7044 1676 7046
rect 1732 7044 1756 7046
rect 1812 7044 1836 7046
rect 1892 7044 1916 7046
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 2292 7044 2316 7046
rect 2372 7044 2396 7046
rect 2452 7044 2476 7046
rect 2532 7044 2556 7046
rect 2612 7044 2636 7046
rect 2692 7044 2706 7046
rect 1502 7035 2706 7044
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1412 4049 1440 6938
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2240 6390 2268 6666
rect 2700 6458 2728 6666
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 2792 6322 2820 6802
rect 2976 6730 3004 7414
rect 3160 6798 3188 9318
rect 3252 6798 3280 12600
rect 3344 10198 3372 15302
rect 3436 15162 3464 15370
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3436 14278 3464 15098
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3436 12238 3464 14010
rect 3528 13161 3556 16050
rect 3514 13152 3570 13161
rect 3514 13087 3570 13096
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3422 11928 3478 11937
rect 3422 11863 3478 11872
rect 3436 11830 3464 11863
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3436 11354 3464 11766
rect 3528 11626 3556 12854
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3528 11200 3556 11562
rect 3436 11172 3556 11200
rect 3436 10674 3464 11172
rect 3620 11098 3648 16458
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3712 15162 3740 16050
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3712 12918 3740 14350
rect 3700 12912 3752 12918
rect 3700 12854 3752 12860
rect 3804 12594 3832 15574
rect 3896 15366 3924 17002
rect 4356 16522 4384 17138
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 4344 16516 4396 16522
rect 4344 16458 4396 16464
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3528 11070 3648 11098
rect 3712 12566 3832 12594
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3332 10192 3384 10198
rect 3332 10134 3384 10140
rect 3344 10062 3372 10134
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3422 10024 3478 10033
rect 3422 9959 3478 9968
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 7002 3372 8774
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 3160 6254 3188 6734
rect 3252 6662 3280 6734
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 1502 6012 2706 6021
rect 1502 6010 1516 6012
rect 1572 6010 1596 6012
rect 1652 6010 1676 6012
rect 1732 6010 1756 6012
rect 1812 6010 1836 6012
rect 1892 6010 1916 6012
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 2292 6010 2316 6012
rect 2372 6010 2396 6012
rect 2452 6010 2476 6012
rect 2532 6010 2556 6012
rect 2612 6010 2636 6012
rect 2692 6010 2706 6012
rect 1746 5958 1756 6010
rect 1812 5958 1822 6010
rect 2066 5958 2076 6010
rect 2132 5958 2142 6010
rect 2386 5958 2396 6010
rect 2452 5958 2462 6010
rect 1502 5956 1516 5958
rect 1572 5956 1596 5958
rect 1652 5956 1676 5958
rect 1732 5956 1756 5958
rect 1812 5956 1836 5958
rect 1892 5956 1916 5958
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 2292 5956 2316 5958
rect 2372 5956 2396 5958
rect 2452 5956 2476 5958
rect 2532 5956 2556 5958
rect 2612 5956 2636 5958
rect 2692 5956 2706 5958
rect 1502 5947 2706 5956
rect 2884 5846 2912 6190
rect 3436 5896 3464 9959
rect 3252 5868 3464 5896
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2320 5636 2372 5642
rect 2320 5578 2372 5584
rect 2332 5234 2360 5578
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 5302 3096 5510
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 1502 4924 2706 4933
rect 1502 4922 1516 4924
rect 1572 4922 1596 4924
rect 1652 4922 1676 4924
rect 1732 4922 1756 4924
rect 1812 4922 1836 4924
rect 1892 4922 1916 4924
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 2292 4922 2316 4924
rect 2372 4922 2396 4924
rect 2452 4922 2476 4924
rect 2532 4922 2556 4924
rect 2612 4922 2636 4924
rect 2692 4922 2706 4924
rect 1746 4870 1756 4922
rect 1812 4870 1822 4922
rect 2066 4870 2076 4922
rect 2132 4870 2142 4922
rect 2386 4870 2396 4922
rect 2452 4870 2462 4922
rect 1502 4868 1516 4870
rect 1572 4868 1596 4870
rect 1652 4868 1676 4870
rect 1732 4868 1756 4870
rect 1812 4868 1836 4870
rect 1892 4868 1916 4870
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 2292 4868 2316 4870
rect 2372 4868 2396 4870
rect 2452 4868 2476 4870
rect 2532 4868 2556 4870
rect 2612 4868 2636 4870
rect 2692 4868 2706 4870
rect 1502 4859 2706 4868
rect 2792 4554 2820 5102
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4146 2360 4422
rect 2700 4282 2728 4490
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 3068 4214 3096 4626
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 3160 4146 3188 4558
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 1398 4040 1454 4049
rect 1398 3975 1454 3984
rect 1400 3936 1452 3942
rect 1320 3884 1400 3890
rect 1320 3878 1452 3884
rect 1320 3862 1440 3878
rect 1502 3836 2706 3845
rect 1502 3834 1516 3836
rect 1572 3834 1596 3836
rect 1652 3834 1676 3836
rect 1732 3834 1756 3836
rect 1812 3834 1836 3836
rect 1892 3834 1916 3836
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 2292 3834 2316 3836
rect 2372 3834 2396 3836
rect 2452 3834 2476 3836
rect 2532 3834 2556 3836
rect 2612 3834 2636 3836
rect 2692 3834 2706 3836
rect 1746 3782 1756 3834
rect 1812 3782 1822 3834
rect 2066 3782 2076 3834
rect 2132 3782 2142 3834
rect 2386 3782 2396 3834
rect 2452 3782 2462 3834
rect 1502 3780 1516 3782
rect 1572 3780 1596 3782
rect 1652 3780 1676 3782
rect 1732 3780 1756 3782
rect 1812 3780 1836 3782
rect 1892 3780 1916 3782
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 2292 3780 2316 3782
rect 2372 3780 2396 3782
rect 2452 3780 2476 3782
rect 2532 3780 2556 3782
rect 2612 3780 2636 3782
rect 2692 3780 2706 3782
rect 1502 3771 2706 3780
rect 2792 3670 2820 4082
rect 1400 3664 1452 3670
rect 1400 3606 1452 3612
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 1122 3496 1178 3505
rect 1122 3431 1178 3440
rect 1030 3224 1086 3233
rect 1030 3159 1086 3168
rect 1124 2984 1176 2990
rect 938 2952 994 2961
rect 1124 2926 1176 2932
rect 938 2887 994 2896
rect 768 2746 1072 2774
rect 124 800 152 2746
rect 940 2576 992 2582
rect 940 2518 992 2524
rect 952 2417 980 2518
rect 938 2408 994 2417
rect 938 2343 994 2352
rect 1044 2145 1072 2746
rect 1030 2136 1086 2145
rect 1030 2071 1086 2080
rect 1136 1329 1164 2926
rect 1412 2650 1440 3606
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 3058 1624 3334
rect 2424 3126 2452 3402
rect 2700 3194 2728 3402
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 2884 2990 2912 3470
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 3252 2774 3280 5868
rect 3528 5794 3556 11070
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3620 10742 3648 10950
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3620 5914 3648 8298
rect 3712 8022 3740 12566
rect 3896 12481 3924 15302
rect 3988 13938 4016 16458
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4080 15094 4108 15438
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3882 12472 3938 12481
rect 3882 12407 3938 12416
rect 3988 12288 4016 13874
rect 4080 13025 4108 14894
rect 4172 14550 4200 15438
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4264 15026 4292 15302
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4252 14884 4304 14890
rect 4252 14826 4304 14832
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 13870 4200 14214
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13433 4200 13806
rect 4158 13424 4214 13433
rect 4158 13359 4214 13368
rect 4264 13376 4292 14826
rect 4356 14618 4384 15030
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4356 13818 4384 14554
rect 4448 14006 4476 17274
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4540 15910 4568 16934
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15366 4568 15846
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4540 14618 4568 14962
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4526 14512 4582 14521
rect 4526 14447 4582 14456
rect 4540 14414 4568 14447
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4540 14249 4568 14350
rect 4526 14240 4582 14249
rect 4526 14175 4582 14184
rect 4526 14104 4582 14113
rect 4526 14039 4528 14048
rect 4580 14039 4582 14048
rect 4528 14010 4580 14016
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4356 13790 4568 13818
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4448 13569 4476 13670
rect 4434 13560 4490 13569
rect 4434 13495 4490 13504
rect 4172 13326 4200 13359
rect 4264 13348 4384 13376
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4250 13288 4306 13297
rect 4250 13223 4306 13232
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4066 13016 4122 13025
rect 4172 12986 4200 13126
rect 4066 12951 4122 12960
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4264 12850 4292 13223
rect 4356 12850 4384 13348
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4252 12844 4304 12850
rect 3896 12260 4016 12288
rect 4080 12804 4252 12832
rect 3896 12102 3924 12260
rect 4080 12152 4108 12804
rect 4252 12786 4304 12792
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4356 12730 4384 12786
rect 4172 12702 4384 12730
rect 4172 12442 4200 12702
rect 4448 12594 4476 12854
rect 4263 12566 4476 12594
rect 4160 12436 4212 12442
rect 4263 12434 4291 12566
rect 4263 12406 4292 12434
rect 4160 12378 4212 12384
rect 4264 12306 4292 12406
rect 4434 12336 4490 12345
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4252 12300 4304 12306
rect 4304 12260 4384 12288
rect 4434 12271 4490 12280
rect 4252 12242 4304 12248
rect 3988 12124 4108 12152
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3790 11792 3846 11801
rect 3790 11727 3792 11736
rect 3844 11727 3846 11736
rect 3792 11698 3844 11704
rect 3804 10674 3832 11698
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3896 10606 3924 11834
rect 3988 11558 4016 12124
rect 4172 12050 4200 12242
rect 4080 12022 4200 12050
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 11121 4016 11494
rect 4080 11150 4108 12022
rect 4264 11914 4292 12038
rect 4172 11886 4292 11914
rect 4068 11144 4120 11150
rect 3974 11112 4030 11121
rect 4068 11086 4120 11092
rect 3974 11047 4030 11056
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10810 4016 10950
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4080 10656 4108 11086
rect 4172 11014 4200 11886
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4158 10840 4214 10849
rect 4158 10775 4214 10784
rect 3988 10628 4108 10656
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3988 10470 4016 10628
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3712 7886 3740 7958
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3344 5766 3556 5794
rect 3344 5710 3372 5766
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3528 5642 3556 5766
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3620 5234 3648 5850
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 1502 2748 2706 2757
rect 1502 2746 1516 2748
rect 1572 2746 1596 2748
rect 1652 2746 1676 2748
rect 1732 2746 1756 2748
rect 1812 2746 1836 2748
rect 1892 2746 1916 2748
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 2292 2746 2316 2748
rect 2372 2746 2396 2748
rect 2452 2746 2476 2748
rect 2532 2746 2556 2748
rect 2612 2746 2636 2748
rect 2692 2746 2706 2748
rect 1746 2694 1756 2746
rect 1812 2694 1822 2746
rect 2066 2694 2076 2746
rect 2132 2694 2142 2746
rect 2386 2694 2396 2746
rect 2452 2694 2462 2746
rect 1502 2692 1516 2694
rect 1572 2692 1596 2694
rect 1652 2692 1676 2694
rect 1732 2692 1756 2694
rect 1812 2692 1836 2694
rect 1892 2692 1916 2694
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 2292 2692 2316 2694
rect 2372 2692 2396 2694
rect 2452 2692 2476 2694
rect 2532 2692 2556 2694
rect 2612 2692 2636 2694
rect 2692 2692 2706 2694
rect 1502 2683 2706 2692
rect 3160 2746 3280 2774
rect 1400 2644 1452 2650
rect 1400 2586 1452 2592
rect 3160 2446 3188 2746
rect 3344 2446 3372 3470
rect 3712 2553 3740 7278
rect 3988 4690 4016 9658
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3988 3534 4016 3674
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3698 2544 3754 2553
rect 3698 2479 3754 2488
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 3422 1864 3478 1873
rect 3422 1799 3424 1808
rect 3476 1799 3478 1808
rect 3424 1770 3476 1776
rect 3528 1601 3556 2042
rect 3514 1592 3570 1601
rect 3514 1527 3570 1536
rect 3424 1352 3476 1358
rect 1122 1320 1178 1329
rect 3424 1294 3476 1300
rect 1122 1255 1178 1264
rect 3332 1216 3384 1222
rect 3332 1158 3384 1164
rect 296 1012 348 1018
rect 296 954 348 960
rect 308 800 336 954
rect 110 0 166 800
rect 294 0 350 800
rect 3344 785 3372 1158
rect 3330 776 3386 785
rect 3330 711 3386 720
rect 3436 513 3464 1294
rect 4080 1290 4108 10503
rect 4172 9081 4200 10775
rect 4158 9072 4214 9081
rect 4158 9007 4214 9016
rect 4172 8294 4200 9007
rect 4264 8566 4292 11698
rect 4356 10849 4384 12260
rect 4448 12238 4476 12271
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4448 11694 4476 12174
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4342 10840 4398 10849
rect 4342 10775 4398 10784
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4172 8266 4292 8294
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4172 5370 4200 5714
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4264 5250 4292 8266
rect 4356 5370 4384 10542
rect 4448 8906 4476 11222
rect 4540 10742 4568 13790
rect 4632 11898 4660 16118
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4632 11218 4660 11494
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4632 10985 4660 11018
rect 4724 11014 4752 15846
rect 4816 14958 4844 16526
rect 4908 15638 4936 17138
rect 5446 16688 5502 16697
rect 5446 16623 5502 16632
rect 5460 16590 5488 16623
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 4988 16516 5040 16522
rect 4988 16458 5040 16464
rect 5000 15910 5028 16458
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 5000 15484 5028 15846
rect 4908 15456 5028 15484
rect 5170 15464 5226 15473
rect 4804 14952 4856 14958
rect 4908 14929 4936 15456
rect 5170 15399 5172 15408
rect 5224 15399 5226 15408
rect 5172 15370 5224 15376
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5000 15065 5028 15302
rect 4986 15056 5042 15065
rect 4986 14991 5042 15000
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 4804 14894 4856 14900
rect 4894 14920 4950 14929
rect 4894 14855 4950 14864
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4816 13870 4844 14486
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4816 13462 4844 13806
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4816 11762 4844 13262
rect 4908 12889 4936 14758
rect 5092 14618 5120 14962
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 5000 13530 5028 14486
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 5092 13938 5120 14350
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5078 13832 5134 13841
rect 5078 13767 5134 13776
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 5092 13376 5120 13767
rect 5184 13530 5212 14962
rect 5276 14634 5304 15982
rect 5368 15858 5396 16526
rect 5502 16348 6706 16357
rect 5502 16346 5516 16348
rect 5572 16346 5596 16348
rect 5652 16346 5676 16348
rect 5732 16346 5756 16348
rect 5812 16346 5836 16348
rect 5892 16346 5916 16348
rect 5972 16346 5996 16348
rect 6052 16346 6076 16348
rect 6132 16346 6156 16348
rect 6212 16346 6236 16348
rect 6292 16346 6316 16348
rect 6372 16346 6396 16348
rect 6452 16346 6476 16348
rect 6532 16346 6556 16348
rect 6612 16346 6636 16348
rect 6692 16346 6706 16348
rect 5746 16294 5756 16346
rect 5812 16294 5822 16346
rect 6066 16294 6076 16346
rect 6132 16294 6142 16346
rect 6386 16294 6396 16346
rect 6452 16294 6462 16346
rect 5502 16292 5516 16294
rect 5572 16292 5596 16294
rect 5652 16292 5676 16294
rect 5732 16292 5756 16294
rect 5812 16292 5836 16294
rect 5892 16292 5916 16294
rect 5972 16292 5996 16294
rect 6052 16292 6076 16294
rect 6132 16292 6156 16294
rect 6212 16292 6236 16294
rect 6292 16292 6316 16294
rect 6372 16292 6396 16294
rect 6452 16292 6476 16294
rect 6532 16292 6556 16294
rect 6612 16292 6636 16294
rect 6692 16292 6706 16294
rect 5502 16283 6706 16292
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 5368 15830 5488 15858
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5368 14804 5396 15642
rect 5460 15609 5488 15830
rect 6182 15736 6238 15745
rect 6288 15706 6316 16118
rect 6748 15910 6776 16526
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6182 15671 6184 15680
rect 6236 15671 6238 15680
rect 6276 15700 6328 15706
rect 6184 15642 6236 15648
rect 6276 15642 6328 15648
rect 5446 15600 5502 15609
rect 5446 15535 5502 15544
rect 6288 15434 6316 15642
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 5502 15260 6706 15269
rect 5502 15258 5516 15260
rect 5572 15258 5596 15260
rect 5652 15258 5676 15260
rect 5732 15258 5756 15260
rect 5812 15258 5836 15260
rect 5892 15258 5916 15260
rect 5972 15258 5996 15260
rect 6052 15258 6076 15260
rect 6132 15258 6156 15260
rect 6212 15258 6236 15260
rect 6292 15258 6316 15260
rect 6372 15258 6396 15260
rect 6452 15258 6476 15260
rect 6532 15258 6556 15260
rect 6612 15258 6636 15260
rect 6692 15258 6706 15260
rect 5746 15206 5756 15258
rect 5812 15206 5822 15258
rect 6066 15206 6076 15258
rect 6132 15206 6142 15258
rect 6386 15206 6396 15258
rect 6452 15206 6462 15258
rect 5502 15204 5516 15206
rect 5572 15204 5596 15206
rect 5652 15204 5676 15206
rect 5732 15204 5756 15206
rect 5812 15204 5836 15206
rect 5892 15204 5916 15206
rect 5972 15204 5996 15206
rect 6052 15204 6076 15206
rect 6132 15204 6156 15206
rect 6212 15204 6236 15206
rect 6292 15204 6316 15206
rect 6372 15204 6396 15206
rect 6452 15204 6476 15206
rect 6532 15204 6556 15206
rect 6612 15204 6636 15206
rect 6692 15204 6706 15206
rect 5502 15195 6706 15204
rect 6552 15088 6604 15094
rect 5630 15056 5686 15065
rect 5630 14991 5686 15000
rect 6550 15056 6552 15065
rect 6604 15056 6606 15065
rect 6550 14991 6606 15000
rect 5540 14816 5592 14822
rect 5368 14776 5540 14804
rect 5540 14758 5592 14764
rect 5446 14648 5502 14657
rect 5276 14606 5396 14634
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5276 13376 5304 14214
rect 5368 14056 5396 14606
rect 5446 14583 5502 14592
rect 5460 14482 5488 14583
rect 5552 14521 5580 14758
rect 5538 14512 5594 14521
rect 5448 14476 5500 14482
rect 5538 14447 5594 14456
rect 5448 14418 5500 14424
rect 5644 14385 5672 14991
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 5816 14816 5868 14822
rect 5722 14784 5778 14793
rect 5816 14758 5868 14764
rect 5722 14719 5778 14728
rect 5736 14414 5764 14719
rect 5828 14550 5856 14758
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 5724 14408 5776 14414
rect 5630 14376 5686 14385
rect 5724 14350 5776 14356
rect 6012 14346 6040 14894
rect 6644 14816 6696 14822
rect 6458 14784 6514 14793
rect 6644 14758 6696 14764
rect 6458 14719 6514 14728
rect 6274 14512 6330 14521
rect 6274 14447 6276 14456
rect 6328 14447 6330 14456
rect 6276 14418 6328 14424
rect 6472 14414 6500 14719
rect 6656 14657 6684 14758
rect 6642 14648 6698 14657
rect 6642 14583 6698 14592
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 5630 14311 5686 14320
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 5502 14172 6706 14181
rect 5502 14170 5516 14172
rect 5572 14170 5596 14172
rect 5652 14170 5676 14172
rect 5732 14170 5756 14172
rect 5812 14170 5836 14172
rect 5892 14170 5916 14172
rect 5972 14170 5996 14172
rect 6052 14170 6076 14172
rect 6132 14170 6156 14172
rect 6212 14170 6236 14172
rect 6292 14170 6316 14172
rect 6372 14170 6396 14172
rect 6452 14170 6476 14172
rect 6532 14170 6556 14172
rect 6612 14170 6636 14172
rect 6692 14170 6706 14172
rect 5746 14118 5756 14170
rect 5812 14118 5822 14170
rect 6066 14118 6076 14170
rect 6132 14118 6142 14170
rect 6386 14118 6396 14170
rect 6452 14118 6462 14170
rect 5502 14116 5516 14118
rect 5572 14116 5596 14118
rect 5652 14116 5676 14118
rect 5732 14116 5756 14118
rect 5812 14116 5836 14118
rect 5892 14116 5916 14118
rect 5972 14116 5996 14118
rect 6052 14116 6076 14118
rect 6132 14116 6156 14118
rect 6212 14116 6236 14118
rect 6292 14116 6316 14118
rect 6372 14116 6396 14118
rect 6452 14116 6476 14118
rect 6532 14116 6556 14118
rect 6612 14116 6636 14118
rect 6692 14116 6706 14118
rect 5502 14107 6706 14116
rect 5368 14028 5764 14056
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5538 13560 5594 13569
rect 5448 13524 5500 13530
rect 5538 13495 5540 13504
rect 5448 13466 5500 13472
rect 5592 13495 5594 13504
rect 5540 13466 5592 13472
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5000 13348 5120 13376
rect 5184 13348 5304 13376
rect 5000 13025 5028 13348
rect 5184 13297 5212 13348
rect 5170 13288 5226 13297
rect 5080 13252 5132 13258
rect 5368 13240 5396 13398
rect 5170 13223 5226 13232
rect 5080 13194 5132 13200
rect 5276 13212 5396 13240
rect 4986 13016 5042 13025
rect 4986 12951 5042 12960
rect 5000 12918 5028 12951
rect 4988 12912 5040 12918
rect 4894 12880 4950 12889
rect 4988 12854 5040 12860
rect 4894 12815 4950 12824
rect 4894 12472 4950 12481
rect 5092 12424 5120 13194
rect 5276 13172 5304 13212
rect 5460 13190 5488 13466
rect 5644 13462 5672 13670
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 5736 13297 5764 14028
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5920 13569 5948 13942
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 5906 13560 5962 13569
rect 5906 13495 5962 13504
rect 6472 13326 6500 13874
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6656 13326 6684 13738
rect 6460 13320 6512 13326
rect 5722 13288 5778 13297
rect 6644 13320 6696 13326
rect 6460 13262 6512 13268
rect 6642 13288 6644 13297
rect 6696 13288 6698 13297
rect 5722 13223 5778 13232
rect 6642 13223 6698 13232
rect 5448 13184 5500 13190
rect 5276 13144 5396 13172
rect 5170 13016 5226 13025
rect 5170 12951 5226 12960
rect 5368 12968 5396 13144
rect 5448 13126 5500 13132
rect 5502 13084 6706 13093
rect 5502 13082 5516 13084
rect 5572 13082 5596 13084
rect 5652 13082 5676 13084
rect 5732 13082 5756 13084
rect 5812 13082 5836 13084
rect 5892 13082 5916 13084
rect 5972 13082 5996 13084
rect 6052 13082 6076 13084
rect 6132 13082 6156 13084
rect 6212 13082 6236 13084
rect 6292 13082 6316 13084
rect 6372 13082 6396 13084
rect 6452 13082 6476 13084
rect 6532 13082 6556 13084
rect 6612 13082 6636 13084
rect 6692 13082 6706 13084
rect 5746 13030 5756 13082
rect 5812 13030 5822 13082
rect 6066 13030 6076 13082
rect 6132 13030 6142 13082
rect 6386 13030 6396 13082
rect 6452 13030 6462 13082
rect 5502 13028 5516 13030
rect 5572 13028 5596 13030
rect 5652 13028 5676 13030
rect 5732 13028 5756 13030
rect 5812 13028 5836 13030
rect 5892 13028 5916 13030
rect 5972 13028 5996 13030
rect 6052 13028 6076 13030
rect 6132 13028 6156 13030
rect 6212 13028 6236 13030
rect 6292 13028 6316 13030
rect 6372 13028 6396 13030
rect 6452 13028 6476 13030
rect 6532 13028 6556 13030
rect 6612 13028 6636 13030
rect 6692 13028 6706 13030
rect 5502 13019 6706 13028
rect 6184 12980 6236 12986
rect 5184 12832 5212 12951
rect 5368 12940 5580 12968
rect 5552 12850 5580 12940
rect 6184 12922 6236 12928
rect 5814 12880 5870 12889
rect 5540 12844 5592 12850
rect 5184 12804 5396 12832
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5184 12442 5212 12650
rect 4894 12407 4896 12416
rect 4948 12407 4950 12416
rect 4896 12378 4948 12384
rect 5000 12396 5120 12424
rect 5172 12436 5224 12442
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4908 11608 4936 12174
rect 4816 11580 4936 11608
rect 4816 11286 4844 11580
rect 4894 11520 4950 11529
rect 4894 11455 4950 11464
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4712 11008 4764 11014
rect 4618 10976 4674 10985
rect 4712 10950 4764 10956
rect 4618 10911 4674 10920
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4448 6254 4476 8570
rect 4540 8498 4568 9590
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4540 6322 4568 8434
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4264 5222 4476 5250
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4172 2650 4200 3470
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4448 2514 4476 5222
rect 4632 2922 4660 10746
rect 4724 10674 4752 10950
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4724 9654 4752 9998
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 3602 4752 9318
rect 4816 3670 4844 11086
rect 4908 10810 4936 11455
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 5000 10606 5028 12396
rect 5172 12378 5224 12384
rect 5276 12345 5304 12650
rect 5262 12336 5318 12345
rect 5080 12300 5132 12306
rect 5262 12271 5318 12280
rect 5080 12242 5132 12248
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4908 7546 4936 10202
rect 5000 10033 5028 10202
rect 4986 10024 5042 10033
rect 4986 9959 5042 9968
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 5914 4936 6258
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4908 5234 4936 5850
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4908 2774 4936 5170
rect 5000 4078 5028 9862
rect 5092 9722 5120 12242
rect 5172 12164 5224 12170
rect 5172 12106 5224 12112
rect 5184 11762 5212 12106
rect 5276 11762 5304 12271
rect 5368 12170 5396 12804
rect 5448 12810 5500 12816
rect 5814 12815 5870 12824
rect 5540 12786 5592 12792
rect 5448 12752 5500 12758
rect 5460 12345 5488 12752
rect 5552 12374 5580 12786
rect 5722 12744 5778 12753
rect 5722 12679 5778 12688
rect 5540 12368 5592 12374
rect 5446 12336 5502 12345
rect 5632 12368 5684 12374
rect 5540 12310 5592 12316
rect 5630 12336 5632 12345
rect 5684 12336 5686 12345
rect 5446 12271 5502 12280
rect 5630 12271 5686 12280
rect 5540 12232 5592 12238
rect 5736 12186 5764 12679
rect 5828 12238 5856 12815
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12306 5948 12582
rect 6012 12481 6040 12718
rect 5998 12472 6054 12481
rect 5998 12407 6054 12416
rect 6196 12345 6224 12922
rect 6550 12880 6606 12889
rect 6748 12850 6776 15370
rect 6840 14396 6868 16050
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6932 14521 6960 15846
rect 7194 15736 7250 15745
rect 7194 15671 7250 15680
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6918 14512 6974 14521
rect 6918 14447 6974 14456
rect 6840 14368 6960 14396
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 13705 6868 14214
rect 6932 13734 6960 14368
rect 6920 13728 6972 13734
rect 6826 13696 6882 13705
rect 6920 13670 6972 13676
rect 6826 13631 6882 13640
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6840 12850 6868 13466
rect 6550 12815 6606 12824
rect 6736 12844 6788 12850
rect 6564 12714 6592 12815
rect 6736 12786 6788 12792
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6826 12744 6882 12753
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6644 12708 6696 12714
rect 6932 12714 6960 13670
rect 6826 12679 6882 12688
rect 6920 12708 6972 12714
rect 6644 12650 6696 12656
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12458 6408 12582
rect 6276 12436 6328 12442
rect 6380 12430 6500 12458
rect 6276 12378 6328 12384
rect 6182 12336 6238 12345
rect 5908 12300 5960 12306
rect 6182 12271 6238 12280
rect 5908 12242 5960 12248
rect 5592 12180 5764 12186
rect 5540 12174 5764 12180
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5356 12164 5408 12170
rect 5552 12158 5764 12174
rect 6288 12170 6316 12378
rect 6472 12209 6500 12430
rect 6656 12209 6684 12650
rect 6458 12200 6514 12209
rect 6276 12164 6328 12170
rect 5356 12106 5408 12112
rect 6458 12135 6514 12144
rect 6642 12200 6698 12209
rect 6642 12135 6698 12144
rect 6276 12106 6328 12112
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5262 11656 5318 11665
rect 5262 11591 5264 11600
rect 5316 11591 5318 11600
rect 5264 11562 5316 11568
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5078 9616 5134 9625
rect 5078 9551 5134 9560
rect 5092 8498 5120 9551
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 5092 6458 5120 8298
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5092 2938 5120 4422
rect 5184 3058 5212 11222
rect 5276 10713 5304 11562
rect 5262 10704 5318 10713
rect 5262 10639 5318 10648
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 9586 5304 10406
rect 5368 9722 5396 12106
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 5502 11996 6706 12005
rect 5502 11994 5516 11996
rect 5572 11994 5596 11996
rect 5652 11994 5676 11996
rect 5732 11994 5756 11996
rect 5812 11994 5836 11996
rect 5892 11994 5916 11996
rect 5972 11994 5996 11996
rect 6052 11994 6076 11996
rect 6132 11994 6156 11996
rect 6212 11994 6236 11996
rect 6292 11994 6316 11996
rect 6372 11994 6396 11996
rect 6452 11994 6476 11996
rect 6532 11994 6556 11996
rect 6612 11994 6636 11996
rect 6692 11994 6706 11996
rect 5746 11942 5756 11994
rect 5812 11942 5822 11994
rect 6066 11942 6076 11994
rect 6132 11942 6142 11994
rect 6386 11942 6396 11994
rect 6452 11942 6462 11994
rect 5502 11940 5516 11942
rect 5572 11940 5596 11942
rect 5652 11940 5676 11942
rect 5732 11940 5756 11942
rect 5812 11940 5836 11942
rect 5892 11940 5916 11942
rect 5972 11940 5996 11942
rect 6052 11940 6076 11942
rect 6132 11940 6156 11942
rect 6212 11940 6236 11942
rect 6292 11940 6316 11942
rect 6372 11940 6396 11942
rect 6452 11940 6476 11942
rect 6532 11940 6556 11942
rect 6612 11940 6636 11942
rect 6692 11940 6706 11942
rect 5502 11931 6706 11940
rect 6368 11824 6420 11830
rect 5630 11792 5686 11801
rect 6368 11766 6420 11772
rect 5630 11727 5632 11736
rect 5684 11727 5686 11736
rect 5816 11756 5868 11762
rect 5632 11698 5684 11704
rect 5816 11698 5868 11704
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5828 11529 5856 11698
rect 5814 11520 5870 11529
rect 5814 11455 5870 11464
rect 5920 11286 5948 11698
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6012 11393 6040 11630
rect 5998 11384 6054 11393
rect 5998 11319 6054 11328
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 6380 11082 6408 11766
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6472 11286 6500 11562
rect 6550 11520 6606 11529
rect 6550 11455 6606 11464
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6564 10996 6592 11455
rect 6748 11064 6776 12038
rect 6840 11801 6868 12679
rect 6920 12650 6972 12656
rect 6918 12336 6974 12345
rect 6918 12271 6974 12280
rect 6826 11792 6882 11801
rect 6826 11727 6882 11736
rect 6932 11608 6960 12271
rect 7024 12238 7052 15370
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7010 12064 7066 12073
rect 7010 11999 7066 12008
rect 7024 11626 7052 11999
rect 6840 11580 6960 11608
rect 7012 11620 7064 11626
rect 6840 11132 6868 11580
rect 7012 11562 7064 11568
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6840 11104 6960 11132
rect 6748 11036 6868 11064
rect 6564 10968 6776 10996
rect 5502 10908 6706 10917
rect 5502 10906 5516 10908
rect 5572 10906 5596 10908
rect 5652 10906 5676 10908
rect 5732 10906 5756 10908
rect 5812 10906 5836 10908
rect 5892 10906 5916 10908
rect 5972 10906 5996 10908
rect 6052 10906 6076 10908
rect 6132 10906 6156 10908
rect 6212 10906 6236 10908
rect 6292 10906 6316 10908
rect 6372 10906 6396 10908
rect 6452 10906 6476 10908
rect 6532 10906 6556 10908
rect 6612 10906 6636 10908
rect 6692 10906 6706 10908
rect 5746 10854 5756 10906
rect 5812 10854 5822 10906
rect 6066 10854 6076 10906
rect 6132 10854 6142 10906
rect 6386 10854 6396 10906
rect 6452 10854 6462 10906
rect 5502 10852 5516 10854
rect 5572 10852 5596 10854
rect 5652 10852 5676 10854
rect 5732 10852 5756 10854
rect 5812 10852 5836 10854
rect 5892 10852 5916 10854
rect 5972 10852 5996 10854
rect 6052 10852 6076 10854
rect 6132 10852 6156 10854
rect 6212 10852 6236 10854
rect 6292 10852 6316 10854
rect 6372 10852 6396 10854
rect 6452 10852 6476 10854
rect 6532 10852 6556 10854
rect 6612 10852 6636 10854
rect 6692 10852 6706 10854
rect 5502 10843 6706 10852
rect 6748 10792 6776 10968
rect 6564 10764 6776 10792
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10062 5488 10610
rect 5540 10600 5592 10606
rect 5538 10568 5540 10577
rect 5592 10568 5594 10577
rect 6564 10538 6592 10764
rect 6840 10724 6868 11036
rect 6748 10696 6868 10724
rect 5538 10503 5594 10512
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6564 10305 6592 10474
rect 6550 10296 6606 10305
rect 6550 10231 6606 10240
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 6642 10024 6698 10033
rect 6642 9959 6698 9968
rect 6656 9926 6684 9959
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 5502 9820 6706 9829
rect 5502 9818 5516 9820
rect 5572 9818 5596 9820
rect 5652 9818 5676 9820
rect 5732 9818 5756 9820
rect 5812 9818 5836 9820
rect 5892 9818 5916 9820
rect 5972 9818 5996 9820
rect 6052 9818 6076 9820
rect 6132 9818 6156 9820
rect 6212 9818 6236 9820
rect 6292 9818 6316 9820
rect 6372 9818 6396 9820
rect 6452 9818 6476 9820
rect 6532 9818 6556 9820
rect 6612 9818 6636 9820
rect 6692 9818 6706 9820
rect 5746 9766 5756 9818
rect 5812 9766 5822 9818
rect 6066 9766 6076 9818
rect 6132 9766 6142 9818
rect 6386 9766 6396 9818
rect 6452 9766 6462 9818
rect 5502 9764 5516 9766
rect 5572 9764 5596 9766
rect 5652 9764 5676 9766
rect 5732 9764 5756 9766
rect 5812 9764 5836 9766
rect 5892 9764 5916 9766
rect 5972 9764 5996 9766
rect 6052 9764 6076 9766
rect 6132 9764 6156 9766
rect 6212 9764 6236 9766
rect 6292 9764 6316 9766
rect 6372 9764 6396 9766
rect 6452 9764 6476 9766
rect 6532 9764 6556 9766
rect 6612 9764 6636 9766
rect 6692 9764 6706 9766
rect 5502 9755 6706 9764
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5276 8906 5304 9114
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5276 8498 5304 8842
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5276 6390 5304 8298
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5264 6248 5316 6254
rect 5368 6225 5396 9454
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6564 8974 6592 9386
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 5502 8732 6706 8741
rect 5502 8730 5516 8732
rect 5572 8730 5596 8732
rect 5652 8730 5676 8732
rect 5732 8730 5756 8732
rect 5812 8730 5836 8732
rect 5892 8730 5916 8732
rect 5972 8730 5996 8732
rect 6052 8730 6076 8732
rect 6132 8730 6156 8732
rect 6212 8730 6236 8732
rect 6292 8730 6316 8732
rect 6372 8730 6396 8732
rect 6452 8730 6476 8732
rect 6532 8730 6556 8732
rect 6612 8730 6636 8732
rect 6692 8730 6706 8732
rect 5746 8678 5756 8730
rect 5812 8678 5822 8730
rect 6066 8678 6076 8730
rect 6132 8678 6142 8730
rect 6386 8678 6396 8730
rect 6452 8678 6462 8730
rect 5502 8676 5516 8678
rect 5572 8676 5596 8678
rect 5652 8676 5676 8678
rect 5732 8676 5756 8678
rect 5812 8676 5836 8678
rect 5892 8676 5916 8678
rect 5972 8676 5996 8678
rect 6052 8676 6076 8678
rect 6132 8676 6156 8678
rect 6212 8676 6236 8678
rect 6292 8676 6316 8678
rect 6372 8676 6396 8678
rect 6452 8676 6476 8678
rect 6532 8676 6556 8678
rect 6612 8676 6636 8678
rect 6692 8676 6706 8678
rect 5502 8667 6706 8676
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5460 8401 5488 8570
rect 5446 8392 5502 8401
rect 5446 8327 5502 8336
rect 5502 7644 6706 7653
rect 5502 7642 5516 7644
rect 5572 7642 5596 7644
rect 5652 7642 5676 7644
rect 5732 7642 5756 7644
rect 5812 7642 5836 7644
rect 5892 7642 5916 7644
rect 5972 7642 5996 7644
rect 6052 7642 6076 7644
rect 6132 7642 6156 7644
rect 6212 7642 6236 7644
rect 6292 7642 6316 7644
rect 6372 7642 6396 7644
rect 6452 7642 6476 7644
rect 6532 7642 6556 7644
rect 6612 7642 6636 7644
rect 6692 7642 6706 7644
rect 5746 7590 5756 7642
rect 5812 7590 5822 7642
rect 6066 7590 6076 7642
rect 6132 7590 6142 7642
rect 6386 7590 6396 7642
rect 6452 7590 6462 7642
rect 5502 7588 5516 7590
rect 5572 7588 5596 7590
rect 5652 7588 5676 7590
rect 5732 7588 5756 7590
rect 5812 7588 5836 7590
rect 5892 7588 5916 7590
rect 5972 7588 5996 7590
rect 6052 7588 6076 7590
rect 6132 7588 6156 7590
rect 6212 7588 6236 7590
rect 6292 7588 6316 7590
rect 6372 7588 6396 7590
rect 6452 7588 6476 7590
rect 6532 7588 6556 7590
rect 6612 7588 6636 7590
rect 6692 7588 6706 7590
rect 5502 7579 6706 7588
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5644 7342 5672 7482
rect 5722 7440 5778 7449
rect 5722 7375 5778 7384
rect 5736 7342 5764 7375
rect 5540 7336 5592 7342
rect 5538 7304 5540 7313
rect 5632 7336 5684 7342
rect 5592 7304 5594 7313
rect 5632 7278 5684 7284
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5538 7239 5594 7248
rect 5502 6556 6706 6565
rect 5502 6554 5516 6556
rect 5572 6554 5596 6556
rect 5652 6554 5676 6556
rect 5732 6554 5756 6556
rect 5812 6554 5836 6556
rect 5892 6554 5916 6556
rect 5972 6554 5996 6556
rect 6052 6554 6076 6556
rect 6132 6554 6156 6556
rect 6212 6554 6236 6556
rect 6292 6554 6316 6556
rect 6372 6554 6396 6556
rect 6452 6554 6476 6556
rect 6532 6554 6556 6556
rect 6612 6554 6636 6556
rect 6692 6554 6706 6556
rect 5746 6502 5756 6554
rect 5812 6502 5822 6554
rect 6066 6502 6076 6554
rect 6132 6502 6142 6554
rect 6386 6502 6396 6554
rect 6452 6502 6462 6554
rect 5502 6500 5516 6502
rect 5572 6500 5596 6502
rect 5652 6500 5676 6502
rect 5732 6500 5756 6502
rect 5812 6500 5836 6502
rect 5892 6500 5916 6502
rect 5972 6500 5996 6502
rect 6052 6500 6076 6502
rect 6132 6500 6156 6502
rect 6212 6500 6236 6502
rect 6292 6500 6316 6502
rect 6372 6500 6396 6502
rect 6452 6500 6476 6502
rect 6532 6500 6556 6502
rect 6612 6500 6636 6502
rect 6692 6500 6706 6502
rect 5502 6491 6706 6500
rect 5264 6190 5316 6196
rect 5354 6216 5410 6225
rect 5276 4758 5304 6190
rect 5354 6151 5410 6160
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6564 5710 6592 6122
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 5502 5468 6706 5477
rect 5502 5466 5516 5468
rect 5572 5466 5596 5468
rect 5652 5466 5676 5468
rect 5732 5466 5756 5468
rect 5812 5466 5836 5468
rect 5892 5466 5916 5468
rect 5972 5466 5996 5468
rect 6052 5466 6076 5468
rect 6132 5466 6156 5468
rect 6212 5466 6236 5468
rect 6292 5466 6316 5468
rect 6372 5466 6396 5468
rect 6452 5466 6476 5468
rect 6532 5466 6556 5468
rect 6612 5466 6636 5468
rect 6692 5466 6706 5468
rect 5746 5414 5756 5466
rect 5812 5414 5822 5466
rect 6066 5414 6076 5466
rect 6132 5414 6142 5466
rect 6386 5414 6396 5466
rect 6452 5414 6462 5466
rect 5502 5412 5516 5414
rect 5572 5412 5596 5414
rect 5652 5412 5676 5414
rect 5732 5412 5756 5414
rect 5812 5412 5836 5414
rect 5892 5412 5916 5414
rect 5972 5412 5996 5414
rect 6052 5412 6076 5414
rect 6132 5412 6156 5414
rect 6212 5412 6236 5414
rect 6292 5412 6316 5414
rect 6372 5412 6396 5414
rect 6452 5412 6476 5414
rect 6532 5412 6556 5414
rect 6612 5412 6636 5414
rect 6692 5412 6706 5414
rect 5502 5403 6706 5412
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5264 4752 5316 4758
rect 5264 4694 5316 4700
rect 5736 4486 5764 5306
rect 6458 5264 6514 5273
rect 6458 5199 6460 5208
rect 6512 5199 6514 5208
rect 6460 5170 6512 5176
rect 6748 5166 6776 10696
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 7954 6868 10406
rect 6932 10130 6960 11104
rect 7024 10690 7052 11290
rect 7116 10792 7144 15506
rect 7208 13870 7236 15671
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7300 15201 7328 15370
rect 7286 15192 7342 15201
rect 7286 15127 7342 15136
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7300 14346 7328 15030
rect 7392 14793 7420 16458
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7484 15337 7512 16050
rect 7576 15586 7604 17206
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7668 16017 7696 16050
rect 7654 16008 7710 16017
rect 7654 15943 7710 15952
rect 7576 15558 7696 15586
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7470 15328 7526 15337
rect 7470 15263 7526 15272
rect 7472 14816 7524 14822
rect 7378 14784 7434 14793
rect 7472 14758 7524 14764
rect 7378 14719 7434 14728
rect 7484 14482 7512 14758
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7300 14006 7328 14282
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7208 13025 7236 13806
rect 7392 13297 7420 14350
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7484 13530 7512 13874
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7576 13410 7604 15438
rect 7668 15026 7696 15558
rect 7746 15464 7802 15473
rect 7746 15399 7802 15408
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7668 14482 7696 14962
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7654 14376 7710 14385
rect 7654 14311 7710 14320
rect 7484 13382 7604 13410
rect 7378 13288 7434 13297
rect 7378 13223 7434 13232
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7194 13016 7250 13025
rect 7194 12951 7250 12960
rect 7196 12912 7248 12918
rect 7300 12900 7328 13126
rect 7248 12872 7328 12900
rect 7196 12854 7248 12860
rect 7380 12844 7432 12850
rect 7300 12804 7380 12832
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7208 12374 7236 12718
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7208 11830 7236 12310
rect 7300 12306 7328 12804
rect 7380 12786 7432 12792
rect 7484 12730 7512 13382
rect 7562 13152 7618 13161
rect 7562 13087 7618 13096
rect 7576 12918 7604 13087
rect 7564 12912 7616 12918
rect 7564 12854 7616 12860
rect 7668 12764 7696 14311
rect 7392 12702 7512 12730
rect 7576 12736 7696 12764
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7286 12200 7342 12209
rect 7286 12135 7342 12144
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7196 11824 7248 11830
rect 7196 11766 7248 11772
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7208 11286 7236 11630
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7300 10985 7328 12038
rect 7392 11354 7420 12702
rect 7576 12628 7604 12736
rect 7484 12600 7604 12628
rect 7656 12640 7708 12646
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7380 11008 7432 11014
rect 7286 10976 7342 10985
rect 7380 10950 7432 10956
rect 7286 10911 7342 10920
rect 7116 10764 7328 10792
rect 7024 10662 7236 10690
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7116 10418 7144 10542
rect 7024 10390 7144 10418
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 9722 6960 10066
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6840 7410 6868 7890
rect 6932 7546 6960 9454
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6826 6896 6882 6905
rect 6826 6831 6882 6840
rect 6840 6254 6868 6831
rect 6932 6798 6960 7210
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6564 4622 6592 5034
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4690 6776 4966
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5502 4380 6706 4389
rect 5502 4378 5516 4380
rect 5572 4378 5596 4380
rect 5652 4378 5676 4380
rect 5732 4378 5756 4380
rect 5812 4378 5836 4380
rect 5892 4378 5916 4380
rect 5972 4378 5996 4380
rect 6052 4378 6076 4380
rect 6132 4378 6156 4380
rect 6212 4378 6236 4380
rect 6292 4378 6316 4380
rect 6372 4378 6396 4380
rect 6452 4378 6476 4380
rect 6532 4378 6556 4380
rect 6612 4378 6636 4380
rect 6692 4378 6706 4380
rect 5746 4326 5756 4378
rect 5812 4326 5822 4378
rect 6066 4326 6076 4378
rect 6132 4326 6142 4378
rect 6386 4326 6396 4378
rect 6452 4326 6462 4378
rect 5502 4324 5516 4326
rect 5572 4324 5596 4326
rect 5652 4324 5676 4326
rect 5732 4324 5756 4326
rect 5812 4324 5836 4326
rect 5892 4324 5916 4326
rect 5972 4324 5996 4326
rect 6052 4324 6076 4326
rect 6132 4324 6156 4326
rect 6212 4324 6236 4326
rect 6292 4324 6316 4326
rect 6372 4324 6396 4326
rect 6452 4324 6476 4326
rect 6532 4324 6556 4326
rect 6612 4324 6636 4326
rect 6692 4324 6706 4326
rect 5502 4315 6706 4324
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 5736 3641 5764 4150
rect 6656 4026 6684 4150
rect 6748 4146 6776 4626
rect 6840 4282 6868 6054
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6932 5234 6960 5714
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6656 3998 6776 4026
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3738 6132 3878
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 5722 3632 5778 3641
rect 5722 3567 5778 3576
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5092 2910 5212 2938
rect 4908 2746 5120 2774
rect 5092 2582 5120 2746
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 4068 1284 4120 1290
rect 4068 1226 4120 1232
rect 3516 1080 3568 1086
rect 3514 1048 3516 1057
rect 3568 1048 3570 1057
rect 3514 983 3570 992
rect 3422 504 3478 513
rect 3422 439 3478 448
rect 4066 232 4122 241
rect 4172 218 4200 2314
rect 5184 2310 5212 2910
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5276 1018 5304 3334
rect 5368 3126 5396 3402
rect 5502 3292 6706 3301
rect 5502 3290 5516 3292
rect 5572 3290 5596 3292
rect 5652 3290 5676 3292
rect 5732 3290 5756 3292
rect 5812 3290 5836 3292
rect 5892 3290 5916 3292
rect 5972 3290 5996 3292
rect 6052 3290 6076 3292
rect 6132 3290 6156 3292
rect 6212 3290 6236 3292
rect 6292 3290 6316 3292
rect 6372 3290 6396 3292
rect 6452 3290 6476 3292
rect 6532 3290 6556 3292
rect 6612 3290 6636 3292
rect 6692 3290 6706 3292
rect 5746 3238 5756 3290
rect 5812 3238 5822 3290
rect 6066 3238 6076 3290
rect 6132 3238 6142 3290
rect 6386 3238 6396 3290
rect 6452 3238 6462 3290
rect 5502 3236 5516 3238
rect 5572 3236 5596 3238
rect 5652 3236 5676 3238
rect 5732 3236 5756 3238
rect 5812 3236 5836 3238
rect 5892 3236 5916 3238
rect 5972 3236 5996 3238
rect 6052 3236 6076 3238
rect 6132 3236 6156 3238
rect 6212 3236 6236 3238
rect 6292 3236 6316 3238
rect 6372 3236 6396 3238
rect 6452 3236 6476 3238
rect 6532 3236 6556 3238
rect 6612 3236 6636 3238
rect 6692 3236 6706 3238
rect 5502 3227 6706 3236
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5552 2774 5580 3130
rect 6644 2984 6696 2990
rect 6748 2972 6776 3998
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6840 3194 6868 3674
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6696 2944 6776 2972
rect 6644 2926 6696 2932
rect 6828 2916 6880 2922
rect 6828 2858 6880 2864
rect 5368 2746 5580 2774
rect 5368 2446 5396 2746
rect 6840 2650 6868 2858
rect 6932 2650 6960 4694
rect 7024 3602 7052 10390
rect 7102 10296 7158 10305
rect 7102 10231 7158 10240
rect 7116 8673 7144 10231
rect 7102 8664 7158 8673
rect 7102 8599 7158 8608
rect 7208 8378 7236 10662
rect 7300 10146 7328 10764
rect 7392 10690 7420 10950
rect 7484 10810 7512 12600
rect 7656 12582 7708 12588
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7576 11762 7604 12038
rect 7668 11937 7696 12582
rect 7760 12345 7788 15399
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7852 14414 7880 14894
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7852 13938 7880 14350
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 7944 13818 7972 17478
rect 13502 17436 14706 17445
rect 13502 17434 13516 17436
rect 13572 17434 13596 17436
rect 13652 17434 13676 17436
rect 13732 17434 13756 17436
rect 13812 17434 13836 17436
rect 13892 17434 13916 17436
rect 13972 17434 13996 17436
rect 14052 17434 14076 17436
rect 14132 17434 14156 17436
rect 14212 17434 14236 17436
rect 14292 17434 14316 17436
rect 14372 17434 14396 17436
rect 14452 17434 14476 17436
rect 14532 17434 14556 17436
rect 14612 17434 14636 17436
rect 14692 17434 14706 17436
rect 13746 17382 13756 17434
rect 13812 17382 13822 17434
rect 14066 17382 14076 17434
rect 14132 17382 14142 17434
rect 14386 17382 14396 17434
rect 14452 17382 14462 17434
rect 13502 17380 13516 17382
rect 13572 17380 13596 17382
rect 13652 17380 13676 17382
rect 13732 17380 13756 17382
rect 13812 17380 13836 17382
rect 13892 17380 13916 17382
rect 13972 17380 13996 17382
rect 14052 17380 14076 17382
rect 14132 17380 14156 17382
rect 14212 17380 14236 17382
rect 14292 17380 14316 17382
rect 14372 17380 14396 17382
rect 14452 17380 14476 17382
rect 14532 17380 14556 17382
rect 14612 17380 14636 17382
rect 14692 17380 14706 17382
rect 13502 17371 14706 17380
rect 10874 17232 10930 17241
rect 9036 17196 9088 17202
rect 10874 17167 10930 17176
rect 9036 17138 9088 17144
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8220 15434 8248 15642
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 8036 15026 8064 15302
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8036 14278 8064 14554
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7852 13790 7972 13818
rect 7852 13394 7880 13790
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7746 12336 7802 12345
rect 7746 12271 7802 12280
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7654 11928 7710 11937
rect 7654 11863 7710 11872
rect 7760 11812 7788 12106
rect 7852 11830 7880 13194
rect 7944 12850 7972 13670
rect 8036 13569 8064 14214
rect 8022 13560 8078 13569
rect 8022 13495 8078 13504
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12374 7972 12786
rect 8036 12594 8064 13330
rect 8128 12753 8156 15370
rect 8220 15094 8248 15370
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8312 14822 8340 15030
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 14006 8248 14350
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8220 13841 8248 13942
rect 8312 13870 8340 14758
rect 8300 13864 8352 13870
rect 8206 13832 8262 13841
rect 8300 13806 8352 13812
rect 8206 13767 8262 13776
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8220 13297 8248 13398
rect 8206 13288 8262 13297
rect 8206 13223 8262 13232
rect 8312 13138 8340 13806
rect 8220 13110 8340 13138
rect 8220 12782 8248 13110
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8208 12776 8260 12782
rect 8114 12744 8170 12753
rect 8208 12718 8260 12724
rect 8114 12679 8170 12688
rect 8036 12566 8156 12594
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7930 12200 7986 12209
rect 7930 12135 7986 12144
rect 7668 11784 7788 11812
rect 7840 11824 7892 11830
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7668 11665 7696 11784
rect 7840 11766 7892 11772
rect 7654 11656 7710 11665
rect 7654 11591 7710 11600
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7944 11506 7972 12135
rect 8036 11744 8064 12378
rect 8128 11937 8156 12566
rect 8220 12374 8248 12718
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8312 12220 8340 12922
rect 8220 12192 8340 12220
rect 8114 11928 8170 11937
rect 8114 11863 8170 11872
rect 8036 11716 8156 11744
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7392 10662 7512 10690
rect 7484 10588 7512 10662
rect 7392 10560 7512 10588
rect 7392 10470 7420 10560
rect 7380 10464 7432 10470
rect 7576 10418 7604 11018
rect 7380 10406 7432 10412
rect 7484 10390 7604 10418
rect 7300 10118 7420 10146
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7300 9586 7328 9998
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7300 9382 7328 9522
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7300 8498 7328 8910
rect 7392 8537 7420 10118
rect 7378 8528 7434 8537
rect 7288 8492 7340 8498
rect 7378 8463 7434 8472
rect 7288 8434 7340 8440
rect 7208 8350 7420 8378
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7886 7236 8230
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7300 7546 7328 7822
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7300 7410 7328 7482
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7300 6322 7328 6734
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7116 3058 7144 6054
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7300 5234 7328 5646
rect 7392 5370 7420 8350
rect 7484 7449 7512 10390
rect 7562 10296 7618 10305
rect 7562 10231 7618 10240
rect 7470 7440 7526 7449
rect 7470 7375 7526 7384
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7484 6254 7512 6666
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7576 5370 7604 10231
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7576 5166 7604 5306
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4146 7328 4558
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7300 4010 7328 4082
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7668 3194 7696 11494
rect 7760 11218 7788 11494
rect 7944 11478 8064 11506
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7838 10976 7894 10985
rect 7838 10911 7894 10920
rect 7852 10520 7880 10911
rect 7944 10849 7972 11222
rect 8036 11082 8064 11478
rect 8128 11121 8156 11716
rect 8220 11694 8248 12192
rect 8404 12050 8432 15506
rect 8312 12022 8432 12050
rect 8312 11812 8340 12022
rect 8312 11784 8432 11812
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 11354 8248 11630
rect 8404 11506 8432 11784
rect 8496 11665 8524 16662
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8588 15434 8616 15574
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8588 14006 8616 15370
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8482 11656 8538 11665
rect 8588 11626 8616 13670
rect 8680 12850 8708 14486
rect 8772 14414 8800 14826
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8772 14278 8800 14350
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8864 13802 8892 14894
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8758 13560 8814 13569
rect 8758 13495 8814 13504
rect 8772 13462 8800 13495
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8666 12744 8722 12753
rect 8666 12679 8722 12688
rect 8680 12442 8708 12679
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8666 12336 8722 12345
rect 8666 12271 8722 12280
rect 8482 11591 8538 11600
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8404 11478 8524 11506
rect 8390 11384 8446 11393
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 11342 8390 11370
rect 8206 11248 8262 11257
rect 8206 11183 8262 11192
rect 8114 11112 8170 11121
rect 8024 11076 8076 11082
rect 8114 11047 8170 11056
rect 8024 11018 8076 11024
rect 8116 11008 8168 11014
rect 8022 10976 8078 10985
rect 8116 10950 8168 10956
rect 8022 10911 8078 10920
rect 7930 10840 7986 10849
rect 7930 10775 7986 10784
rect 7760 10492 7880 10520
rect 7760 10305 7788 10492
rect 7932 10464 7984 10470
rect 7838 10432 7894 10441
rect 7932 10406 7984 10412
rect 7838 10367 7894 10376
rect 7746 10296 7802 10305
rect 7746 10231 7802 10240
rect 7746 10160 7802 10169
rect 7746 10095 7802 10104
rect 7760 9110 7788 10095
rect 7852 9489 7880 10367
rect 7838 9480 7894 9489
rect 7838 9415 7894 9424
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8634 7788 8910
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7746 8528 7802 8537
rect 7746 8463 7802 8472
rect 7760 7410 7788 8463
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 6458 7788 6734
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7852 5778 7880 7890
rect 7944 6730 7972 10406
rect 8036 9625 8064 10911
rect 8128 10810 8156 10950
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8220 10520 8248 11183
rect 8128 10492 8248 10520
rect 8128 10169 8156 10492
rect 8206 10432 8262 10441
rect 8206 10367 8262 10376
rect 8114 10160 8170 10169
rect 8114 10095 8170 10104
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8128 9654 8156 9930
rect 8116 9648 8168 9654
rect 8022 9616 8078 9625
rect 8116 9590 8168 9596
rect 8022 9551 8078 9560
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8036 9382 8064 9454
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8128 8566 8156 8842
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8128 7478 8156 7754
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 7944 6322 7972 6666
rect 8128 6390 8156 6666
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8036 5234 8064 5306
rect 8128 5302 8156 5578
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8220 4842 8248 10367
rect 8312 5914 8340 11342
rect 8390 11319 8446 11328
rect 8496 11268 8524 11478
rect 8404 11240 8524 11268
rect 8574 11248 8630 11257
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8024 4820 8076 4826
rect 8220 4814 8340 4842
rect 8024 4762 8076 4768
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7746 4040 7802 4049
rect 7746 3975 7802 3984
rect 7760 3466 7788 3975
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7852 3058 7880 3402
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7852 2650 7880 2994
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 5502 2204 6706 2213
rect 5502 2202 5516 2204
rect 5572 2202 5596 2204
rect 5652 2202 5676 2204
rect 5732 2202 5756 2204
rect 5812 2202 5836 2204
rect 5892 2202 5916 2204
rect 5972 2202 5996 2204
rect 6052 2202 6076 2204
rect 6132 2202 6156 2204
rect 6212 2202 6236 2204
rect 6292 2202 6316 2204
rect 6372 2202 6396 2204
rect 6452 2202 6476 2204
rect 6532 2202 6556 2204
rect 6612 2202 6636 2204
rect 6692 2202 6706 2204
rect 5746 2150 5756 2202
rect 5812 2150 5822 2202
rect 6066 2150 6076 2202
rect 6132 2150 6142 2202
rect 6386 2150 6396 2202
rect 6452 2150 6462 2202
rect 5502 2148 5516 2150
rect 5572 2148 5596 2150
rect 5652 2148 5676 2150
rect 5732 2148 5756 2150
rect 5812 2148 5836 2150
rect 5892 2148 5916 2150
rect 5972 2148 5996 2150
rect 6052 2148 6076 2150
rect 6132 2148 6156 2150
rect 6212 2148 6236 2150
rect 6292 2148 6316 2150
rect 6372 2148 6396 2150
rect 6452 2148 6476 2150
rect 6532 2148 6556 2150
rect 6612 2148 6636 2150
rect 6692 2148 6706 2150
rect 5502 2139 6706 2148
rect 7576 1698 7604 2246
rect 7944 2038 7972 4218
rect 8036 3194 8064 4762
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8128 4214 8156 4490
rect 8220 4214 8248 4626
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8312 4026 8340 4814
rect 8128 3998 8340 4026
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7932 2032 7984 2038
rect 7932 1974 7984 1980
rect 8128 1970 8156 3998
rect 8404 3194 8432 11240
rect 8574 11183 8576 11192
rect 8628 11183 8630 11192
rect 8576 11154 8628 11160
rect 8482 11112 8538 11121
rect 8482 11047 8538 11056
rect 8496 10470 8524 11047
rect 8680 10606 8708 12271
rect 8772 12050 8800 13262
rect 8864 12918 8892 13738
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8864 12170 8892 12854
rect 8956 12238 8984 14758
rect 9048 14113 9076 17138
rect 9502 16892 10706 16901
rect 9502 16890 9516 16892
rect 9572 16890 9596 16892
rect 9652 16890 9676 16892
rect 9732 16890 9756 16892
rect 9812 16890 9836 16892
rect 9892 16890 9916 16892
rect 9972 16890 9996 16892
rect 10052 16890 10076 16892
rect 10132 16890 10156 16892
rect 10212 16890 10236 16892
rect 10292 16890 10316 16892
rect 10372 16890 10396 16892
rect 10452 16890 10476 16892
rect 10532 16890 10556 16892
rect 10612 16890 10636 16892
rect 10692 16890 10706 16892
rect 9746 16838 9756 16890
rect 9812 16838 9822 16890
rect 10066 16838 10076 16890
rect 10132 16838 10142 16890
rect 10386 16838 10396 16890
rect 10452 16838 10462 16890
rect 9502 16836 9516 16838
rect 9572 16836 9596 16838
rect 9652 16836 9676 16838
rect 9732 16836 9756 16838
rect 9812 16836 9836 16838
rect 9892 16836 9916 16838
rect 9972 16836 9996 16838
rect 10052 16836 10076 16838
rect 10132 16836 10156 16838
rect 10212 16836 10236 16838
rect 10292 16836 10316 16838
rect 10372 16836 10396 16838
rect 10452 16836 10476 16838
rect 10532 16836 10556 16838
rect 10612 16836 10636 16838
rect 10692 16836 10706 16838
rect 9502 16827 10706 16836
rect 9220 16176 9272 16182
rect 9220 16118 9272 16124
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 9140 14958 9168 15982
rect 9232 15026 9260 16118
rect 9502 15804 10706 15813
rect 9502 15802 9516 15804
rect 9572 15802 9596 15804
rect 9652 15802 9676 15804
rect 9732 15802 9756 15804
rect 9812 15802 9836 15804
rect 9892 15802 9916 15804
rect 9972 15802 9996 15804
rect 10052 15802 10076 15804
rect 10132 15802 10156 15804
rect 10212 15802 10236 15804
rect 10292 15802 10316 15804
rect 10372 15802 10396 15804
rect 10452 15802 10476 15804
rect 10532 15802 10556 15804
rect 10612 15802 10636 15804
rect 10692 15802 10706 15804
rect 9746 15750 9756 15802
rect 9812 15750 9822 15802
rect 10066 15750 10076 15802
rect 10132 15750 10142 15802
rect 10386 15750 10396 15802
rect 10452 15750 10462 15802
rect 9502 15748 9516 15750
rect 9572 15748 9596 15750
rect 9652 15748 9676 15750
rect 9732 15748 9756 15750
rect 9812 15748 9836 15750
rect 9892 15748 9916 15750
rect 9972 15748 9996 15750
rect 10052 15748 10076 15750
rect 10132 15748 10156 15750
rect 10212 15748 10236 15750
rect 10292 15748 10316 15750
rect 10372 15748 10396 15750
rect 10452 15748 10476 15750
rect 10532 15748 10556 15750
rect 10612 15748 10636 15750
rect 10692 15748 10706 15750
rect 9502 15739 10706 15748
rect 9404 15496 9456 15502
rect 9324 15456 9404 15484
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9034 14104 9090 14113
rect 9034 14039 9090 14048
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 9048 12782 9076 13942
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9034 12200 9090 12209
rect 8852 12164 8904 12170
rect 9034 12135 9090 12144
rect 8852 12106 8904 12112
rect 8772 12022 8984 12050
rect 8956 11778 8984 12022
rect 8864 11750 8984 11778
rect 8864 11540 8892 11750
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8772 11512 8892 11540
rect 8956 11529 8984 11562
rect 9048 11540 9076 12135
rect 9140 11937 9168 14894
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9232 13530 9260 14350
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9232 12714 9260 13466
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9126 11928 9182 11937
rect 9126 11863 9182 11872
rect 9232 11801 9260 12378
rect 9324 11937 9352 15456
rect 9404 15438 9456 15444
rect 9402 14920 9458 14929
rect 9402 14855 9404 14864
rect 9456 14855 9458 14864
rect 9404 14826 9456 14832
rect 9502 14716 10706 14725
rect 9502 14714 9516 14716
rect 9572 14714 9596 14716
rect 9652 14714 9676 14716
rect 9732 14714 9756 14716
rect 9812 14714 9836 14716
rect 9892 14714 9916 14716
rect 9972 14714 9996 14716
rect 10052 14714 10076 14716
rect 10132 14714 10156 14716
rect 10212 14714 10236 14716
rect 10292 14714 10316 14716
rect 10372 14714 10396 14716
rect 10452 14714 10476 14716
rect 10532 14714 10556 14716
rect 10612 14714 10636 14716
rect 10692 14714 10706 14716
rect 9746 14662 9756 14714
rect 9812 14662 9822 14714
rect 10066 14662 10076 14714
rect 10132 14662 10142 14714
rect 10386 14662 10396 14714
rect 10452 14662 10462 14714
rect 9502 14660 9516 14662
rect 9572 14660 9596 14662
rect 9652 14660 9676 14662
rect 9732 14660 9756 14662
rect 9812 14660 9836 14662
rect 9892 14660 9916 14662
rect 9972 14660 9996 14662
rect 10052 14660 10076 14662
rect 10132 14660 10156 14662
rect 10212 14660 10236 14662
rect 10292 14660 10316 14662
rect 10372 14660 10396 14662
rect 10452 14660 10476 14662
rect 10532 14660 10556 14662
rect 10612 14660 10636 14662
rect 10692 14660 10706 14662
rect 9502 14651 10706 14660
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9416 12753 9444 14214
rect 10322 14104 10378 14113
rect 9496 14068 9548 14074
rect 10322 14039 10378 14048
rect 9496 14010 9548 14016
rect 9508 13938 9536 14010
rect 10336 13938 10364 14039
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 9502 13628 10706 13637
rect 9502 13626 9516 13628
rect 9572 13626 9596 13628
rect 9652 13626 9676 13628
rect 9732 13626 9756 13628
rect 9812 13626 9836 13628
rect 9892 13626 9916 13628
rect 9972 13626 9996 13628
rect 10052 13626 10076 13628
rect 10132 13626 10156 13628
rect 10212 13626 10236 13628
rect 10292 13626 10316 13628
rect 10372 13626 10396 13628
rect 10452 13626 10476 13628
rect 10532 13626 10556 13628
rect 10612 13626 10636 13628
rect 10692 13626 10706 13628
rect 9746 13574 9756 13626
rect 9812 13574 9822 13626
rect 10066 13574 10076 13626
rect 10132 13574 10142 13626
rect 10386 13574 10396 13626
rect 10452 13574 10462 13626
rect 9502 13572 9516 13574
rect 9572 13572 9596 13574
rect 9652 13572 9676 13574
rect 9732 13572 9756 13574
rect 9812 13572 9836 13574
rect 9892 13572 9916 13574
rect 9972 13572 9996 13574
rect 10052 13572 10076 13574
rect 10132 13572 10156 13574
rect 10212 13572 10236 13574
rect 10292 13572 10316 13574
rect 10372 13572 10396 13574
rect 10452 13572 10476 13574
rect 10532 13572 10556 13574
rect 10612 13572 10636 13574
rect 10692 13572 10706 13574
rect 9502 13563 10706 13572
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10416 13320 10468 13326
rect 10796 13297 10824 14350
rect 10416 13262 10468 13268
rect 10782 13288 10838 13297
rect 9600 12850 9628 13262
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9402 12744 9458 12753
rect 9402 12679 9458 12688
rect 9508 12628 9536 12786
rect 9784 12782 9812 13262
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9968 12918 9996 13126
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 9772 12776 9824 12782
rect 10152 12753 10180 13262
rect 9772 12718 9824 12724
rect 10138 12744 10194 12753
rect 10428 12714 10456 13262
rect 10782 13223 10838 13232
rect 10600 13184 10652 13190
rect 10784 13184 10836 13190
rect 10652 13144 10732 13172
rect 10600 13126 10652 13132
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10138 12679 10194 12688
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 9416 12600 9536 12628
rect 10520 12628 10548 12718
rect 10600 12640 10652 12646
rect 10520 12600 10600 12628
rect 9416 12434 9444 12600
rect 10704 12628 10732 13144
rect 10784 13126 10836 13132
rect 10796 12850 10824 13126
rect 10888 12889 10916 17167
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10874 12880 10930 12889
rect 10784 12844 10836 12850
rect 10874 12815 10930 12824
rect 10784 12786 10836 12792
rect 10876 12640 10928 12646
rect 10704 12600 10824 12628
rect 10600 12582 10652 12588
rect 9502 12540 10706 12549
rect 9502 12538 9516 12540
rect 9572 12538 9596 12540
rect 9652 12538 9676 12540
rect 9732 12538 9756 12540
rect 9812 12538 9836 12540
rect 9892 12538 9916 12540
rect 9972 12538 9996 12540
rect 10052 12538 10076 12540
rect 10132 12538 10156 12540
rect 10212 12538 10236 12540
rect 10292 12538 10316 12540
rect 10372 12538 10396 12540
rect 10452 12538 10476 12540
rect 10532 12538 10556 12540
rect 10612 12538 10636 12540
rect 10692 12538 10706 12540
rect 9746 12486 9756 12538
rect 9812 12486 9822 12538
rect 10066 12486 10076 12538
rect 10132 12486 10142 12538
rect 10386 12486 10396 12538
rect 10452 12486 10462 12538
rect 9502 12484 9516 12486
rect 9572 12484 9596 12486
rect 9652 12484 9676 12486
rect 9732 12484 9756 12486
rect 9812 12484 9836 12486
rect 9892 12484 9916 12486
rect 9972 12484 9996 12486
rect 10052 12484 10076 12486
rect 10132 12484 10156 12486
rect 10212 12484 10236 12486
rect 10292 12484 10316 12486
rect 10372 12484 10396 12486
rect 10452 12484 10476 12486
rect 10532 12484 10556 12486
rect 10612 12484 10636 12486
rect 10692 12484 10706 12486
rect 9502 12475 10706 12484
rect 10416 12436 10468 12442
rect 9416 12406 9628 12434
rect 9402 12336 9458 12345
rect 9402 12271 9404 12280
rect 9456 12271 9458 12280
rect 9404 12242 9456 12248
rect 9310 11928 9366 11937
rect 9310 11863 9366 11872
rect 9218 11792 9274 11801
rect 9402 11792 9458 11801
rect 9218 11727 9274 11736
rect 9324 11736 9402 11744
rect 9324 11716 9404 11736
rect 8942 11520 8998 11529
rect 8668 10600 8720 10606
rect 8574 10568 8630 10577
rect 8668 10542 8720 10548
rect 8574 10503 8630 10512
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8588 10248 8616 10503
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8496 10220 8616 10248
rect 8496 7002 8524 10220
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8496 3670 8524 4966
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8588 3534 8616 10066
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8404 2514 8432 3130
rect 8680 3126 8708 10406
rect 8772 3738 8800 11512
rect 9048 11512 9260 11540
rect 8942 11455 8998 11464
rect 9034 11384 9090 11393
rect 9232 11354 9260 11512
rect 9034 11319 9090 11328
rect 9128 11348 9180 11354
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8864 10985 8892 11086
rect 9048 11014 9076 11319
rect 9128 11290 9180 11296
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9140 11132 9168 11290
rect 9220 11144 9272 11150
rect 9140 11104 9220 11132
rect 8944 11008 8996 11014
rect 8850 10976 8906 10985
rect 8944 10950 8996 10956
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 8850 10911 8906 10920
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8864 7857 8892 10542
rect 8850 7848 8906 7857
rect 8850 7783 8906 7792
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8588 2650 8616 2994
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8116 1964 8168 1970
rect 8116 1906 8168 1912
rect 7564 1692 7616 1698
rect 7564 1634 7616 1640
rect 8864 1086 8892 3878
rect 8956 3505 8984 10950
rect 9034 10296 9090 10305
rect 9034 10231 9090 10240
rect 9048 8498 9076 10231
rect 9140 10130 9168 11104
rect 9220 11086 9272 11092
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 9140 9654 9168 9930
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9232 9024 9260 10746
rect 9324 10606 9352 11716
rect 9456 11727 9458 11736
rect 9404 11698 9456 11704
rect 9600 11694 9628 12406
rect 10416 12378 10468 12384
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 10322 12336 10378 12345
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9770 12200 9826 12209
rect 9692 11830 9720 12174
rect 9770 12135 9826 12144
rect 9864 12164 9916 12170
rect 9784 11830 9812 12135
rect 9864 12106 9916 12112
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9772 11824 9824 11830
rect 9876 11801 9904 12106
rect 10060 11898 10088 12310
rect 10232 12300 10284 12306
rect 10322 12271 10378 12280
rect 10232 12242 10284 12248
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9772 11766 9824 11772
rect 9862 11792 9918 11801
rect 9784 11694 9812 11766
rect 9862 11727 9918 11736
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9772 11688 9824 11694
rect 10060 11665 10088 11834
rect 10244 11665 10272 12242
rect 10336 11762 10364 12271
rect 10428 12238 10456 12378
rect 10612 12306 10640 12378
rect 10690 12336 10746 12345
rect 10600 12300 10652 12306
rect 10690 12271 10746 12280
rect 10600 12242 10652 12248
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 9772 11630 9824 11636
rect 10046 11656 10102 11665
rect 10046 11591 10102 11600
rect 10230 11656 10286 11665
rect 10230 11591 10286 11600
rect 9404 11552 9456 11558
rect 10428 11540 10456 12174
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11898 10548 12106
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10704 11762 10732 12271
rect 10796 12209 10824 12600
rect 10876 12582 10928 12588
rect 10782 12200 10838 12209
rect 10782 12135 10838 12144
rect 10888 12102 10916 12582
rect 10980 12152 11008 14214
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11072 12434 11100 12786
rect 11164 12617 11192 17002
rect 17502 16892 18706 16901
rect 17502 16890 17516 16892
rect 17572 16890 17596 16892
rect 17652 16890 17676 16892
rect 17732 16890 17756 16892
rect 17812 16890 17836 16892
rect 17892 16890 17916 16892
rect 17972 16890 17996 16892
rect 18052 16890 18076 16892
rect 18132 16890 18156 16892
rect 18212 16890 18236 16892
rect 18292 16890 18316 16892
rect 18372 16890 18396 16892
rect 18452 16890 18476 16892
rect 18532 16890 18556 16892
rect 18612 16890 18636 16892
rect 18692 16890 18706 16892
rect 17746 16838 17756 16890
rect 17812 16838 17822 16890
rect 18066 16838 18076 16890
rect 18132 16838 18142 16890
rect 18386 16838 18396 16890
rect 18452 16838 18462 16890
rect 17502 16836 17516 16838
rect 17572 16836 17596 16838
rect 17652 16836 17676 16838
rect 17732 16836 17756 16838
rect 17812 16836 17836 16838
rect 17892 16836 17916 16838
rect 17972 16836 17996 16838
rect 18052 16836 18076 16838
rect 18132 16836 18156 16838
rect 18212 16836 18236 16838
rect 18292 16836 18316 16838
rect 18372 16836 18396 16838
rect 18452 16836 18476 16838
rect 18532 16836 18556 16838
rect 18612 16836 18636 16838
rect 18692 16836 18706 16838
rect 17502 16827 18706 16836
rect 18786 16688 18842 16697
rect 18786 16623 18842 16632
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 11426 15600 11482 15609
rect 11426 15535 11482 15544
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11150 12608 11206 12617
rect 11150 12543 11206 12552
rect 11072 12406 11192 12434
rect 11164 12220 11192 12406
rect 11256 12374 11284 13262
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11348 12442 11376 12718
rect 11440 12442 11468 15535
rect 11518 15328 11574 15337
rect 11518 15263 11574 15272
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11164 12192 11376 12220
rect 10980 12124 11284 12152
rect 10876 12096 10928 12102
rect 10928 12056 11008 12084
rect 10876 12038 10928 12044
rect 10784 11824 10836 11830
rect 10782 11792 10784 11801
rect 10836 11792 10838 11801
rect 10692 11756 10744 11762
rect 10782 11727 10838 11736
rect 10692 11698 10744 11704
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10428 11512 10824 11540
rect 9404 11494 9456 11500
rect 9312 10600 9364 10606
rect 9416 10577 9444 11494
rect 9502 11452 10706 11461
rect 9502 11450 9516 11452
rect 9572 11450 9596 11452
rect 9652 11450 9676 11452
rect 9732 11450 9756 11452
rect 9812 11450 9836 11452
rect 9892 11450 9916 11452
rect 9972 11450 9996 11452
rect 10052 11450 10076 11452
rect 10132 11450 10156 11452
rect 10212 11450 10236 11452
rect 10292 11450 10316 11452
rect 10372 11450 10396 11452
rect 10452 11450 10476 11452
rect 10532 11450 10556 11452
rect 10612 11450 10636 11452
rect 10692 11450 10706 11452
rect 9746 11398 9756 11450
rect 9812 11398 9822 11450
rect 10066 11398 10076 11450
rect 10132 11398 10142 11450
rect 10386 11398 10396 11450
rect 10452 11398 10462 11450
rect 9502 11396 9516 11398
rect 9572 11396 9596 11398
rect 9652 11396 9676 11398
rect 9732 11396 9756 11398
rect 9812 11396 9836 11398
rect 9892 11396 9916 11398
rect 9972 11396 9996 11398
rect 10052 11396 10076 11398
rect 10132 11396 10156 11398
rect 10212 11396 10236 11398
rect 10292 11396 10316 11398
rect 10372 11396 10396 11398
rect 10452 11396 10476 11398
rect 10532 11396 10556 11398
rect 10612 11396 10636 11398
rect 10692 11396 10706 11398
rect 9502 11387 10706 11396
rect 9496 11348 9548 11354
rect 10796 11336 10824 11512
rect 9496 11290 9548 11296
rect 10704 11308 10824 11336
rect 9508 11082 9536 11290
rect 9954 11248 10010 11257
rect 9954 11183 9956 11192
rect 10008 11183 10010 11192
rect 10598 11248 10654 11257
rect 10704 11218 10732 11308
rect 10598 11183 10654 11192
rect 10692 11212 10744 11218
rect 9956 11154 10008 11160
rect 9864 11144 9916 11150
rect 9678 11112 9734 11121
rect 9496 11076 9548 11082
rect 9864 11086 9916 11092
rect 9678 11047 9734 11056
rect 9496 11018 9548 11024
rect 9692 10810 9720 11047
rect 9772 11008 9824 11014
rect 9876 10985 9904 11086
rect 9772 10950 9824 10956
rect 9862 10976 9918 10985
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9600 10577 9628 10678
rect 9312 10542 9364 10548
rect 9402 10568 9458 10577
rect 9324 9092 9352 10542
rect 9402 10503 9458 10512
rect 9586 10568 9642 10577
rect 9586 10503 9642 10512
rect 9784 10470 9812 10950
rect 9862 10911 9918 10920
rect 9968 10538 9996 11154
rect 10138 10568 10194 10577
rect 9956 10532 10008 10538
rect 10138 10503 10194 10512
rect 9956 10474 10008 10480
rect 10152 10470 10180 10503
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 10140 10464 10192 10470
rect 10612 10452 10640 11183
rect 10692 11154 10744 11160
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10704 10577 10732 11018
rect 10888 10606 10916 11630
rect 10980 11098 11008 12056
rect 11058 12064 11114 12073
rect 11058 11999 11114 12008
rect 11072 11218 11100 11999
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10980 11070 11100 11098
rect 10966 10976 11022 10985
rect 10966 10911 11022 10920
rect 10876 10600 10928 10606
rect 10690 10568 10746 10577
rect 10876 10542 10928 10548
rect 10690 10503 10746 10512
rect 10612 10441 10824 10452
rect 10612 10432 10838 10441
rect 10612 10424 10782 10432
rect 10140 10406 10192 10412
rect 9502 10364 10706 10373
rect 10782 10367 10838 10376
rect 9502 10362 9516 10364
rect 9572 10362 9596 10364
rect 9652 10362 9676 10364
rect 9732 10362 9756 10364
rect 9812 10362 9836 10364
rect 9892 10362 9916 10364
rect 9972 10362 9996 10364
rect 10052 10362 10076 10364
rect 10132 10362 10156 10364
rect 10212 10362 10236 10364
rect 10292 10362 10316 10364
rect 10372 10362 10396 10364
rect 10452 10362 10476 10364
rect 10532 10362 10556 10364
rect 10612 10362 10636 10364
rect 10692 10362 10706 10364
rect 9746 10310 9756 10362
rect 9812 10310 9822 10362
rect 10066 10310 10076 10362
rect 10132 10310 10142 10362
rect 10386 10310 10396 10362
rect 10452 10310 10462 10362
rect 9502 10308 9516 10310
rect 9572 10308 9596 10310
rect 9652 10308 9676 10310
rect 9732 10308 9756 10310
rect 9812 10308 9836 10310
rect 9892 10308 9916 10310
rect 9972 10308 9996 10310
rect 10052 10308 10076 10310
rect 10132 10308 10156 10310
rect 10212 10308 10236 10310
rect 10292 10308 10316 10310
rect 10372 10308 10396 10310
rect 10452 10308 10476 10310
rect 10532 10308 10556 10310
rect 10612 10308 10636 10310
rect 10692 10308 10706 10310
rect 9502 10299 10706 10308
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 9402 10160 9458 10169
rect 9402 10095 9458 10104
rect 9770 10160 9826 10169
rect 9770 10095 9826 10104
rect 9416 9160 9444 10095
rect 9784 10062 9812 10095
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 10520 9654 10548 10202
rect 10876 9988 10928 9994
rect 10876 9930 10928 9936
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10690 9480 10746 9489
rect 10690 9415 10692 9424
rect 10744 9415 10746 9424
rect 10692 9386 10744 9392
rect 9502 9276 10706 9285
rect 9502 9274 9516 9276
rect 9572 9274 9596 9276
rect 9652 9274 9676 9276
rect 9732 9274 9756 9276
rect 9812 9274 9836 9276
rect 9892 9274 9916 9276
rect 9972 9274 9996 9276
rect 10052 9274 10076 9276
rect 10132 9274 10156 9276
rect 10212 9274 10236 9276
rect 10292 9274 10316 9276
rect 10372 9274 10396 9276
rect 10452 9274 10476 9276
rect 10532 9274 10556 9276
rect 10612 9274 10636 9276
rect 10692 9274 10706 9276
rect 9746 9222 9756 9274
rect 9812 9222 9822 9274
rect 10066 9222 10076 9274
rect 10132 9222 10142 9274
rect 10386 9222 10396 9274
rect 10452 9222 10462 9274
rect 9502 9220 9516 9222
rect 9572 9220 9596 9222
rect 9652 9220 9676 9222
rect 9732 9220 9756 9222
rect 9812 9220 9836 9222
rect 9892 9220 9916 9222
rect 9972 9220 9996 9222
rect 10052 9220 10076 9222
rect 10132 9220 10156 9222
rect 10212 9220 10236 9222
rect 10292 9220 10316 9222
rect 10372 9220 10396 9222
rect 10452 9220 10476 9222
rect 10532 9220 10556 9222
rect 10612 9220 10636 9222
rect 10692 9220 10706 9222
rect 9502 9211 10706 9220
rect 9956 9172 10008 9178
rect 9416 9132 9536 9160
rect 9324 9064 9444 9092
rect 9232 8996 9352 9024
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9232 8566 9260 8774
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9232 7478 9260 7686
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 6390 9260 6598
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9140 5302 9168 5578
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9220 3664 9272 3670
rect 9126 3632 9182 3641
rect 9220 3606 9272 3612
rect 9126 3567 9182 3576
rect 8942 3496 8998 3505
rect 8942 3431 8998 3440
rect 8956 2990 8984 3431
rect 9140 3398 9168 3567
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9232 3194 9260 3606
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9048 2514 9076 2858
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 9140 2446 9168 2790
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9140 1766 9168 2382
rect 9232 2378 9260 3130
rect 9324 3058 9352 8996
rect 9416 7818 9444 9064
rect 9508 9042 9536 9132
rect 10796 9160 10824 9658
rect 9956 9114 10008 9120
rect 10704 9132 10824 9160
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9968 8430 9996 9114
rect 10704 9042 10732 9132
rect 10692 9036 10744 9042
rect 10888 9024 10916 9930
rect 10692 8978 10744 8984
rect 10796 8996 10916 9024
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9502 8188 10706 8197
rect 9502 8186 9516 8188
rect 9572 8186 9596 8188
rect 9652 8186 9676 8188
rect 9732 8186 9756 8188
rect 9812 8186 9836 8188
rect 9892 8186 9916 8188
rect 9972 8186 9996 8188
rect 10052 8186 10076 8188
rect 10132 8186 10156 8188
rect 10212 8186 10236 8188
rect 10292 8186 10316 8188
rect 10372 8186 10396 8188
rect 10452 8186 10476 8188
rect 10532 8186 10556 8188
rect 10612 8186 10636 8188
rect 10692 8186 10706 8188
rect 9746 8134 9756 8186
rect 9812 8134 9822 8186
rect 10066 8134 10076 8186
rect 10132 8134 10142 8186
rect 10386 8134 10396 8186
rect 10452 8134 10462 8186
rect 9502 8132 9516 8134
rect 9572 8132 9596 8134
rect 9652 8132 9676 8134
rect 9732 8132 9756 8134
rect 9812 8132 9836 8134
rect 9892 8132 9916 8134
rect 9972 8132 9996 8134
rect 10052 8132 10076 8134
rect 10132 8132 10156 8134
rect 10212 8132 10236 8134
rect 10292 8132 10316 8134
rect 10372 8132 10396 8134
rect 10452 8132 10476 8134
rect 10532 8132 10556 8134
rect 10612 8132 10636 8134
rect 10692 8132 10706 8134
rect 9502 8123 10706 8132
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9784 7478 9812 7822
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9968 7410 9996 7754
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9502 7100 10706 7109
rect 9502 7098 9516 7100
rect 9572 7098 9596 7100
rect 9652 7098 9676 7100
rect 9732 7098 9756 7100
rect 9812 7098 9836 7100
rect 9892 7098 9916 7100
rect 9972 7098 9996 7100
rect 10052 7098 10076 7100
rect 10132 7098 10156 7100
rect 10212 7098 10236 7100
rect 10292 7098 10316 7100
rect 10372 7098 10396 7100
rect 10452 7098 10476 7100
rect 10532 7098 10556 7100
rect 10612 7098 10636 7100
rect 10692 7098 10706 7100
rect 9746 7046 9756 7098
rect 9812 7046 9822 7098
rect 10066 7046 10076 7098
rect 10132 7046 10142 7098
rect 10386 7046 10396 7098
rect 10452 7046 10462 7098
rect 9502 7044 9516 7046
rect 9572 7044 9596 7046
rect 9652 7044 9676 7046
rect 9732 7044 9756 7046
rect 9812 7044 9836 7046
rect 9892 7044 9916 7046
rect 9972 7044 9996 7046
rect 10052 7044 10076 7046
rect 10132 7044 10156 7046
rect 10212 7044 10236 7046
rect 10292 7044 10316 7046
rect 10372 7044 10396 7046
rect 10452 7044 10476 7046
rect 10532 7044 10556 7046
rect 10612 7044 10636 7046
rect 10692 7044 10706 7046
rect 9502 7035 10706 7044
rect 9502 6012 10706 6021
rect 9502 6010 9516 6012
rect 9572 6010 9596 6012
rect 9652 6010 9676 6012
rect 9732 6010 9756 6012
rect 9812 6010 9836 6012
rect 9892 6010 9916 6012
rect 9972 6010 9996 6012
rect 10052 6010 10076 6012
rect 10132 6010 10156 6012
rect 10212 6010 10236 6012
rect 10292 6010 10316 6012
rect 10372 6010 10396 6012
rect 10452 6010 10476 6012
rect 10532 6010 10556 6012
rect 10612 6010 10636 6012
rect 10692 6010 10706 6012
rect 9746 5958 9756 6010
rect 9812 5958 9822 6010
rect 10066 5958 10076 6010
rect 10132 5958 10142 6010
rect 10386 5958 10396 6010
rect 10452 5958 10462 6010
rect 9502 5956 9516 5958
rect 9572 5956 9596 5958
rect 9652 5956 9676 5958
rect 9732 5956 9756 5958
rect 9812 5956 9836 5958
rect 9892 5956 9916 5958
rect 9972 5956 9996 5958
rect 10052 5956 10076 5958
rect 10132 5956 10156 5958
rect 10212 5956 10236 5958
rect 10292 5956 10316 5958
rect 10372 5956 10396 5958
rect 10452 5956 10476 5958
rect 10532 5956 10556 5958
rect 10612 5956 10636 5958
rect 10692 5956 10706 5958
rect 9502 5947 10706 5956
rect 9502 4924 10706 4933
rect 9502 4922 9516 4924
rect 9572 4922 9596 4924
rect 9652 4922 9676 4924
rect 9732 4922 9756 4924
rect 9812 4922 9836 4924
rect 9892 4922 9916 4924
rect 9972 4922 9996 4924
rect 10052 4922 10076 4924
rect 10132 4922 10156 4924
rect 10212 4922 10236 4924
rect 10292 4922 10316 4924
rect 10372 4922 10396 4924
rect 10452 4922 10476 4924
rect 10532 4922 10556 4924
rect 10612 4922 10636 4924
rect 10692 4922 10706 4924
rect 9746 4870 9756 4922
rect 9812 4870 9822 4922
rect 10066 4870 10076 4922
rect 10132 4870 10142 4922
rect 10386 4870 10396 4922
rect 10452 4870 10462 4922
rect 9502 4868 9516 4870
rect 9572 4868 9596 4870
rect 9652 4868 9676 4870
rect 9732 4868 9756 4870
rect 9812 4868 9836 4870
rect 9892 4868 9916 4870
rect 9972 4868 9996 4870
rect 10052 4868 10076 4870
rect 10132 4868 10156 4870
rect 10212 4868 10236 4870
rect 10292 4868 10316 4870
rect 10372 4868 10396 4870
rect 10452 4868 10476 4870
rect 10532 4868 10556 4870
rect 10612 4868 10636 4870
rect 10692 4868 10706 4870
rect 9502 4859 10706 4868
rect 10690 4584 10746 4593
rect 10690 4519 10692 4528
rect 10744 4519 10746 4528
rect 10692 4490 10744 4496
rect 9502 3836 10706 3845
rect 9502 3834 9516 3836
rect 9572 3834 9596 3836
rect 9652 3834 9676 3836
rect 9732 3834 9756 3836
rect 9812 3834 9836 3836
rect 9892 3834 9916 3836
rect 9972 3834 9996 3836
rect 10052 3834 10076 3836
rect 10132 3834 10156 3836
rect 10212 3834 10236 3836
rect 10292 3834 10316 3836
rect 10372 3834 10396 3836
rect 10452 3834 10476 3836
rect 10532 3834 10556 3836
rect 10612 3834 10636 3836
rect 10692 3834 10706 3836
rect 9746 3782 9756 3834
rect 9812 3782 9822 3834
rect 10066 3782 10076 3834
rect 10132 3782 10142 3834
rect 10386 3782 10396 3834
rect 10452 3782 10462 3834
rect 9502 3780 9516 3782
rect 9572 3780 9596 3782
rect 9652 3780 9676 3782
rect 9732 3780 9756 3782
rect 9812 3780 9836 3782
rect 9892 3780 9916 3782
rect 9972 3780 9996 3782
rect 10052 3780 10076 3782
rect 10132 3780 10156 3782
rect 10212 3780 10236 3782
rect 10292 3780 10316 3782
rect 10372 3780 10396 3782
rect 10452 3780 10476 3782
rect 10532 3780 10556 3782
rect 10612 3780 10636 3782
rect 10692 3780 10706 3782
rect 9502 3771 10706 3780
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 9416 3534 9444 3674
rect 10416 3664 10468 3670
rect 9586 3632 9642 3641
rect 10416 3606 10468 3612
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 9586 3567 9642 3576
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9324 2514 9352 2994
rect 9416 2530 9444 3470
rect 9600 3126 9628 3567
rect 10428 3369 10456 3606
rect 10520 3534 10548 3606
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10508 3392 10560 3398
rect 10414 3360 10470 3369
rect 10508 3334 10560 3340
rect 10414 3295 10470 3304
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 10520 2922 10548 3334
rect 10612 3233 10640 3470
rect 10598 3224 10654 3233
rect 10598 3159 10654 3168
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10704 2854 10732 3674
rect 10796 3058 10824 8996
rect 10980 8922 11008 10911
rect 11072 9926 11100 11070
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11072 9217 11100 9386
rect 11058 9208 11114 9217
rect 11058 9143 11114 9152
rect 11058 9072 11114 9081
rect 11058 9007 11114 9016
rect 11072 8974 11100 9007
rect 10888 8894 11008 8922
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10888 2922 10916 8894
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 9502 2748 10706 2757
rect 9502 2746 9516 2748
rect 9572 2746 9596 2748
rect 9652 2746 9676 2748
rect 9732 2746 9756 2748
rect 9812 2746 9836 2748
rect 9892 2746 9916 2748
rect 9972 2746 9996 2748
rect 10052 2746 10076 2748
rect 10132 2746 10156 2748
rect 10212 2746 10236 2748
rect 10292 2746 10316 2748
rect 10372 2746 10396 2748
rect 10452 2746 10476 2748
rect 10532 2746 10556 2748
rect 10612 2746 10636 2748
rect 10692 2746 10706 2748
rect 9746 2694 9756 2746
rect 9812 2694 9822 2746
rect 10066 2694 10076 2746
rect 10132 2694 10142 2746
rect 10386 2694 10396 2746
rect 10452 2694 10462 2746
rect 9502 2692 9516 2694
rect 9572 2692 9596 2694
rect 9652 2692 9676 2694
rect 9732 2692 9756 2694
rect 9812 2692 9836 2694
rect 9892 2692 9916 2694
rect 9972 2692 9996 2694
rect 10052 2692 10076 2694
rect 10132 2692 10156 2694
rect 10212 2692 10236 2694
rect 10292 2692 10316 2694
rect 10372 2692 10396 2694
rect 10452 2692 10476 2694
rect 10532 2692 10556 2694
rect 10612 2692 10636 2694
rect 10692 2692 10706 2694
rect 9502 2683 10706 2692
rect 9416 2514 9812 2530
rect 9312 2508 9364 2514
rect 9416 2508 9824 2514
rect 9416 2502 9772 2508
rect 9312 2450 9364 2456
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9128 1760 9180 1766
rect 9128 1702 9180 1708
rect 9600 1222 9628 2502
rect 9772 2450 9824 2456
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 2106 9720 2382
rect 10600 2372 10652 2378
rect 10600 2314 10652 2320
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 10612 1834 10640 2314
rect 10796 2310 10824 2858
rect 10874 2816 10930 2825
rect 10874 2751 10930 2760
rect 10888 2446 10916 2751
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10600 1828 10652 1834
rect 10600 1770 10652 1776
rect 10980 1358 11008 8774
rect 11072 7478 11100 8774
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11072 6905 11100 7278
rect 11164 7002 11192 11494
rect 11256 9994 11284 12124
rect 11348 10742 11376 12192
rect 11532 12186 11560 15263
rect 11702 14920 11758 14929
rect 11702 14855 11758 14864
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11440 12158 11560 12186
rect 11440 10985 11468 12158
rect 11520 12096 11572 12102
rect 11624 12084 11652 13262
rect 11716 13002 11744 14855
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11808 13938 11836 14350
rect 11980 14000 12032 14006
rect 11900 13960 11980 13988
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13394 11836 13670
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11794 13016 11850 13025
rect 11716 12974 11794 13002
rect 11794 12951 11850 12960
rect 11900 12850 11928 13960
rect 11980 13942 12032 13948
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11794 12608 11850 12617
rect 11794 12543 11850 12552
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11572 12056 11652 12084
rect 11520 12038 11572 12044
rect 11532 11150 11560 12038
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11624 11082 11652 11834
rect 11716 11801 11744 12378
rect 11702 11792 11758 11801
rect 11702 11727 11758 11736
rect 11808 11676 11836 12543
rect 11900 12238 11928 12786
rect 11992 12238 12020 13126
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11900 11830 11928 12174
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11808 11648 11928 11676
rect 11794 11350 11850 11359
rect 11794 11285 11850 11294
rect 11702 11112 11758 11121
rect 11612 11076 11664 11082
rect 11702 11047 11758 11056
rect 11612 11018 11664 11024
rect 11426 10976 11482 10985
rect 11426 10911 11482 10920
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11348 10062 11376 10678
rect 11428 10532 11480 10538
rect 11428 10474 11480 10480
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11242 9888 11298 9897
rect 11242 9823 11298 9832
rect 11256 7721 11284 9823
rect 11348 9722 11376 9998
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11334 9616 11390 9625
rect 11440 9586 11468 10474
rect 11334 9551 11390 9560
rect 11428 9580 11480 9586
rect 11242 7712 11298 7721
rect 11242 7647 11298 7656
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11256 7206 11284 7482
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11058 6896 11114 6905
rect 11058 6831 11114 6840
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11072 4049 11100 6326
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11164 5778 11192 6258
rect 11256 6254 11284 7142
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 11058 3632 11114 3641
rect 11058 3567 11114 3576
rect 11072 3369 11100 3567
rect 11058 3360 11114 3369
rect 11058 3295 11114 3304
rect 11164 3108 11192 4218
rect 11348 4026 11376 9551
rect 11428 9522 11480 9528
rect 11440 7954 11468 9522
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11426 7712 11482 7721
rect 11426 7647 11482 7656
rect 11440 6390 11468 7647
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11440 5914 11468 6190
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11532 4146 11560 10678
rect 11624 8090 11652 11018
rect 11716 10169 11744 11047
rect 11808 10713 11836 11285
rect 11900 11014 11928 11648
rect 12084 11354 12112 12854
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12070 11248 12126 11257
rect 12070 11183 12126 11192
rect 11978 11112 12034 11121
rect 11978 11047 12034 11056
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11794 10704 11850 10713
rect 11794 10639 11850 10648
rect 11794 10568 11850 10577
rect 11794 10503 11850 10512
rect 11888 10532 11940 10538
rect 11702 10160 11758 10169
rect 11702 10095 11758 10104
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11716 9722 11744 9930
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11716 8362 11744 9386
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11624 7002 11652 7346
rect 11702 7032 11758 7041
rect 11612 6996 11664 7002
rect 11702 6967 11758 6976
rect 11612 6938 11664 6944
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11624 4622 11652 5102
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11348 3998 11468 4026
rect 11336 3936 11388 3942
rect 11242 3904 11298 3913
rect 11336 3878 11388 3884
rect 11242 3839 11298 3848
rect 11256 3534 11284 3839
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11348 3380 11376 3878
rect 11440 3398 11468 3998
rect 11072 3080 11192 3108
rect 11256 3352 11376 3380
rect 11428 3392 11480 3398
rect 11072 2514 11100 3080
rect 11256 3040 11284 3352
rect 11428 3334 11480 3340
rect 11164 3012 11284 3040
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11164 2106 11192 3012
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11256 2378 11284 2858
rect 11532 2446 11560 4082
rect 11624 3602 11652 4558
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11716 2825 11744 6967
rect 11808 6746 11836 10503
rect 11888 10474 11940 10480
rect 11900 8906 11928 10474
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11808 6718 11928 6746
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 5778 11836 6598
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11900 4486 11928 6718
rect 11992 5914 12020 11047
rect 12084 10742 12112 11183
rect 12176 11150 12204 13330
rect 12268 12617 12296 16390
rect 13502 16348 14706 16357
rect 13502 16346 13516 16348
rect 13572 16346 13596 16348
rect 13652 16346 13676 16348
rect 13732 16346 13756 16348
rect 13812 16346 13836 16348
rect 13892 16346 13916 16348
rect 13972 16346 13996 16348
rect 14052 16346 14076 16348
rect 14132 16346 14156 16348
rect 14212 16346 14236 16348
rect 14292 16346 14316 16348
rect 14372 16346 14396 16348
rect 14452 16346 14476 16348
rect 14532 16346 14556 16348
rect 14612 16346 14636 16348
rect 14692 16346 14706 16348
rect 13746 16294 13756 16346
rect 13812 16294 13822 16346
rect 14066 16294 14076 16346
rect 14132 16294 14142 16346
rect 14386 16294 14396 16346
rect 14452 16294 14462 16346
rect 13502 16292 13516 16294
rect 13572 16292 13596 16294
rect 13652 16292 13676 16294
rect 13732 16292 13756 16294
rect 13812 16292 13836 16294
rect 13892 16292 13916 16294
rect 13972 16292 13996 16294
rect 14052 16292 14076 16294
rect 14132 16292 14156 16294
rect 14212 16292 14236 16294
rect 14292 16292 14316 16294
rect 14372 16292 14396 16294
rect 14452 16292 14476 16294
rect 14532 16292 14556 16294
rect 14612 16292 14636 16294
rect 14692 16292 14706 16294
rect 13502 16283 14706 16292
rect 16578 16008 16634 16017
rect 12348 15972 12400 15978
rect 16578 15943 16634 15952
rect 12348 15914 12400 15920
rect 12254 12608 12310 12617
rect 12254 12543 12310 12552
rect 12360 12481 12388 15914
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12452 13870 12480 14282
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12346 12472 12402 12481
rect 12346 12407 12402 12416
rect 12346 12200 12402 12209
rect 12346 12135 12402 12144
rect 12254 12064 12310 12073
rect 12254 11999 12310 12008
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12176 10266 12204 10542
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12162 10160 12218 10169
rect 12162 10095 12218 10104
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12084 7818 12112 9930
rect 12176 9722 12204 10095
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12268 9568 12296 11999
rect 12360 11393 12388 12135
rect 12452 12102 12480 13466
rect 12624 13456 12676 13462
rect 12728 13444 12756 13806
rect 12676 13416 12756 13444
rect 12624 13398 12676 13404
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12636 12986 12664 13262
rect 12728 13258 12756 13416
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12728 12866 12756 13194
rect 12636 12838 12756 12866
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12544 11778 12572 12242
rect 12636 12170 12664 12838
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12728 12238 12756 12718
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12452 11750 12572 11778
rect 12346 11384 12402 11393
rect 12346 11319 12402 11328
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12360 10674 12388 11222
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12452 10577 12480 11750
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12544 10674 12572 11562
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12438 10568 12494 10577
rect 12438 10503 12494 10512
rect 12438 10432 12494 10441
rect 12438 10367 12494 10376
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12176 9540 12296 9568
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12084 5710 12112 6734
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11992 5302 12020 5510
rect 12084 5370 12112 5646
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 12084 5166 12112 5306
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 12072 4140 12124 4146
rect 12176 4128 12204 9540
rect 12360 9466 12388 9590
rect 12452 9518 12480 10367
rect 12544 10062 12572 10610
rect 12636 10606 12664 12106
rect 12728 11762 12756 12174
rect 12820 11801 12848 15302
rect 13502 15260 14706 15269
rect 13502 15258 13516 15260
rect 13572 15258 13596 15260
rect 13652 15258 13676 15260
rect 13732 15258 13756 15260
rect 13812 15258 13836 15260
rect 13892 15258 13916 15260
rect 13972 15258 13996 15260
rect 14052 15258 14076 15260
rect 14132 15258 14156 15260
rect 14212 15258 14236 15260
rect 14292 15258 14316 15260
rect 14372 15258 14396 15260
rect 14452 15258 14476 15260
rect 14532 15258 14556 15260
rect 14612 15258 14636 15260
rect 14692 15258 14706 15260
rect 13746 15206 13756 15258
rect 13812 15206 13822 15258
rect 14066 15206 14076 15258
rect 14132 15206 14142 15258
rect 14386 15206 14396 15258
rect 14452 15206 14462 15258
rect 13502 15204 13516 15206
rect 13572 15204 13596 15206
rect 13652 15204 13676 15206
rect 13732 15204 13756 15206
rect 13812 15204 13836 15206
rect 13892 15204 13916 15206
rect 13972 15204 13996 15206
rect 14052 15204 14076 15206
rect 14132 15204 14156 15206
rect 14212 15204 14236 15206
rect 14292 15204 14316 15206
rect 14372 15204 14396 15206
rect 14452 15204 14476 15206
rect 14532 15204 14556 15206
rect 14612 15204 14636 15206
rect 14692 15204 14706 15206
rect 13502 15195 14706 15204
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 13176 14476 13228 14482
rect 13228 14436 13308 14464
rect 13176 14418 13228 14424
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12912 12850 12940 13874
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12806 11792 12862 11801
rect 12716 11756 12768 11762
rect 12806 11727 12862 11736
rect 12716 11698 12768 11704
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12728 11014 12756 11494
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12544 9586 12572 9998
rect 12636 9586 12664 10406
rect 12728 10010 12756 10950
rect 12820 10674 12848 11494
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12728 9982 12848 10010
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12268 9438 12388 9466
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12268 8294 12296 9438
rect 12348 9376 12400 9382
rect 12544 9364 12572 9522
rect 12348 9318 12400 9324
rect 12452 9336 12572 9364
rect 12360 9178 12388 9318
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12452 8129 12480 9336
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12438 8120 12494 8129
rect 12544 8090 12572 9114
rect 12636 8566 12664 9522
rect 12728 8673 12756 9658
rect 12820 9382 12848 9982
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12714 8664 12770 8673
rect 12820 8634 12848 9318
rect 12714 8599 12770 8608
rect 12808 8628 12860 8634
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12438 8055 12494 8064
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12636 8022 12664 8230
rect 12728 8090 12756 8599
rect 12808 8570 12860 8576
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12268 6746 12296 7414
rect 12544 6934 12572 7890
rect 12636 7274 12664 7958
rect 12820 7886 12848 8570
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12622 7168 12678 7177
rect 12622 7103 12678 7112
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12440 6792 12492 6798
rect 12438 6760 12440 6769
rect 12532 6792 12584 6798
rect 12492 6760 12494 6769
rect 12268 6718 12388 6746
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 6254 12296 6598
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12268 5302 12296 5850
rect 12360 5846 12388 6718
rect 12532 6734 12584 6740
rect 12438 6695 12494 6704
rect 12452 6254 12480 6695
rect 12544 6361 12572 6734
rect 12530 6352 12586 6361
rect 12530 6287 12532 6296
rect 12584 6287 12586 6296
rect 12532 6258 12584 6264
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12636 6118 12664 7103
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12124 4100 12204 4128
rect 12072 4082 12124 4088
rect 11702 2816 11758 2825
rect 11702 2751 11758 2760
rect 11808 2514 11836 4082
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11900 2990 11928 3946
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11992 3398 12020 3674
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 12084 3058 12112 3402
rect 12176 3194 12204 3402
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 12268 2446 12296 4014
rect 12360 3913 12388 4422
rect 12452 4214 12480 4422
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12346 3904 12402 3913
rect 12346 3839 12402 3848
rect 12360 2990 12388 3839
rect 12728 3777 12756 7686
rect 12912 5778 12940 12786
rect 13004 12782 13032 13942
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 11898 13032 12038
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13004 9654 13032 11698
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 13004 6458 13032 9114
rect 13096 7970 13124 13806
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13188 12730 13216 12922
rect 13280 12832 13308 14436
rect 13372 14346 13584 14362
rect 13372 14340 13596 14346
rect 13372 14334 13544 14340
rect 13372 14006 13400 14334
rect 13544 14282 13596 14288
rect 13502 14172 14706 14181
rect 13502 14170 13516 14172
rect 13572 14170 13596 14172
rect 13652 14170 13676 14172
rect 13732 14170 13756 14172
rect 13812 14170 13836 14172
rect 13892 14170 13916 14172
rect 13972 14170 13996 14172
rect 14052 14170 14076 14172
rect 14132 14170 14156 14172
rect 14212 14170 14236 14172
rect 14292 14170 14316 14172
rect 14372 14170 14396 14172
rect 14452 14170 14476 14172
rect 14532 14170 14556 14172
rect 14612 14170 14636 14172
rect 14692 14170 14706 14172
rect 13746 14118 13756 14170
rect 13812 14118 13822 14170
rect 14066 14118 14076 14170
rect 14132 14118 14142 14170
rect 14386 14118 14396 14170
rect 14452 14118 14462 14170
rect 13502 14116 13516 14118
rect 13572 14116 13596 14118
rect 13652 14116 13676 14118
rect 13732 14116 13756 14118
rect 13812 14116 13836 14118
rect 13892 14116 13916 14118
rect 13972 14116 13996 14118
rect 14052 14116 14076 14118
rect 14132 14116 14156 14118
rect 14212 14116 14236 14118
rect 14292 14116 14316 14118
rect 14372 14116 14396 14118
rect 14452 14116 14476 14118
rect 14532 14116 14556 14118
rect 14612 14116 14636 14118
rect 14692 14116 14706 14118
rect 13502 14107 14706 14116
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 14752 13326 14780 15030
rect 15750 14512 15806 14521
rect 15016 14476 15068 14482
rect 15750 14447 15806 14456
rect 15016 14418 15068 14424
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 12968 13400 13126
rect 13502 13084 14706 13093
rect 13502 13082 13516 13084
rect 13572 13082 13596 13084
rect 13652 13082 13676 13084
rect 13732 13082 13756 13084
rect 13812 13082 13836 13084
rect 13892 13082 13916 13084
rect 13972 13082 13996 13084
rect 14052 13082 14076 13084
rect 14132 13082 14156 13084
rect 14212 13082 14236 13084
rect 14292 13082 14316 13084
rect 14372 13082 14396 13084
rect 14452 13082 14476 13084
rect 14532 13082 14556 13084
rect 14612 13082 14636 13084
rect 14692 13082 14706 13084
rect 13746 13030 13756 13082
rect 13812 13030 13822 13082
rect 14066 13030 14076 13082
rect 14132 13030 14142 13082
rect 14386 13030 14396 13082
rect 14452 13030 14462 13082
rect 13502 13028 13516 13030
rect 13572 13028 13596 13030
rect 13652 13028 13676 13030
rect 13732 13028 13756 13030
rect 13812 13028 13836 13030
rect 13892 13028 13916 13030
rect 13972 13028 13996 13030
rect 14052 13028 14076 13030
rect 14132 13028 14156 13030
rect 14212 13028 14236 13030
rect 14292 13028 14316 13030
rect 14372 13028 14396 13030
rect 14452 13028 14476 13030
rect 14532 13028 14556 13030
rect 14612 13028 14636 13030
rect 14692 13028 14706 13030
rect 13502 13019 14706 13028
rect 13372 12940 13492 12968
rect 13280 12804 13400 12832
rect 13188 12702 13308 12730
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13188 11830 13216 12582
rect 13280 11830 13308 12702
rect 13372 12374 13400 12804
rect 13464 12714 13492 12940
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13464 12442 13492 12650
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 14384 12306 14412 12582
rect 14844 12434 14872 13942
rect 14936 13802 14964 13942
rect 14924 13796 14976 13802
rect 14924 13738 14976 13744
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14752 12406 14872 12434
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11898 13400 12038
rect 13502 11996 14706 12005
rect 13502 11994 13516 11996
rect 13572 11994 13596 11996
rect 13652 11994 13676 11996
rect 13732 11994 13756 11996
rect 13812 11994 13836 11996
rect 13892 11994 13916 11996
rect 13972 11994 13996 11996
rect 14052 11994 14076 11996
rect 14132 11994 14156 11996
rect 14212 11994 14236 11996
rect 14292 11994 14316 11996
rect 14372 11994 14396 11996
rect 14452 11994 14476 11996
rect 14532 11994 14556 11996
rect 14612 11994 14636 11996
rect 14692 11994 14706 11996
rect 13746 11942 13756 11994
rect 13812 11942 13822 11994
rect 14066 11942 14076 11994
rect 14132 11942 14142 11994
rect 14386 11942 14396 11994
rect 14452 11942 14462 11994
rect 13502 11940 13516 11942
rect 13572 11940 13596 11942
rect 13652 11940 13676 11942
rect 13732 11940 13756 11942
rect 13812 11940 13836 11942
rect 13892 11940 13916 11942
rect 13972 11940 13996 11942
rect 14052 11940 14076 11942
rect 14132 11940 14156 11942
rect 14212 11940 14236 11942
rect 14292 11940 14316 11942
rect 14372 11940 14396 11942
rect 14452 11940 14476 11942
rect 14532 11940 14556 11942
rect 14612 11940 14636 11942
rect 14692 11940 14706 11942
rect 13502 11931 14706 11940
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13188 11082 13216 11766
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13280 10010 13308 11494
rect 14292 11354 14320 11562
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14462 11248 14518 11257
rect 14462 11183 14464 11192
rect 14516 11183 14518 11192
rect 14464 11154 14516 11160
rect 14568 11082 14596 11834
rect 14646 11792 14702 11801
rect 14646 11727 14702 11736
rect 14660 11150 14688 11727
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10606 13400 10950
rect 13502 10908 14706 10917
rect 13502 10906 13516 10908
rect 13572 10906 13596 10908
rect 13652 10906 13676 10908
rect 13732 10906 13756 10908
rect 13812 10906 13836 10908
rect 13892 10906 13916 10908
rect 13972 10906 13996 10908
rect 14052 10906 14076 10908
rect 14132 10906 14156 10908
rect 14212 10906 14236 10908
rect 14292 10906 14316 10908
rect 14372 10906 14396 10908
rect 14452 10906 14476 10908
rect 14532 10906 14556 10908
rect 14612 10906 14636 10908
rect 14692 10906 14706 10908
rect 13746 10854 13756 10906
rect 13812 10854 13822 10906
rect 14066 10854 14076 10906
rect 14132 10854 14142 10906
rect 14386 10854 14396 10906
rect 14452 10854 14462 10906
rect 13502 10852 13516 10854
rect 13572 10852 13596 10854
rect 13652 10852 13676 10854
rect 13732 10852 13756 10854
rect 13812 10852 13836 10854
rect 13892 10852 13916 10854
rect 13972 10852 13996 10854
rect 14052 10852 14076 10854
rect 14132 10852 14156 10854
rect 14212 10852 14236 10854
rect 14292 10852 14316 10854
rect 14372 10852 14396 10854
rect 14452 10852 14476 10854
rect 14532 10852 14556 10854
rect 14612 10852 14636 10854
rect 14692 10852 14706 10854
rect 13502 10843 14706 10852
rect 14752 10690 14780 12406
rect 14936 12186 14964 13262
rect 15028 12850 15056 14418
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14832 12164 14884 12170
rect 14936 12158 15056 12186
rect 14832 12106 14884 12112
rect 14844 11898 14872 12106
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14660 10662 14780 10690
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13188 9982 13308 10010
rect 13188 9704 13216 9982
rect 13268 9920 13320 9926
rect 13266 9888 13268 9897
rect 13320 9888 13322 9897
rect 13266 9823 13322 9832
rect 13372 9704 13400 10406
rect 14292 10033 14320 10542
rect 14476 10169 14504 10542
rect 14660 10266 14688 10662
rect 14738 10568 14794 10577
rect 14738 10503 14794 10512
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14462 10160 14518 10169
rect 14462 10095 14518 10104
rect 14476 10062 14504 10095
rect 14464 10056 14516 10062
rect 14278 10024 14334 10033
rect 14464 9998 14516 10004
rect 14278 9959 14334 9968
rect 13502 9820 14706 9829
rect 13502 9818 13516 9820
rect 13572 9818 13596 9820
rect 13652 9818 13676 9820
rect 13732 9818 13756 9820
rect 13812 9818 13836 9820
rect 13892 9818 13916 9820
rect 13972 9818 13996 9820
rect 14052 9818 14076 9820
rect 14132 9818 14156 9820
rect 14212 9818 14236 9820
rect 14292 9818 14316 9820
rect 14372 9818 14396 9820
rect 14452 9818 14476 9820
rect 14532 9818 14556 9820
rect 14612 9818 14636 9820
rect 14692 9818 14706 9820
rect 13746 9766 13756 9818
rect 13812 9766 13822 9818
rect 14066 9766 14076 9818
rect 14132 9766 14142 9818
rect 14386 9766 14396 9818
rect 14452 9766 14462 9818
rect 13502 9764 13516 9766
rect 13572 9764 13596 9766
rect 13652 9764 13676 9766
rect 13732 9764 13756 9766
rect 13812 9764 13836 9766
rect 13892 9764 13916 9766
rect 13972 9764 13996 9766
rect 14052 9764 14076 9766
rect 14132 9764 14156 9766
rect 14212 9764 14236 9766
rect 14292 9764 14316 9766
rect 14372 9764 14396 9766
rect 14452 9764 14476 9766
rect 14532 9764 14556 9766
rect 14612 9764 14636 9766
rect 14692 9764 14706 9766
rect 13502 9755 14706 9764
rect 14752 9704 14780 10503
rect 14844 9926 14872 11562
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 13188 9676 13308 9704
rect 13372 9676 13492 9704
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 9110 13216 9386
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13174 8936 13230 8945
rect 13174 8871 13176 8880
rect 13228 8871 13230 8880
rect 13176 8842 13228 8848
rect 13174 8800 13230 8809
rect 13174 8735 13230 8744
rect 13188 8294 13216 8735
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13096 7942 13216 7970
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13096 7546 13124 7822
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13096 5778 13124 6802
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12912 5250 12940 5714
rect 12912 5222 13032 5250
rect 13004 5166 13032 5222
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13096 4690 13124 5714
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12714 3768 12770 3777
rect 12714 3703 12770 3712
rect 12990 3224 13046 3233
rect 12990 3159 13046 3168
rect 12348 2984 12400 2990
rect 12716 2984 12768 2990
rect 12348 2926 12400 2932
rect 12714 2952 12716 2961
rect 12768 2952 12770 2961
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 12256 2440 12308 2446
rect 12360 2428 12388 2926
rect 12714 2887 12770 2896
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12912 2650 12940 2858
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13004 2530 13032 3159
rect 13096 2990 13124 4626
rect 13188 4162 13216 7942
rect 13280 7342 13308 9676
rect 13358 9616 13414 9625
rect 13358 9551 13414 9560
rect 13372 8634 13400 9551
rect 13464 9110 13492 9676
rect 14568 9676 14780 9704
rect 14464 9512 14516 9518
rect 13818 9480 13874 9489
rect 13544 9444 13596 9450
rect 14464 9454 14516 9460
rect 13818 9415 13874 9424
rect 14188 9444 14240 9450
rect 13544 9386 13596 9392
rect 13556 9217 13584 9386
rect 13542 9208 13598 9217
rect 13542 9143 13598 9152
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13832 8945 13860 9415
rect 14188 9386 14240 9392
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 13818 8936 13874 8945
rect 14108 8906 14136 9318
rect 14200 8974 14228 9386
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 13818 8871 13874 8880
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 14476 8838 14504 9454
rect 14568 8945 14596 9676
rect 14646 9616 14702 9625
rect 14646 9551 14702 9560
rect 14832 9580 14884 9586
rect 14554 8936 14610 8945
rect 14660 8906 14688 9551
rect 14832 9522 14884 9528
rect 14554 8871 14610 8880
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 13502 8732 14706 8741
rect 13502 8730 13516 8732
rect 13572 8730 13596 8732
rect 13652 8730 13676 8732
rect 13732 8730 13756 8732
rect 13812 8730 13836 8732
rect 13892 8730 13916 8732
rect 13972 8730 13996 8732
rect 14052 8730 14076 8732
rect 14132 8730 14156 8732
rect 14212 8730 14236 8732
rect 14292 8730 14316 8732
rect 14372 8730 14396 8732
rect 14452 8730 14476 8732
rect 14532 8730 14556 8732
rect 14612 8730 14636 8732
rect 14692 8730 14706 8732
rect 13746 8678 13756 8730
rect 13812 8678 13822 8730
rect 14066 8678 14076 8730
rect 14132 8678 14142 8730
rect 14386 8678 14396 8730
rect 14452 8678 14462 8730
rect 13502 8676 13516 8678
rect 13572 8676 13596 8678
rect 13652 8676 13676 8678
rect 13732 8676 13756 8678
rect 13812 8676 13836 8678
rect 13892 8676 13916 8678
rect 13972 8676 13996 8678
rect 14052 8676 14076 8678
rect 14132 8676 14156 8678
rect 14212 8676 14236 8678
rect 14292 8676 14316 8678
rect 14372 8676 14396 8678
rect 14452 8676 14476 8678
rect 14532 8676 14556 8678
rect 14612 8676 14636 8678
rect 14692 8676 14706 8678
rect 13502 8667 14706 8676
rect 14844 8650 14872 9522
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 14752 8622 14872 8650
rect 14094 8528 14150 8537
rect 14094 8463 14150 8472
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13280 6254 13308 6870
rect 13372 6798 13400 8230
rect 13556 7954 13584 8366
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 14108 7750 14136 8463
rect 14556 7880 14608 7886
rect 14554 7848 14556 7857
rect 14608 7848 14610 7857
rect 14554 7783 14610 7792
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 13502 7644 14706 7653
rect 13502 7642 13516 7644
rect 13572 7642 13596 7644
rect 13652 7642 13676 7644
rect 13732 7642 13756 7644
rect 13812 7642 13836 7644
rect 13892 7642 13916 7644
rect 13972 7642 13996 7644
rect 14052 7642 14076 7644
rect 14132 7642 14156 7644
rect 14212 7642 14236 7644
rect 14292 7642 14316 7644
rect 14372 7642 14396 7644
rect 14452 7642 14476 7644
rect 14532 7642 14556 7644
rect 14612 7642 14636 7644
rect 14692 7642 14706 7644
rect 13746 7590 13756 7642
rect 13812 7590 13822 7642
rect 14066 7590 14076 7642
rect 14132 7590 14142 7642
rect 14386 7590 14396 7642
rect 14452 7590 14462 7642
rect 13502 7588 13516 7590
rect 13572 7588 13596 7590
rect 13652 7588 13676 7590
rect 13732 7588 13756 7590
rect 13812 7588 13836 7590
rect 13892 7588 13916 7590
rect 13972 7588 13996 7590
rect 14052 7588 14076 7590
rect 14132 7588 14156 7590
rect 14212 7588 14236 7590
rect 14292 7588 14316 7590
rect 14372 7588 14396 7590
rect 14452 7588 14476 7590
rect 14532 7588 14556 7590
rect 14612 7588 14636 7590
rect 14692 7588 14706 7590
rect 13502 7579 14706 7588
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14016 6934 14044 7278
rect 14752 7206 14780 8622
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14844 8401 14872 8434
rect 14830 8392 14886 8401
rect 14830 8327 14886 8336
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14004 6928 14056 6934
rect 14844 6916 14872 8230
rect 14004 6870 14056 6876
rect 14752 6888 14872 6916
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13372 6118 13400 6734
rect 13502 6556 14706 6565
rect 13502 6554 13516 6556
rect 13572 6554 13596 6556
rect 13652 6554 13676 6556
rect 13732 6554 13756 6556
rect 13812 6554 13836 6556
rect 13892 6554 13916 6556
rect 13972 6554 13996 6556
rect 14052 6554 14076 6556
rect 14132 6554 14156 6556
rect 14212 6554 14236 6556
rect 14292 6554 14316 6556
rect 14372 6554 14396 6556
rect 14452 6554 14476 6556
rect 14532 6554 14556 6556
rect 14612 6554 14636 6556
rect 14692 6554 14706 6556
rect 13746 6502 13756 6554
rect 13812 6502 13822 6554
rect 14066 6502 14076 6554
rect 14132 6502 14142 6554
rect 14386 6502 14396 6554
rect 14452 6502 14462 6554
rect 13502 6500 13516 6502
rect 13572 6500 13596 6502
rect 13652 6500 13676 6502
rect 13732 6500 13756 6502
rect 13812 6500 13836 6502
rect 13892 6500 13916 6502
rect 13972 6500 13996 6502
rect 14052 6500 14076 6502
rect 14132 6500 14156 6502
rect 14212 6500 14236 6502
rect 14292 6500 14316 6502
rect 14372 6500 14396 6502
rect 14452 6500 14476 6502
rect 14532 6500 14556 6502
rect 14612 6500 14636 6502
rect 14692 6500 14706 6502
rect 13502 6491 14706 6500
rect 14556 6384 14608 6390
rect 14554 6352 14556 6361
rect 14608 6352 14610 6361
rect 14372 6316 14424 6322
rect 14554 6287 14610 6296
rect 14372 6258 14424 6264
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 14384 5914 14412 6258
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14554 6080 14610 6089
rect 14554 6015 14610 6024
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13372 4758 13400 5646
rect 14568 5574 14596 6015
rect 14660 5642 14688 6122
rect 14752 5710 14780 6888
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 13502 5468 14706 5477
rect 13502 5466 13516 5468
rect 13572 5466 13596 5468
rect 13652 5466 13676 5468
rect 13732 5466 13756 5468
rect 13812 5466 13836 5468
rect 13892 5466 13916 5468
rect 13972 5466 13996 5468
rect 14052 5466 14076 5468
rect 14132 5466 14156 5468
rect 14212 5466 14236 5468
rect 14292 5466 14316 5468
rect 14372 5466 14396 5468
rect 14452 5466 14476 5468
rect 14532 5466 14556 5468
rect 14612 5466 14636 5468
rect 14692 5466 14706 5468
rect 13746 5414 13756 5466
rect 13812 5414 13822 5466
rect 14066 5414 14076 5466
rect 14132 5414 14142 5466
rect 14386 5414 14396 5466
rect 14452 5414 14462 5466
rect 13502 5412 13516 5414
rect 13572 5412 13596 5414
rect 13652 5412 13676 5414
rect 13732 5412 13756 5414
rect 13812 5412 13836 5414
rect 13892 5412 13916 5414
rect 13972 5412 13996 5414
rect 14052 5412 14076 5414
rect 14132 5412 14156 5414
rect 14212 5412 14236 5414
rect 14292 5412 14316 5414
rect 14372 5412 14396 5414
rect 14452 5412 14476 5414
rect 14532 5412 14556 5414
rect 14612 5412 14636 5414
rect 14692 5412 14706 5414
rect 13502 5403 14706 5412
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14292 4758 14320 5102
rect 13360 4752 13412 4758
rect 13360 4694 13412 4700
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 14568 4622 14596 5306
rect 14752 4842 14780 5510
rect 14844 5030 14872 6666
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14660 4826 14780 4842
rect 14648 4820 14780 4826
rect 14700 4814 14780 4820
rect 14648 4762 14700 4768
rect 14556 4616 14608 4622
rect 14608 4564 14780 4570
rect 14556 4558 14780 4564
rect 14568 4542 14780 4558
rect 13502 4380 14706 4389
rect 13502 4378 13516 4380
rect 13572 4378 13596 4380
rect 13652 4378 13676 4380
rect 13732 4378 13756 4380
rect 13812 4378 13836 4380
rect 13892 4378 13916 4380
rect 13972 4378 13996 4380
rect 14052 4378 14076 4380
rect 14132 4378 14156 4380
rect 14212 4378 14236 4380
rect 14292 4378 14316 4380
rect 14372 4378 14396 4380
rect 14452 4378 14476 4380
rect 14532 4378 14556 4380
rect 14612 4378 14636 4380
rect 14692 4378 14706 4380
rect 13746 4326 13756 4378
rect 13812 4326 13822 4378
rect 14066 4326 14076 4378
rect 14132 4326 14142 4378
rect 14386 4326 14396 4378
rect 14452 4326 14462 4378
rect 13502 4324 13516 4326
rect 13572 4324 13596 4326
rect 13652 4324 13676 4326
rect 13732 4324 13756 4326
rect 13812 4324 13836 4326
rect 13892 4324 13916 4326
rect 13972 4324 13996 4326
rect 14052 4324 14076 4326
rect 14132 4324 14156 4326
rect 14212 4324 14236 4326
rect 14292 4324 14316 4326
rect 14372 4324 14396 4326
rect 14452 4324 14476 4326
rect 14532 4324 14556 4326
rect 14612 4324 14636 4326
rect 14692 4324 14706 4326
rect 13502 4315 14706 4324
rect 14752 4282 14780 4542
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14832 4208 14884 4214
rect 13188 4146 13400 4162
rect 14832 4150 14884 4156
rect 13188 4140 13412 4146
rect 13188 4134 13360 4140
rect 13360 4082 13412 4088
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13188 3738 13216 4014
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13280 3058 13308 4014
rect 13372 3670 13400 4082
rect 14186 4040 14242 4049
rect 14186 3975 14242 3984
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13372 3194 13400 3606
rect 14200 3466 14228 3975
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14646 3768 14702 3777
rect 14646 3703 14702 3712
rect 14660 3670 14688 3703
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14464 3528 14516 3534
rect 14278 3496 14334 3505
rect 14188 3460 14240 3466
rect 14278 3431 14280 3440
rect 14188 3402 14240 3408
rect 14332 3431 14334 3440
rect 14462 3496 14464 3505
rect 14516 3496 14518 3505
rect 14462 3431 14518 3440
rect 14280 3402 14332 3408
rect 14660 3398 14688 3606
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 13502 3292 14706 3301
rect 13502 3290 13516 3292
rect 13572 3290 13596 3292
rect 13652 3290 13676 3292
rect 13732 3290 13756 3292
rect 13812 3290 13836 3292
rect 13892 3290 13916 3292
rect 13972 3290 13996 3292
rect 14052 3290 14076 3292
rect 14132 3290 14156 3292
rect 14212 3290 14236 3292
rect 14292 3290 14316 3292
rect 14372 3290 14396 3292
rect 14452 3290 14476 3292
rect 14532 3290 14556 3292
rect 14612 3290 14636 3292
rect 14692 3290 14706 3292
rect 13746 3238 13756 3290
rect 13812 3238 13822 3290
rect 14066 3238 14076 3290
rect 14132 3238 14142 3290
rect 14386 3238 14396 3290
rect 14452 3238 14462 3290
rect 13502 3236 13516 3238
rect 13572 3236 13596 3238
rect 13652 3236 13676 3238
rect 13732 3236 13756 3238
rect 13812 3236 13836 3238
rect 13892 3236 13916 3238
rect 13972 3236 13996 3238
rect 14052 3236 14076 3238
rect 14132 3236 14156 3238
rect 14212 3236 14236 3238
rect 14292 3236 14316 3238
rect 14372 3236 14396 3238
rect 14452 3236 14476 3238
rect 14532 3236 14556 3238
rect 14612 3236 14636 3238
rect 14692 3236 14706 3238
rect 13502 3227 14706 3236
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 14752 3126 14780 3878
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13082 2544 13138 2553
rect 13004 2502 13082 2530
rect 13082 2479 13084 2488
rect 13136 2479 13138 2488
rect 13084 2450 13136 2456
rect 12440 2440 12492 2446
rect 12360 2400 12440 2428
rect 12256 2382 12308 2388
rect 13280 2428 13308 2994
rect 13924 2650 13952 2994
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 13360 2440 13412 2446
rect 13280 2400 13360 2428
rect 12440 2382 12492 2388
rect 13360 2382 13412 2388
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 2106 12296 2246
rect 13502 2204 14706 2213
rect 13502 2202 13516 2204
rect 13572 2202 13596 2204
rect 13652 2202 13676 2204
rect 13732 2202 13756 2204
rect 13812 2202 13836 2204
rect 13892 2202 13916 2204
rect 13972 2202 13996 2204
rect 14052 2202 14076 2204
rect 14132 2202 14156 2204
rect 14212 2202 14236 2204
rect 14292 2202 14316 2204
rect 14372 2202 14396 2204
rect 14452 2202 14476 2204
rect 14532 2202 14556 2204
rect 14612 2202 14636 2204
rect 14692 2202 14706 2204
rect 13746 2150 13756 2202
rect 13812 2150 13822 2202
rect 14066 2150 14076 2202
rect 14132 2150 14142 2202
rect 14386 2150 14396 2202
rect 14452 2150 14462 2202
rect 13502 2148 13516 2150
rect 13572 2148 13596 2150
rect 13652 2148 13676 2150
rect 13732 2148 13756 2150
rect 13812 2148 13836 2150
rect 13892 2148 13916 2150
rect 13972 2148 13996 2150
rect 14052 2148 14076 2150
rect 14132 2148 14156 2150
rect 14212 2148 14236 2150
rect 14292 2148 14316 2150
rect 14372 2148 14396 2150
rect 14452 2148 14476 2150
rect 14532 2148 14556 2150
rect 14612 2148 14636 2150
rect 14692 2148 14706 2150
rect 13502 2139 14706 2148
rect 14844 2106 14872 4150
rect 14936 2446 14964 12038
rect 15028 10470 15056 12158
rect 15120 11257 15148 13330
rect 15212 12238 15240 14010
rect 15304 13394 15332 14350
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15304 12850 15332 13330
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15396 12102 15424 13126
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15106 11248 15162 11257
rect 15106 11183 15162 11192
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15028 8634 15056 10066
rect 15120 9722 15148 11086
rect 15212 11082 15240 11630
rect 15290 11248 15346 11257
rect 15290 11183 15346 11192
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15212 10742 15240 11018
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15304 10010 15332 11183
rect 15396 11150 15424 11766
rect 15488 11762 15516 12854
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15396 10674 15424 11086
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15396 10130 15424 10610
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15120 8362 15148 9114
rect 15212 9042 15240 9998
rect 15304 9982 15424 10010
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15212 8430 15240 8978
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 15304 8242 15332 9862
rect 15396 8294 15424 9982
rect 15028 8214 15332 8242
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15028 6458 15056 8214
rect 15382 8120 15438 8129
rect 15382 8055 15438 8064
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15304 6866 15332 7822
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15198 6760 15254 6769
rect 15198 6695 15254 6704
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15028 4214 15056 6054
rect 15120 5778 15148 6326
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15120 4622 15148 5714
rect 15212 5710 15240 6695
rect 15304 5778 15332 6802
rect 15396 6458 15424 8055
rect 15488 7041 15516 11290
rect 15474 7032 15530 7041
rect 15474 6967 15530 6976
rect 15580 6730 15608 11562
rect 15672 11354 15700 12106
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15672 8974 15700 10474
rect 15764 9625 15792 14447
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15750 9616 15806 9625
rect 15750 9551 15806 9560
rect 15752 9512 15804 9518
rect 15750 9480 15752 9489
rect 15804 9480 15806 9489
rect 15750 9415 15806 9424
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15672 6610 15700 8570
rect 15580 6582 15700 6610
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15580 6361 15608 6582
rect 15566 6352 15622 6361
rect 15384 6316 15436 6322
rect 15566 6287 15622 6296
rect 15660 6316 15712 6322
rect 15384 6258 15436 6264
rect 15660 6258 15712 6264
rect 15396 6089 15424 6258
rect 15382 6080 15438 6089
rect 15382 6015 15438 6024
rect 15292 5772 15344 5778
rect 15344 5732 15424 5760
rect 15292 5714 15344 5720
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15304 4690 15332 4966
rect 15396 4690 15424 5732
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15488 5166 15516 5578
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15672 4690 15700 6258
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15028 3942 15056 4014
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 15028 2650 15056 3878
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15120 2825 15148 3606
rect 15212 2854 15240 4014
rect 15396 3534 15424 4626
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15580 4078 15608 4490
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 3194 15424 3470
rect 15764 3466 15792 9318
rect 15856 7954 15884 11562
rect 15948 9926 15976 13194
rect 16224 12850 16252 13330
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16028 12368 16080 12374
rect 16028 12310 16080 12316
rect 16040 10577 16068 12310
rect 16224 12238 16252 12786
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16026 10568 16082 10577
rect 16026 10503 16082 10512
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15856 5370 15884 6870
rect 15948 6322 15976 9862
rect 16040 6769 16068 10406
rect 16026 6760 16082 6769
rect 16026 6695 16082 6704
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16040 6322 16068 6598
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16040 5778 16068 6258
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 16132 5642 16160 12038
rect 16224 11762 16252 12174
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16224 9586 16252 10610
rect 16316 10470 16344 13670
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16408 12918 16436 13262
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16408 12238 16436 12854
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16592 12170 16620 15943
rect 17502 15804 18706 15813
rect 17502 15802 17516 15804
rect 17572 15802 17596 15804
rect 17652 15802 17676 15804
rect 17732 15802 17756 15804
rect 17812 15802 17836 15804
rect 17892 15802 17916 15804
rect 17972 15802 17996 15804
rect 18052 15802 18076 15804
rect 18132 15802 18156 15804
rect 18212 15802 18236 15804
rect 18292 15802 18316 15804
rect 18372 15802 18396 15804
rect 18452 15802 18476 15804
rect 18532 15802 18556 15804
rect 18612 15802 18636 15804
rect 18692 15802 18706 15804
rect 17746 15750 17756 15802
rect 17812 15750 17822 15802
rect 18066 15750 18076 15802
rect 18132 15750 18142 15802
rect 18386 15750 18396 15802
rect 18452 15750 18462 15802
rect 17502 15748 17516 15750
rect 17572 15748 17596 15750
rect 17652 15748 17676 15750
rect 17732 15748 17756 15750
rect 17812 15748 17836 15750
rect 17892 15748 17916 15750
rect 17972 15748 17996 15750
rect 18052 15748 18076 15750
rect 18132 15748 18156 15750
rect 18212 15748 18236 15750
rect 18292 15748 18316 15750
rect 18372 15748 18396 15750
rect 18452 15748 18476 15750
rect 18532 15748 18556 15750
rect 18612 15748 18636 15750
rect 18692 15748 18706 15750
rect 17502 15739 18706 15748
rect 17502 14716 18706 14725
rect 17502 14714 17516 14716
rect 17572 14714 17596 14716
rect 17652 14714 17676 14716
rect 17732 14714 17756 14716
rect 17812 14714 17836 14716
rect 17892 14714 17916 14716
rect 17972 14714 17996 14716
rect 18052 14714 18076 14716
rect 18132 14714 18156 14716
rect 18212 14714 18236 14716
rect 18292 14714 18316 14716
rect 18372 14714 18396 14716
rect 18452 14714 18476 14716
rect 18532 14714 18556 14716
rect 18612 14714 18636 14716
rect 18692 14714 18706 14716
rect 17746 14662 17756 14714
rect 17812 14662 17822 14714
rect 18066 14662 18076 14714
rect 18132 14662 18142 14714
rect 18386 14662 18396 14714
rect 18452 14662 18462 14714
rect 17502 14660 17516 14662
rect 17572 14660 17596 14662
rect 17652 14660 17676 14662
rect 17732 14660 17756 14662
rect 17812 14660 17836 14662
rect 17892 14660 17916 14662
rect 17972 14660 17996 14662
rect 18052 14660 18076 14662
rect 18132 14660 18156 14662
rect 18212 14660 18236 14662
rect 18292 14660 18316 14662
rect 18372 14660 18396 14662
rect 18452 14660 18476 14662
rect 18532 14660 18556 14662
rect 18612 14660 18636 14662
rect 18692 14660 18706 14662
rect 17502 14651 18706 14660
rect 17502 13628 18706 13637
rect 17502 13626 17516 13628
rect 17572 13626 17596 13628
rect 17652 13626 17676 13628
rect 17732 13626 17756 13628
rect 17812 13626 17836 13628
rect 17892 13626 17916 13628
rect 17972 13626 17996 13628
rect 18052 13626 18076 13628
rect 18132 13626 18156 13628
rect 18212 13626 18236 13628
rect 18292 13626 18316 13628
rect 18372 13626 18396 13628
rect 18452 13626 18476 13628
rect 18532 13626 18556 13628
rect 18612 13626 18636 13628
rect 18692 13626 18706 13628
rect 17746 13574 17756 13626
rect 17812 13574 17822 13626
rect 18066 13574 18076 13626
rect 18132 13574 18142 13626
rect 18386 13574 18396 13626
rect 18452 13574 18462 13626
rect 17502 13572 17516 13574
rect 17572 13572 17596 13574
rect 17652 13572 17676 13574
rect 17732 13572 17756 13574
rect 17812 13572 17836 13574
rect 17892 13572 17916 13574
rect 17972 13572 17996 13574
rect 18052 13572 18076 13574
rect 18132 13572 18156 13574
rect 18212 13572 18236 13574
rect 18292 13572 18316 13574
rect 18372 13572 18396 13574
rect 18452 13572 18476 13574
rect 18532 13572 18556 13574
rect 18612 13572 18636 13574
rect 18692 13572 18706 13574
rect 17502 13563 18706 13572
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 12850 17172 13262
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16210 9344 16266 9353
rect 16210 9279 16266 9288
rect 16224 7177 16252 9279
rect 16210 7168 16266 7177
rect 16210 7103 16266 7112
rect 16316 6934 16344 10202
rect 16408 9926 16436 10610
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16408 8906 16436 9454
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16408 8634 16436 8842
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16224 6390 16252 6802
rect 16408 6780 16436 8298
rect 16500 7478 16528 11630
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16316 6752 16436 6780
rect 16486 6760 16542 6769
rect 16212 6384 16264 6390
rect 16212 6326 16264 6332
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15752 3460 15804 3466
rect 15752 3402 15804 3408
rect 15580 3194 15608 3402
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15200 2848 15252 2854
rect 15106 2816 15162 2825
rect 15200 2790 15252 2796
rect 15106 2751 15162 2760
rect 15016 2644 15068 2650
rect 15016 2586 15068 2592
rect 15396 2514 15424 3130
rect 15856 3040 15884 5306
rect 16316 4826 16344 6752
rect 16486 6695 16542 6704
rect 16394 5536 16450 5545
rect 16394 5471 16450 5480
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16408 3126 16436 5471
rect 16500 5234 16528 6695
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16592 5098 16620 11494
rect 16670 10976 16726 10985
rect 16670 10911 16726 10920
rect 16684 9586 16712 10911
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16684 8974 16712 9386
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16684 8566 16712 8774
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 5370 16712 8230
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16592 4486 16620 5034
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16684 3641 16712 4626
rect 16776 4622 16804 12106
rect 16868 11257 16896 12718
rect 17144 12238 17172 12786
rect 17502 12540 18706 12549
rect 17502 12538 17516 12540
rect 17572 12538 17596 12540
rect 17652 12538 17676 12540
rect 17732 12538 17756 12540
rect 17812 12538 17836 12540
rect 17892 12538 17916 12540
rect 17972 12538 17996 12540
rect 18052 12538 18076 12540
rect 18132 12538 18156 12540
rect 18212 12538 18236 12540
rect 18292 12538 18316 12540
rect 18372 12538 18396 12540
rect 18452 12538 18476 12540
rect 18532 12538 18556 12540
rect 18612 12538 18636 12540
rect 18692 12538 18706 12540
rect 17746 12486 17756 12538
rect 17812 12486 17822 12538
rect 18066 12486 18076 12538
rect 18132 12486 18142 12538
rect 18386 12486 18396 12538
rect 18452 12486 18462 12538
rect 17502 12484 17516 12486
rect 17572 12484 17596 12486
rect 17652 12484 17676 12486
rect 17732 12484 17756 12486
rect 17812 12484 17836 12486
rect 17892 12484 17916 12486
rect 17972 12484 17996 12486
rect 18052 12484 18076 12486
rect 18132 12484 18156 12486
rect 18212 12484 18236 12486
rect 18292 12484 18316 12486
rect 18372 12484 18396 12486
rect 18452 12484 18476 12486
rect 18532 12484 18556 12486
rect 18612 12484 18636 12486
rect 18692 12484 18706 12486
rect 17502 12475 18706 12484
rect 18800 12434 18828 16623
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18984 12434 19012 14214
rect 18708 12406 18828 12434
rect 18892 12406 19012 12434
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 16960 11762 16988 12174
rect 17144 11762 17172 12174
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16854 11248 16910 11257
rect 16854 11183 16910 11192
rect 16960 11150 16988 11698
rect 17144 11218 17172 11698
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 16868 7818 16896 11018
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16960 9874 16988 10542
rect 17052 9994 17080 11018
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10266 17172 10950
rect 17236 10606 17264 12242
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17236 10198 17264 10406
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 16960 9846 17080 9874
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16960 6440 16988 9454
rect 17052 9450 17080 9846
rect 17040 9444 17092 9450
rect 17040 9386 17092 9392
rect 17052 9058 17080 9386
rect 17144 9178 17172 10066
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17052 9030 17172 9058
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 17052 7954 17080 8842
rect 17144 8294 17172 9030
rect 17236 8974 17264 9862
rect 17328 9654 17356 12106
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17420 10606 17448 11698
rect 17880 11558 17908 12106
rect 18708 11665 18736 12406
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18694 11656 18750 11665
rect 18694 11591 18750 11600
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17502 11452 18706 11461
rect 17502 11450 17516 11452
rect 17572 11450 17596 11452
rect 17652 11450 17676 11452
rect 17732 11450 17756 11452
rect 17812 11450 17836 11452
rect 17892 11450 17916 11452
rect 17972 11450 17996 11452
rect 18052 11450 18076 11452
rect 18132 11450 18156 11452
rect 18212 11450 18236 11452
rect 18292 11450 18316 11452
rect 18372 11450 18396 11452
rect 18452 11450 18476 11452
rect 18532 11450 18556 11452
rect 18612 11450 18636 11452
rect 18692 11450 18706 11452
rect 17746 11398 17756 11450
rect 17812 11398 17822 11450
rect 18066 11398 18076 11450
rect 18132 11398 18142 11450
rect 18386 11398 18396 11450
rect 18452 11398 18462 11450
rect 17502 11396 17516 11398
rect 17572 11396 17596 11398
rect 17652 11396 17676 11398
rect 17732 11396 17756 11398
rect 17812 11396 17836 11398
rect 17892 11396 17916 11398
rect 17972 11396 17996 11398
rect 18052 11396 18076 11398
rect 18132 11396 18156 11398
rect 18212 11396 18236 11398
rect 18292 11396 18316 11398
rect 18372 11396 18396 11398
rect 18452 11396 18476 11398
rect 18532 11396 18556 11398
rect 18612 11396 18636 11398
rect 18692 11396 18706 11398
rect 17502 11387 18706 11396
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17420 9994 17448 10542
rect 17502 10364 18706 10373
rect 17502 10362 17516 10364
rect 17572 10362 17596 10364
rect 17652 10362 17676 10364
rect 17732 10362 17756 10364
rect 17812 10362 17836 10364
rect 17892 10362 17916 10364
rect 17972 10362 17996 10364
rect 18052 10362 18076 10364
rect 18132 10362 18156 10364
rect 18212 10362 18236 10364
rect 18292 10362 18316 10364
rect 18372 10362 18396 10364
rect 18452 10362 18476 10364
rect 18532 10362 18556 10364
rect 18612 10362 18636 10364
rect 18692 10362 18706 10364
rect 17746 10310 17756 10362
rect 17812 10310 17822 10362
rect 18066 10310 18076 10362
rect 18132 10310 18142 10362
rect 18386 10310 18396 10362
rect 18452 10310 18462 10362
rect 17502 10308 17516 10310
rect 17572 10308 17596 10310
rect 17652 10308 17676 10310
rect 17732 10308 17756 10310
rect 17812 10308 17836 10310
rect 17892 10308 17916 10310
rect 17972 10308 17996 10310
rect 18052 10308 18076 10310
rect 18132 10308 18156 10310
rect 18212 10308 18236 10310
rect 18292 10308 18316 10310
rect 18372 10308 18396 10310
rect 18452 10308 18476 10310
rect 18532 10308 18556 10310
rect 18612 10308 18636 10310
rect 18692 10308 18706 10310
rect 17502 10299 18706 10308
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17512 9586 17540 10202
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17500 9580 17552 9586
rect 17420 9540 17500 9568
rect 17420 9160 17448 9540
rect 17500 9522 17552 9528
rect 17958 9480 18014 9489
rect 17958 9415 17960 9424
rect 18012 9415 18014 9424
rect 17960 9386 18012 9392
rect 18064 9382 18092 9862
rect 18708 9489 18736 10134
rect 18800 10130 18828 12106
rect 18892 10713 18920 12406
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 18878 10704 18934 10713
rect 18878 10639 18934 10648
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18788 9988 18840 9994
rect 18788 9930 18840 9936
rect 18694 9480 18750 9489
rect 18694 9415 18750 9424
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17502 9276 18706 9285
rect 17502 9274 17516 9276
rect 17572 9274 17596 9276
rect 17652 9274 17676 9276
rect 17732 9274 17756 9276
rect 17812 9274 17836 9276
rect 17892 9274 17916 9276
rect 17972 9274 17996 9276
rect 18052 9274 18076 9276
rect 18132 9274 18156 9276
rect 18212 9274 18236 9276
rect 18292 9274 18316 9276
rect 18372 9274 18396 9276
rect 18452 9274 18476 9276
rect 18532 9274 18556 9276
rect 18612 9274 18636 9276
rect 18692 9274 18706 9276
rect 17746 9222 17756 9274
rect 17812 9222 17822 9274
rect 18066 9222 18076 9274
rect 18132 9222 18142 9274
rect 18386 9222 18396 9274
rect 18452 9222 18462 9274
rect 17502 9220 17516 9222
rect 17572 9220 17596 9222
rect 17652 9220 17676 9222
rect 17732 9220 17756 9222
rect 17812 9220 17836 9222
rect 17892 9220 17916 9222
rect 17972 9220 17996 9222
rect 18052 9220 18076 9222
rect 18132 9220 18156 9222
rect 18212 9220 18236 9222
rect 18292 9220 18316 9222
rect 18372 9220 18396 9222
rect 18452 9220 18476 9222
rect 18532 9220 18556 9222
rect 18612 9220 18636 9222
rect 18692 9220 18706 9222
rect 17502 9211 18706 9220
rect 17420 9132 17540 9160
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 16868 6412 16988 6440
rect 16868 6089 16896 6412
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 16948 6112 17000 6118
rect 16854 6080 16910 6089
rect 16948 6054 17000 6060
rect 16854 6015 16910 6024
rect 16868 5216 16896 6015
rect 16960 5574 16988 6054
rect 17052 5914 17080 6122
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 17040 5228 17092 5234
rect 16868 5188 17040 5216
rect 16868 4826 16896 5188
rect 17040 5170 17092 5176
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16868 4146 16896 4762
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16670 3632 16726 3641
rect 16670 3567 16726 3576
rect 16960 3534 16988 3946
rect 17052 3602 17080 4150
rect 17144 4010 17172 8026
rect 17236 7478 17264 8910
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17328 8090 17356 8570
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17420 7206 17448 8434
rect 17512 8362 17540 9132
rect 18142 9072 18198 9081
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 18052 9036 18104 9042
rect 18142 9007 18198 9016
rect 18052 8978 18104 8984
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 8566 17632 8910
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17696 8294 17724 8978
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17972 8634 18000 8910
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18064 8498 18092 8978
rect 18156 8634 18184 9007
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18800 8498 18828 9930
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17502 8188 18706 8197
rect 17502 8186 17516 8188
rect 17572 8186 17596 8188
rect 17652 8186 17676 8188
rect 17732 8186 17756 8188
rect 17812 8186 17836 8188
rect 17892 8186 17916 8188
rect 17972 8186 17996 8188
rect 18052 8186 18076 8188
rect 18132 8186 18156 8188
rect 18212 8186 18236 8188
rect 18292 8186 18316 8188
rect 18372 8186 18396 8188
rect 18452 8186 18476 8188
rect 18532 8186 18556 8188
rect 18612 8186 18636 8188
rect 18692 8186 18706 8188
rect 17746 8134 17756 8186
rect 17812 8134 17822 8186
rect 18066 8134 18076 8186
rect 18132 8134 18142 8186
rect 18386 8134 18396 8186
rect 18452 8134 18462 8186
rect 17502 8132 17516 8134
rect 17572 8132 17596 8134
rect 17652 8132 17676 8134
rect 17732 8132 17756 8134
rect 17812 8132 17836 8134
rect 17892 8132 17916 8134
rect 17972 8132 17996 8134
rect 18052 8132 18076 8134
rect 18132 8132 18156 8134
rect 18212 8132 18236 8134
rect 18292 8132 18316 8134
rect 18372 8132 18396 8134
rect 18452 8132 18476 8134
rect 18532 8132 18556 8134
rect 18612 8132 18636 8134
rect 18692 8132 18706 8134
rect 17502 8123 18706 8132
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7546 18000 7686
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17502 7100 18706 7109
rect 17502 7098 17516 7100
rect 17572 7098 17596 7100
rect 17652 7098 17676 7100
rect 17732 7098 17756 7100
rect 17812 7098 17836 7100
rect 17892 7098 17916 7100
rect 17972 7098 17996 7100
rect 18052 7098 18076 7100
rect 18132 7098 18156 7100
rect 18212 7098 18236 7100
rect 18292 7098 18316 7100
rect 18372 7098 18396 7100
rect 18452 7098 18476 7100
rect 18532 7098 18556 7100
rect 18612 7098 18636 7100
rect 18692 7098 18706 7100
rect 17746 7046 17756 7098
rect 17812 7046 17822 7098
rect 18066 7046 18076 7098
rect 18132 7046 18142 7098
rect 18386 7046 18396 7098
rect 18452 7046 18462 7098
rect 17502 7044 17516 7046
rect 17572 7044 17596 7046
rect 17652 7044 17676 7046
rect 17732 7044 17756 7046
rect 17812 7044 17836 7046
rect 17892 7044 17916 7046
rect 17972 7044 17996 7046
rect 18052 7044 18076 7046
rect 18132 7044 18156 7046
rect 18212 7044 18236 7046
rect 18292 7044 18316 7046
rect 18372 7044 18396 7046
rect 18452 7044 18476 7046
rect 18532 7044 18556 7046
rect 18612 7044 18636 7046
rect 18692 7044 18706 7046
rect 17502 7035 18706 7044
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17236 5914 17264 6394
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17420 5846 17448 6938
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17788 6322 17816 6734
rect 18800 6390 18828 8434
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 18786 6216 18842 6225
rect 18786 6151 18842 6160
rect 17502 6012 18706 6021
rect 17502 6010 17516 6012
rect 17572 6010 17596 6012
rect 17652 6010 17676 6012
rect 17732 6010 17756 6012
rect 17812 6010 17836 6012
rect 17892 6010 17916 6012
rect 17972 6010 17996 6012
rect 18052 6010 18076 6012
rect 18132 6010 18156 6012
rect 18212 6010 18236 6012
rect 18292 6010 18316 6012
rect 18372 6010 18396 6012
rect 18452 6010 18476 6012
rect 18532 6010 18556 6012
rect 18612 6010 18636 6012
rect 18692 6010 18706 6012
rect 17746 5958 17756 6010
rect 17812 5958 17822 6010
rect 18066 5958 18076 6010
rect 18132 5958 18142 6010
rect 18386 5958 18396 6010
rect 18452 5958 18462 6010
rect 17502 5956 17516 5958
rect 17572 5956 17596 5958
rect 17652 5956 17676 5958
rect 17732 5956 17756 5958
rect 17812 5956 17836 5958
rect 17892 5956 17916 5958
rect 17972 5956 17996 5958
rect 18052 5956 18076 5958
rect 18132 5956 18156 5958
rect 18212 5956 18236 5958
rect 18292 5956 18316 5958
rect 18372 5956 18396 5958
rect 18452 5956 18476 5958
rect 18532 5956 18556 5958
rect 18612 5956 18636 5958
rect 18692 5956 18706 5958
rect 17502 5947 18706 5956
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 18050 5808 18106 5817
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17236 5030 17264 5306
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17236 4214 17264 4966
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 17328 4146 17356 5102
rect 17420 4758 17448 5782
rect 18050 5743 18106 5752
rect 17868 5296 17920 5302
rect 17868 5238 17920 5244
rect 17880 5030 17908 5238
rect 18064 5166 18092 5743
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18064 5030 18092 5102
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17502 4924 18706 4933
rect 17502 4922 17516 4924
rect 17572 4922 17596 4924
rect 17652 4922 17676 4924
rect 17732 4922 17756 4924
rect 17812 4922 17836 4924
rect 17892 4922 17916 4924
rect 17972 4922 17996 4924
rect 18052 4922 18076 4924
rect 18132 4922 18156 4924
rect 18212 4922 18236 4924
rect 18292 4922 18316 4924
rect 18372 4922 18396 4924
rect 18452 4922 18476 4924
rect 18532 4922 18556 4924
rect 18612 4922 18636 4924
rect 18692 4922 18706 4924
rect 17746 4870 17756 4922
rect 17812 4870 17822 4922
rect 18066 4870 18076 4922
rect 18132 4870 18142 4922
rect 18386 4870 18396 4922
rect 18452 4870 18462 4922
rect 17502 4868 17516 4870
rect 17572 4868 17596 4870
rect 17652 4868 17676 4870
rect 17732 4868 17756 4870
rect 17812 4868 17836 4870
rect 17892 4868 17916 4870
rect 17972 4868 17996 4870
rect 18052 4868 18076 4870
rect 18132 4868 18156 4870
rect 18212 4868 18236 4870
rect 18292 4868 18316 4870
rect 18372 4868 18396 4870
rect 18452 4868 18476 4870
rect 18532 4868 18556 4870
rect 18612 4868 18636 4870
rect 18692 4868 18706 4870
rect 17502 4859 18706 4868
rect 17408 4752 17460 4758
rect 18800 4706 18828 6151
rect 17408 4694 17460 4700
rect 18708 4678 18828 4706
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 17328 3942 17356 4082
rect 18708 4049 18736 4678
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 18694 4040 18750 4049
rect 18694 3975 18750 3984
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17502 3836 18706 3845
rect 17502 3834 17516 3836
rect 17572 3834 17596 3836
rect 17652 3834 17676 3836
rect 17732 3834 17756 3836
rect 17812 3834 17836 3836
rect 17892 3834 17916 3836
rect 17972 3834 17996 3836
rect 18052 3834 18076 3836
rect 18132 3834 18156 3836
rect 18212 3834 18236 3836
rect 18292 3834 18316 3836
rect 18372 3834 18396 3836
rect 18452 3834 18476 3836
rect 18532 3834 18556 3836
rect 18612 3834 18636 3836
rect 18692 3834 18706 3836
rect 17746 3782 17756 3834
rect 17812 3782 17822 3834
rect 18066 3782 18076 3834
rect 18132 3782 18142 3834
rect 18386 3782 18396 3834
rect 18452 3782 18462 3834
rect 17502 3780 17516 3782
rect 17572 3780 17596 3782
rect 17652 3780 17676 3782
rect 17732 3780 17756 3782
rect 17812 3780 17836 3782
rect 17892 3780 17916 3782
rect 17972 3780 17996 3782
rect 18052 3780 18076 3782
rect 18132 3780 18156 3782
rect 18212 3780 18236 3782
rect 18292 3780 18316 3782
rect 18372 3780 18396 3782
rect 18452 3780 18476 3782
rect 18532 3780 18556 3782
rect 18612 3780 18636 3782
rect 18692 3780 18706 3782
rect 17502 3771 18706 3780
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 17038 3496 17094 3505
rect 17038 3431 17094 3440
rect 17052 3194 17080 3431
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16396 3120 16448 3126
rect 16396 3062 16448 3068
rect 16028 3052 16080 3058
rect 15856 3012 16028 3040
rect 16028 2994 16080 3000
rect 16670 2816 16726 2825
rect 16670 2751 16726 2760
rect 16684 2514 16712 2751
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15028 2106 15056 2450
rect 16868 2446 16896 3130
rect 17052 2990 17080 3130
rect 17236 3058 17264 3334
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 17144 2514 17172 2858
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17328 2310 17356 3538
rect 17502 2748 18706 2757
rect 17502 2746 17516 2748
rect 17572 2746 17596 2748
rect 17652 2746 17676 2748
rect 17732 2746 17756 2748
rect 17812 2746 17836 2748
rect 17892 2746 17916 2748
rect 17972 2746 17996 2748
rect 18052 2746 18076 2748
rect 18132 2746 18156 2748
rect 18212 2746 18236 2748
rect 18292 2746 18316 2748
rect 18372 2746 18396 2748
rect 18452 2746 18476 2748
rect 18532 2746 18556 2748
rect 18612 2746 18636 2748
rect 18692 2746 18706 2748
rect 17746 2694 17756 2746
rect 17812 2694 17822 2746
rect 18066 2694 18076 2746
rect 18132 2694 18142 2746
rect 18386 2694 18396 2746
rect 18452 2694 18462 2746
rect 17502 2692 17516 2694
rect 17572 2692 17596 2694
rect 17652 2692 17676 2694
rect 17732 2692 17756 2694
rect 17812 2692 17836 2694
rect 17892 2692 17916 2694
rect 17972 2692 17996 2694
rect 18052 2692 18076 2694
rect 18132 2692 18156 2694
rect 18212 2692 18236 2694
rect 18292 2692 18316 2694
rect 18372 2692 18396 2694
rect 18452 2692 18476 2694
rect 18532 2692 18556 2694
rect 18612 2692 18636 2694
rect 18692 2692 18706 2694
rect 17502 2683 18706 2692
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17052 2106 17080 2246
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 12256 2100 12308 2106
rect 12256 2042 12308 2048
rect 14832 2100 14884 2106
rect 14832 2042 14884 2048
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 15844 2032 15896 2038
rect 15844 1974 15896 1980
rect 15856 1601 15884 1974
rect 17880 1902 17908 2382
rect 17868 1896 17920 1902
rect 17868 1838 17920 1844
rect 18800 1698 18828 4490
rect 18892 4146 18920 10542
rect 18984 8974 19012 11766
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18984 5692 19012 8366
rect 19076 7585 19104 15506
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19260 10962 19288 12922
rect 19168 10934 19288 10962
rect 19062 7576 19118 7585
rect 19062 7511 19118 7520
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 19076 5817 19104 7414
rect 19062 5808 19118 5817
rect 19062 5743 19118 5752
rect 18984 5664 19104 5692
rect 18970 5264 19026 5273
rect 18970 5199 19026 5208
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18788 1692 18840 1698
rect 18788 1634 18840 1640
rect 15842 1592 15898 1601
rect 15842 1527 15898 1536
rect 10968 1352 11020 1358
rect 10968 1294 11020 1300
rect 15382 1320 15438 1329
rect 15382 1255 15384 1264
rect 15436 1255 15438 1264
rect 15384 1226 15436 1232
rect 9588 1216 9640 1222
rect 9588 1158 9640 1164
rect 8852 1080 8904 1086
rect 8852 1022 8904 1028
rect 5264 1012 5316 1018
rect 5264 954 5316 960
rect 18892 785 18920 3946
rect 18878 776 18934 785
rect 18878 711 18934 720
rect 18984 513 19012 5199
rect 19076 1057 19104 5664
rect 19168 5545 19196 10934
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19154 5536 19210 5545
rect 19154 5471 19210 5480
rect 19154 4040 19210 4049
rect 19154 3975 19210 3984
rect 19062 1048 19118 1057
rect 19062 983 19118 992
rect 18970 504 19026 513
rect 18970 439 19026 448
rect 4122 190 4200 218
rect 19062 232 19118 241
rect 4066 167 4122 176
rect 19168 218 19196 3975
rect 19260 2650 19288 10746
rect 19352 9654 19380 13942
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19430 13424 19486 13433
rect 19430 13359 19486 13368
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19352 7682 19380 9590
rect 19340 7676 19392 7682
rect 19340 7618 19392 7624
rect 19338 7576 19394 7585
rect 19338 7511 19394 7520
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19352 1766 19380 7511
rect 19444 4486 19472 13359
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19536 3466 19564 12650
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19628 3194 19656 13806
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19720 5370 19748 12582
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19706 5128 19762 5137
rect 19706 5063 19762 5072
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 19720 2961 19748 5063
rect 19706 2952 19762 2961
rect 19706 2887 19762 2896
rect 19720 2446 19748 2887
rect 19812 2553 19840 14282
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 19904 3058 19932 13874
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 19798 2544 19854 2553
rect 19798 2479 19854 2488
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 19340 1760 19392 1766
rect 19340 1702 19392 1708
rect 19118 190 19196 218
rect 19062 167 19118 176
<< via2 >>
rect 110 12688 166 12744
rect 18 10104 74 10160
rect 570 14320 626 14376
rect 754 14456 810 14512
rect 662 13096 718 13152
rect 754 11056 810 11112
rect 662 4528 718 4584
rect 5516 17434 5572 17436
rect 5596 17434 5652 17436
rect 5676 17434 5732 17436
rect 5756 17434 5812 17436
rect 5836 17434 5892 17436
rect 5916 17434 5972 17436
rect 5996 17434 6052 17436
rect 6076 17434 6132 17436
rect 6156 17434 6212 17436
rect 6236 17434 6292 17436
rect 6316 17434 6372 17436
rect 6396 17434 6452 17436
rect 6476 17434 6532 17436
rect 6556 17434 6612 17436
rect 6636 17434 6692 17436
rect 5516 17382 5554 17434
rect 5554 17382 5566 17434
rect 5566 17382 5572 17434
rect 5596 17382 5618 17434
rect 5618 17382 5630 17434
rect 5630 17382 5652 17434
rect 5676 17382 5682 17434
rect 5682 17382 5694 17434
rect 5694 17382 5732 17434
rect 5756 17382 5758 17434
rect 5758 17382 5810 17434
rect 5810 17382 5812 17434
rect 5836 17382 5874 17434
rect 5874 17382 5886 17434
rect 5886 17382 5892 17434
rect 5916 17382 5938 17434
rect 5938 17382 5950 17434
rect 5950 17382 5972 17434
rect 5996 17382 6002 17434
rect 6002 17382 6014 17434
rect 6014 17382 6052 17434
rect 6076 17382 6078 17434
rect 6078 17382 6130 17434
rect 6130 17382 6132 17434
rect 6156 17382 6194 17434
rect 6194 17382 6206 17434
rect 6206 17382 6212 17434
rect 6236 17382 6258 17434
rect 6258 17382 6270 17434
rect 6270 17382 6292 17434
rect 6316 17382 6322 17434
rect 6322 17382 6334 17434
rect 6334 17382 6372 17434
rect 6396 17382 6398 17434
rect 6398 17382 6450 17434
rect 6450 17382 6452 17434
rect 6476 17382 6514 17434
rect 6514 17382 6526 17434
rect 6526 17382 6532 17434
rect 6556 17382 6578 17434
rect 6578 17382 6590 17434
rect 6590 17382 6612 17434
rect 6636 17382 6642 17434
rect 6642 17382 6654 17434
rect 6654 17382 6692 17434
rect 5516 17380 5572 17382
rect 5596 17380 5652 17382
rect 5676 17380 5732 17382
rect 5756 17380 5812 17382
rect 5836 17380 5892 17382
rect 5916 17380 5972 17382
rect 5996 17380 6052 17382
rect 6076 17380 6132 17382
rect 6156 17380 6212 17382
rect 6236 17380 6292 17382
rect 6316 17380 6372 17382
rect 6396 17380 6452 17382
rect 6476 17380 6532 17382
rect 6556 17380 6612 17382
rect 6636 17380 6692 17382
rect 3330 17196 3386 17232
rect 3330 17176 3332 17196
rect 3332 17176 3384 17196
rect 3384 17176 3386 17196
rect 1516 16890 1572 16892
rect 1596 16890 1652 16892
rect 1676 16890 1732 16892
rect 1756 16890 1812 16892
rect 1836 16890 1892 16892
rect 1916 16890 1972 16892
rect 1996 16890 2052 16892
rect 2076 16890 2132 16892
rect 2156 16890 2212 16892
rect 2236 16890 2292 16892
rect 2316 16890 2372 16892
rect 2396 16890 2452 16892
rect 2476 16890 2532 16892
rect 2556 16890 2612 16892
rect 2636 16890 2692 16892
rect 1516 16838 1554 16890
rect 1554 16838 1566 16890
rect 1566 16838 1572 16890
rect 1596 16838 1618 16890
rect 1618 16838 1630 16890
rect 1630 16838 1652 16890
rect 1676 16838 1682 16890
rect 1682 16838 1694 16890
rect 1694 16838 1732 16890
rect 1756 16838 1758 16890
rect 1758 16838 1810 16890
rect 1810 16838 1812 16890
rect 1836 16838 1874 16890
rect 1874 16838 1886 16890
rect 1886 16838 1892 16890
rect 1916 16838 1938 16890
rect 1938 16838 1950 16890
rect 1950 16838 1972 16890
rect 1996 16838 2002 16890
rect 2002 16838 2014 16890
rect 2014 16838 2052 16890
rect 2076 16838 2078 16890
rect 2078 16838 2130 16890
rect 2130 16838 2132 16890
rect 2156 16838 2194 16890
rect 2194 16838 2206 16890
rect 2206 16838 2212 16890
rect 2236 16838 2258 16890
rect 2258 16838 2270 16890
rect 2270 16838 2292 16890
rect 2316 16838 2322 16890
rect 2322 16838 2334 16890
rect 2334 16838 2372 16890
rect 2396 16838 2398 16890
rect 2398 16838 2450 16890
rect 2450 16838 2452 16890
rect 2476 16838 2514 16890
rect 2514 16838 2526 16890
rect 2526 16838 2532 16890
rect 2556 16838 2578 16890
rect 2578 16838 2590 16890
rect 2590 16838 2612 16890
rect 2636 16838 2642 16890
rect 2642 16838 2654 16890
rect 2654 16838 2692 16890
rect 1516 16836 1572 16838
rect 1596 16836 1652 16838
rect 1676 16836 1732 16838
rect 1756 16836 1812 16838
rect 1836 16836 1892 16838
rect 1916 16836 1972 16838
rect 1996 16836 2052 16838
rect 2076 16836 2132 16838
rect 2156 16836 2212 16838
rect 2236 16836 2292 16838
rect 2316 16836 2372 16838
rect 2396 16836 2452 16838
rect 2476 16836 2532 16838
rect 2556 16836 2612 16838
rect 2636 16836 2692 16838
rect 1516 15802 1572 15804
rect 1596 15802 1652 15804
rect 1676 15802 1732 15804
rect 1756 15802 1812 15804
rect 1836 15802 1892 15804
rect 1916 15802 1972 15804
rect 1996 15802 2052 15804
rect 2076 15802 2132 15804
rect 2156 15802 2212 15804
rect 2236 15802 2292 15804
rect 2316 15802 2372 15804
rect 2396 15802 2452 15804
rect 2476 15802 2532 15804
rect 2556 15802 2612 15804
rect 2636 15802 2692 15804
rect 1516 15750 1554 15802
rect 1554 15750 1566 15802
rect 1566 15750 1572 15802
rect 1596 15750 1618 15802
rect 1618 15750 1630 15802
rect 1630 15750 1652 15802
rect 1676 15750 1682 15802
rect 1682 15750 1694 15802
rect 1694 15750 1732 15802
rect 1756 15750 1758 15802
rect 1758 15750 1810 15802
rect 1810 15750 1812 15802
rect 1836 15750 1874 15802
rect 1874 15750 1886 15802
rect 1886 15750 1892 15802
rect 1916 15750 1938 15802
rect 1938 15750 1950 15802
rect 1950 15750 1972 15802
rect 1996 15750 2002 15802
rect 2002 15750 2014 15802
rect 2014 15750 2052 15802
rect 2076 15750 2078 15802
rect 2078 15750 2130 15802
rect 2130 15750 2132 15802
rect 2156 15750 2194 15802
rect 2194 15750 2206 15802
rect 2206 15750 2212 15802
rect 2236 15750 2258 15802
rect 2258 15750 2270 15802
rect 2270 15750 2292 15802
rect 2316 15750 2322 15802
rect 2322 15750 2334 15802
rect 2334 15750 2372 15802
rect 2396 15750 2398 15802
rect 2398 15750 2450 15802
rect 2450 15750 2452 15802
rect 2476 15750 2514 15802
rect 2514 15750 2526 15802
rect 2526 15750 2532 15802
rect 2556 15750 2578 15802
rect 2578 15750 2590 15802
rect 2590 15750 2612 15802
rect 2636 15750 2642 15802
rect 2642 15750 2654 15802
rect 2654 15750 2692 15802
rect 1516 15748 1572 15750
rect 1596 15748 1652 15750
rect 1676 15748 1732 15750
rect 1756 15748 1812 15750
rect 1836 15748 1892 15750
rect 1916 15748 1972 15750
rect 1996 15748 2052 15750
rect 2076 15748 2132 15750
rect 2156 15748 2212 15750
rect 2236 15748 2292 15750
rect 2316 15748 2372 15750
rect 2396 15748 2452 15750
rect 2476 15748 2532 15750
rect 2556 15748 2612 15750
rect 2636 15748 2692 15750
rect 2778 14864 2834 14920
rect 1516 14714 1572 14716
rect 1596 14714 1652 14716
rect 1676 14714 1732 14716
rect 1756 14714 1812 14716
rect 1836 14714 1892 14716
rect 1916 14714 1972 14716
rect 1996 14714 2052 14716
rect 2076 14714 2132 14716
rect 2156 14714 2212 14716
rect 2236 14714 2292 14716
rect 2316 14714 2372 14716
rect 2396 14714 2452 14716
rect 2476 14714 2532 14716
rect 2556 14714 2612 14716
rect 2636 14714 2692 14716
rect 1516 14662 1554 14714
rect 1554 14662 1566 14714
rect 1566 14662 1572 14714
rect 1596 14662 1618 14714
rect 1618 14662 1630 14714
rect 1630 14662 1652 14714
rect 1676 14662 1682 14714
rect 1682 14662 1694 14714
rect 1694 14662 1732 14714
rect 1756 14662 1758 14714
rect 1758 14662 1810 14714
rect 1810 14662 1812 14714
rect 1836 14662 1874 14714
rect 1874 14662 1886 14714
rect 1886 14662 1892 14714
rect 1916 14662 1938 14714
rect 1938 14662 1950 14714
rect 1950 14662 1972 14714
rect 1996 14662 2002 14714
rect 2002 14662 2014 14714
rect 2014 14662 2052 14714
rect 2076 14662 2078 14714
rect 2078 14662 2130 14714
rect 2130 14662 2132 14714
rect 2156 14662 2194 14714
rect 2194 14662 2206 14714
rect 2206 14662 2212 14714
rect 2236 14662 2258 14714
rect 2258 14662 2270 14714
rect 2270 14662 2292 14714
rect 2316 14662 2322 14714
rect 2322 14662 2334 14714
rect 2334 14662 2372 14714
rect 2396 14662 2398 14714
rect 2398 14662 2450 14714
rect 2450 14662 2452 14714
rect 2476 14662 2514 14714
rect 2514 14662 2526 14714
rect 2526 14662 2532 14714
rect 2556 14662 2578 14714
rect 2578 14662 2590 14714
rect 2590 14662 2612 14714
rect 2636 14662 2642 14714
rect 2642 14662 2654 14714
rect 2654 14662 2692 14714
rect 1516 14660 1572 14662
rect 1596 14660 1652 14662
rect 1676 14660 1732 14662
rect 1756 14660 1812 14662
rect 1836 14660 1892 14662
rect 1916 14660 1972 14662
rect 1996 14660 2052 14662
rect 2076 14660 2132 14662
rect 2156 14660 2212 14662
rect 2236 14660 2292 14662
rect 2316 14660 2372 14662
rect 2396 14660 2452 14662
rect 2476 14660 2532 14662
rect 2556 14660 2612 14662
rect 2636 14660 2692 14662
rect 1582 14456 1638 14512
rect 1858 13776 1914 13832
rect 2226 13776 2282 13832
rect 1516 13626 1572 13628
rect 1596 13626 1652 13628
rect 1676 13626 1732 13628
rect 1756 13626 1812 13628
rect 1836 13626 1892 13628
rect 1916 13626 1972 13628
rect 1996 13626 2052 13628
rect 2076 13626 2132 13628
rect 2156 13626 2212 13628
rect 2236 13626 2292 13628
rect 2316 13626 2372 13628
rect 2396 13626 2452 13628
rect 2476 13626 2532 13628
rect 2556 13626 2612 13628
rect 2636 13626 2692 13628
rect 1516 13574 1554 13626
rect 1554 13574 1566 13626
rect 1566 13574 1572 13626
rect 1596 13574 1618 13626
rect 1618 13574 1630 13626
rect 1630 13574 1652 13626
rect 1676 13574 1682 13626
rect 1682 13574 1694 13626
rect 1694 13574 1732 13626
rect 1756 13574 1758 13626
rect 1758 13574 1810 13626
rect 1810 13574 1812 13626
rect 1836 13574 1874 13626
rect 1874 13574 1886 13626
rect 1886 13574 1892 13626
rect 1916 13574 1938 13626
rect 1938 13574 1950 13626
rect 1950 13574 1972 13626
rect 1996 13574 2002 13626
rect 2002 13574 2014 13626
rect 2014 13574 2052 13626
rect 2076 13574 2078 13626
rect 2078 13574 2130 13626
rect 2130 13574 2132 13626
rect 2156 13574 2194 13626
rect 2194 13574 2206 13626
rect 2206 13574 2212 13626
rect 2236 13574 2258 13626
rect 2258 13574 2270 13626
rect 2270 13574 2292 13626
rect 2316 13574 2322 13626
rect 2322 13574 2334 13626
rect 2334 13574 2372 13626
rect 2396 13574 2398 13626
rect 2398 13574 2450 13626
rect 2450 13574 2452 13626
rect 2476 13574 2514 13626
rect 2514 13574 2526 13626
rect 2526 13574 2532 13626
rect 2556 13574 2578 13626
rect 2578 13574 2590 13626
rect 2590 13574 2612 13626
rect 2636 13574 2642 13626
rect 2642 13574 2654 13626
rect 2654 13574 2692 13626
rect 1516 13572 1572 13574
rect 1596 13572 1652 13574
rect 1676 13572 1732 13574
rect 1756 13572 1812 13574
rect 1836 13572 1892 13574
rect 1916 13572 1972 13574
rect 1996 13572 2052 13574
rect 2076 13572 2132 13574
rect 2156 13572 2212 13574
rect 2236 13572 2292 13574
rect 2316 13572 2372 13574
rect 2396 13572 2452 13574
rect 2476 13572 2532 13574
rect 2556 13572 2612 13574
rect 2636 13572 2692 13574
rect 1766 13368 1822 13424
rect 1950 13252 2006 13288
rect 1950 13232 1952 13252
rect 1952 13232 2004 13252
rect 2004 13232 2006 13252
rect 2318 13368 2374 13424
rect 2318 12824 2374 12880
rect 2962 13640 3018 13696
rect 2870 12824 2926 12880
rect 2686 12688 2742 12744
rect 1516 12538 1572 12540
rect 1596 12538 1652 12540
rect 1676 12538 1732 12540
rect 1756 12538 1812 12540
rect 1836 12538 1892 12540
rect 1916 12538 1972 12540
rect 1996 12538 2052 12540
rect 2076 12538 2132 12540
rect 2156 12538 2212 12540
rect 2236 12538 2292 12540
rect 2316 12538 2372 12540
rect 2396 12538 2452 12540
rect 2476 12538 2532 12540
rect 2556 12538 2612 12540
rect 2636 12538 2692 12540
rect 1516 12486 1554 12538
rect 1554 12486 1566 12538
rect 1566 12486 1572 12538
rect 1596 12486 1618 12538
rect 1618 12486 1630 12538
rect 1630 12486 1652 12538
rect 1676 12486 1682 12538
rect 1682 12486 1694 12538
rect 1694 12486 1732 12538
rect 1756 12486 1758 12538
rect 1758 12486 1810 12538
rect 1810 12486 1812 12538
rect 1836 12486 1874 12538
rect 1874 12486 1886 12538
rect 1886 12486 1892 12538
rect 1916 12486 1938 12538
rect 1938 12486 1950 12538
rect 1950 12486 1972 12538
rect 1996 12486 2002 12538
rect 2002 12486 2014 12538
rect 2014 12486 2052 12538
rect 2076 12486 2078 12538
rect 2078 12486 2130 12538
rect 2130 12486 2132 12538
rect 2156 12486 2194 12538
rect 2194 12486 2206 12538
rect 2206 12486 2212 12538
rect 2236 12486 2258 12538
rect 2258 12486 2270 12538
rect 2270 12486 2292 12538
rect 2316 12486 2322 12538
rect 2322 12486 2334 12538
rect 2334 12486 2372 12538
rect 2396 12486 2398 12538
rect 2398 12486 2450 12538
rect 2450 12486 2452 12538
rect 2476 12486 2514 12538
rect 2514 12486 2526 12538
rect 2526 12486 2532 12538
rect 2556 12486 2578 12538
rect 2578 12486 2590 12538
rect 2590 12486 2612 12538
rect 2636 12486 2642 12538
rect 2642 12486 2654 12538
rect 2654 12486 2692 12538
rect 1516 12484 1572 12486
rect 1596 12484 1652 12486
rect 1676 12484 1732 12486
rect 1756 12484 1812 12486
rect 1836 12484 1892 12486
rect 1916 12484 1972 12486
rect 1996 12484 2052 12486
rect 2076 12484 2132 12486
rect 2156 12484 2212 12486
rect 2236 12484 2292 12486
rect 2316 12484 2372 12486
rect 2396 12484 2452 12486
rect 2476 12484 2532 12486
rect 2556 12484 2612 12486
rect 2636 12484 2692 12486
rect 2318 12300 2374 12336
rect 2318 12280 2320 12300
rect 2320 12280 2372 12300
rect 2372 12280 2374 12300
rect 2226 12144 2282 12200
rect 2410 11600 2466 11656
rect 2870 12280 2926 12336
rect 2594 11772 2596 11792
rect 2596 11772 2648 11792
rect 2648 11772 2650 11792
rect 2594 11736 2650 11772
rect 1516 11450 1572 11452
rect 1596 11450 1652 11452
rect 1676 11450 1732 11452
rect 1756 11450 1812 11452
rect 1836 11450 1892 11452
rect 1916 11450 1972 11452
rect 1996 11450 2052 11452
rect 2076 11450 2132 11452
rect 2156 11450 2212 11452
rect 2236 11450 2292 11452
rect 2316 11450 2372 11452
rect 2396 11450 2452 11452
rect 2476 11450 2532 11452
rect 2556 11450 2612 11452
rect 2636 11450 2692 11452
rect 1516 11398 1554 11450
rect 1554 11398 1566 11450
rect 1566 11398 1572 11450
rect 1596 11398 1618 11450
rect 1618 11398 1630 11450
rect 1630 11398 1652 11450
rect 1676 11398 1682 11450
rect 1682 11398 1694 11450
rect 1694 11398 1732 11450
rect 1756 11398 1758 11450
rect 1758 11398 1810 11450
rect 1810 11398 1812 11450
rect 1836 11398 1874 11450
rect 1874 11398 1886 11450
rect 1886 11398 1892 11450
rect 1916 11398 1938 11450
rect 1938 11398 1950 11450
rect 1950 11398 1972 11450
rect 1996 11398 2002 11450
rect 2002 11398 2014 11450
rect 2014 11398 2052 11450
rect 2076 11398 2078 11450
rect 2078 11398 2130 11450
rect 2130 11398 2132 11450
rect 2156 11398 2194 11450
rect 2194 11398 2206 11450
rect 2206 11398 2212 11450
rect 2236 11398 2258 11450
rect 2258 11398 2270 11450
rect 2270 11398 2292 11450
rect 2316 11398 2322 11450
rect 2322 11398 2334 11450
rect 2334 11398 2372 11450
rect 2396 11398 2398 11450
rect 2398 11398 2450 11450
rect 2450 11398 2452 11450
rect 2476 11398 2514 11450
rect 2514 11398 2526 11450
rect 2526 11398 2532 11450
rect 2556 11398 2578 11450
rect 2578 11398 2590 11450
rect 2590 11398 2612 11450
rect 2636 11398 2642 11450
rect 2642 11398 2654 11450
rect 2654 11398 2692 11450
rect 1516 11396 1572 11398
rect 1596 11396 1652 11398
rect 1676 11396 1732 11398
rect 1756 11396 1812 11398
rect 1836 11396 1892 11398
rect 1916 11396 1972 11398
rect 1996 11396 2052 11398
rect 2076 11396 2132 11398
rect 2156 11396 2212 11398
rect 2236 11396 2292 11398
rect 2316 11396 2372 11398
rect 2396 11396 2452 11398
rect 2476 11396 2532 11398
rect 2556 11396 2612 11398
rect 2636 11396 2692 11398
rect 1858 10920 1914 10976
rect 938 3712 994 3768
rect 1516 10362 1572 10364
rect 1596 10362 1652 10364
rect 1676 10362 1732 10364
rect 1756 10362 1812 10364
rect 1836 10362 1892 10364
rect 1916 10362 1972 10364
rect 1996 10362 2052 10364
rect 2076 10362 2132 10364
rect 2156 10362 2212 10364
rect 2236 10362 2292 10364
rect 2316 10362 2372 10364
rect 2396 10362 2452 10364
rect 2476 10362 2532 10364
rect 2556 10362 2612 10364
rect 2636 10362 2692 10364
rect 1516 10310 1554 10362
rect 1554 10310 1566 10362
rect 1566 10310 1572 10362
rect 1596 10310 1618 10362
rect 1618 10310 1630 10362
rect 1630 10310 1652 10362
rect 1676 10310 1682 10362
rect 1682 10310 1694 10362
rect 1694 10310 1732 10362
rect 1756 10310 1758 10362
rect 1758 10310 1810 10362
rect 1810 10310 1812 10362
rect 1836 10310 1874 10362
rect 1874 10310 1886 10362
rect 1886 10310 1892 10362
rect 1916 10310 1938 10362
rect 1938 10310 1950 10362
rect 1950 10310 1972 10362
rect 1996 10310 2002 10362
rect 2002 10310 2014 10362
rect 2014 10310 2052 10362
rect 2076 10310 2078 10362
rect 2078 10310 2130 10362
rect 2130 10310 2132 10362
rect 2156 10310 2194 10362
rect 2194 10310 2206 10362
rect 2206 10310 2212 10362
rect 2236 10310 2258 10362
rect 2258 10310 2270 10362
rect 2270 10310 2292 10362
rect 2316 10310 2322 10362
rect 2322 10310 2334 10362
rect 2334 10310 2372 10362
rect 2396 10310 2398 10362
rect 2398 10310 2450 10362
rect 2450 10310 2452 10362
rect 2476 10310 2514 10362
rect 2514 10310 2526 10362
rect 2526 10310 2532 10362
rect 2556 10310 2578 10362
rect 2578 10310 2590 10362
rect 2590 10310 2612 10362
rect 2636 10310 2642 10362
rect 2642 10310 2654 10362
rect 2654 10310 2692 10362
rect 1516 10308 1572 10310
rect 1596 10308 1652 10310
rect 1676 10308 1732 10310
rect 1756 10308 1812 10310
rect 1836 10308 1892 10310
rect 1916 10308 1972 10310
rect 1996 10308 2052 10310
rect 2076 10308 2132 10310
rect 2156 10308 2212 10310
rect 2236 10308 2292 10310
rect 2316 10308 2372 10310
rect 2396 10308 2452 10310
rect 2476 10308 2532 10310
rect 2556 10308 2612 10310
rect 2636 10308 2692 10310
rect 1516 9274 1572 9276
rect 1596 9274 1652 9276
rect 1676 9274 1732 9276
rect 1756 9274 1812 9276
rect 1836 9274 1892 9276
rect 1916 9274 1972 9276
rect 1996 9274 2052 9276
rect 2076 9274 2132 9276
rect 2156 9274 2212 9276
rect 2236 9274 2292 9276
rect 2316 9274 2372 9276
rect 2396 9274 2452 9276
rect 2476 9274 2532 9276
rect 2556 9274 2612 9276
rect 2636 9274 2692 9276
rect 1516 9222 1554 9274
rect 1554 9222 1566 9274
rect 1566 9222 1572 9274
rect 1596 9222 1618 9274
rect 1618 9222 1630 9274
rect 1630 9222 1652 9274
rect 1676 9222 1682 9274
rect 1682 9222 1694 9274
rect 1694 9222 1732 9274
rect 1756 9222 1758 9274
rect 1758 9222 1810 9274
rect 1810 9222 1812 9274
rect 1836 9222 1874 9274
rect 1874 9222 1886 9274
rect 1886 9222 1892 9274
rect 1916 9222 1938 9274
rect 1938 9222 1950 9274
rect 1950 9222 1972 9274
rect 1996 9222 2002 9274
rect 2002 9222 2014 9274
rect 2014 9222 2052 9274
rect 2076 9222 2078 9274
rect 2078 9222 2130 9274
rect 2130 9222 2132 9274
rect 2156 9222 2194 9274
rect 2194 9222 2206 9274
rect 2206 9222 2212 9274
rect 2236 9222 2258 9274
rect 2258 9222 2270 9274
rect 2270 9222 2292 9274
rect 2316 9222 2322 9274
rect 2322 9222 2334 9274
rect 2334 9222 2372 9274
rect 2396 9222 2398 9274
rect 2398 9222 2450 9274
rect 2450 9222 2452 9274
rect 2476 9222 2514 9274
rect 2514 9222 2526 9274
rect 2526 9222 2532 9274
rect 2556 9222 2578 9274
rect 2578 9222 2590 9274
rect 2590 9222 2612 9274
rect 2636 9222 2642 9274
rect 2642 9222 2654 9274
rect 2654 9222 2692 9274
rect 1516 9220 1572 9222
rect 1596 9220 1652 9222
rect 1676 9220 1732 9222
rect 1756 9220 1812 9222
rect 1836 9220 1892 9222
rect 1916 9220 1972 9222
rect 1996 9220 2052 9222
rect 2076 9220 2132 9222
rect 2156 9220 2212 9222
rect 2236 9220 2292 9222
rect 2316 9220 2372 9222
rect 2396 9220 2452 9222
rect 2476 9220 2532 9222
rect 2556 9220 2612 9222
rect 2636 9220 2692 9222
rect 3146 12416 3202 12472
rect 3146 12008 3202 12064
rect 3146 11600 3202 11656
rect 1516 8186 1572 8188
rect 1596 8186 1652 8188
rect 1676 8186 1732 8188
rect 1756 8186 1812 8188
rect 1836 8186 1892 8188
rect 1916 8186 1972 8188
rect 1996 8186 2052 8188
rect 2076 8186 2132 8188
rect 2156 8186 2212 8188
rect 2236 8186 2292 8188
rect 2316 8186 2372 8188
rect 2396 8186 2452 8188
rect 2476 8186 2532 8188
rect 2556 8186 2612 8188
rect 2636 8186 2692 8188
rect 1516 8134 1554 8186
rect 1554 8134 1566 8186
rect 1566 8134 1572 8186
rect 1596 8134 1618 8186
rect 1618 8134 1630 8186
rect 1630 8134 1652 8186
rect 1676 8134 1682 8186
rect 1682 8134 1694 8186
rect 1694 8134 1732 8186
rect 1756 8134 1758 8186
rect 1758 8134 1810 8186
rect 1810 8134 1812 8186
rect 1836 8134 1874 8186
rect 1874 8134 1886 8186
rect 1886 8134 1892 8186
rect 1916 8134 1938 8186
rect 1938 8134 1950 8186
rect 1950 8134 1972 8186
rect 1996 8134 2002 8186
rect 2002 8134 2014 8186
rect 2014 8134 2052 8186
rect 2076 8134 2078 8186
rect 2078 8134 2130 8186
rect 2130 8134 2132 8186
rect 2156 8134 2194 8186
rect 2194 8134 2206 8186
rect 2206 8134 2212 8186
rect 2236 8134 2258 8186
rect 2258 8134 2270 8186
rect 2270 8134 2292 8186
rect 2316 8134 2322 8186
rect 2322 8134 2334 8186
rect 2334 8134 2372 8186
rect 2396 8134 2398 8186
rect 2398 8134 2450 8186
rect 2450 8134 2452 8186
rect 2476 8134 2514 8186
rect 2514 8134 2526 8186
rect 2526 8134 2532 8186
rect 2556 8134 2578 8186
rect 2578 8134 2590 8186
rect 2590 8134 2612 8186
rect 2636 8134 2642 8186
rect 2642 8134 2654 8186
rect 2654 8134 2692 8186
rect 1516 8132 1572 8134
rect 1596 8132 1652 8134
rect 1676 8132 1732 8134
rect 1756 8132 1812 8134
rect 1836 8132 1892 8134
rect 1916 8132 1972 8134
rect 1996 8132 2052 8134
rect 2076 8132 2132 8134
rect 2156 8132 2212 8134
rect 2236 8132 2292 8134
rect 2316 8132 2372 8134
rect 2396 8132 2452 8134
rect 2476 8132 2532 8134
rect 2556 8132 2612 8134
rect 2636 8132 2692 8134
rect 1516 7098 1572 7100
rect 1596 7098 1652 7100
rect 1676 7098 1732 7100
rect 1756 7098 1812 7100
rect 1836 7098 1892 7100
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 2316 7098 2372 7100
rect 2396 7098 2452 7100
rect 2476 7098 2532 7100
rect 2556 7098 2612 7100
rect 2636 7098 2692 7100
rect 1516 7046 1554 7098
rect 1554 7046 1566 7098
rect 1566 7046 1572 7098
rect 1596 7046 1618 7098
rect 1618 7046 1630 7098
rect 1630 7046 1652 7098
rect 1676 7046 1682 7098
rect 1682 7046 1694 7098
rect 1694 7046 1732 7098
rect 1756 7046 1758 7098
rect 1758 7046 1810 7098
rect 1810 7046 1812 7098
rect 1836 7046 1874 7098
rect 1874 7046 1886 7098
rect 1886 7046 1892 7098
rect 1916 7046 1938 7098
rect 1938 7046 1950 7098
rect 1950 7046 1972 7098
rect 1996 7046 2002 7098
rect 2002 7046 2014 7098
rect 2014 7046 2052 7098
rect 2076 7046 2078 7098
rect 2078 7046 2130 7098
rect 2130 7046 2132 7098
rect 2156 7046 2194 7098
rect 2194 7046 2206 7098
rect 2206 7046 2212 7098
rect 2236 7046 2258 7098
rect 2258 7046 2270 7098
rect 2270 7046 2292 7098
rect 2316 7046 2322 7098
rect 2322 7046 2334 7098
rect 2334 7046 2372 7098
rect 2396 7046 2398 7098
rect 2398 7046 2450 7098
rect 2450 7046 2452 7098
rect 2476 7046 2514 7098
rect 2514 7046 2526 7098
rect 2526 7046 2532 7098
rect 2556 7046 2578 7098
rect 2578 7046 2590 7098
rect 2590 7046 2612 7098
rect 2636 7046 2642 7098
rect 2642 7046 2654 7098
rect 2654 7046 2692 7098
rect 1516 7044 1572 7046
rect 1596 7044 1652 7046
rect 1676 7044 1732 7046
rect 1756 7044 1812 7046
rect 1836 7044 1892 7046
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 2316 7044 2372 7046
rect 2396 7044 2452 7046
rect 2476 7044 2532 7046
rect 2556 7044 2612 7046
rect 2636 7044 2692 7046
rect 3514 13096 3570 13152
rect 3422 11872 3478 11928
rect 3422 9968 3478 10024
rect 1516 6010 1572 6012
rect 1596 6010 1652 6012
rect 1676 6010 1732 6012
rect 1756 6010 1812 6012
rect 1836 6010 1892 6012
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 2316 6010 2372 6012
rect 2396 6010 2452 6012
rect 2476 6010 2532 6012
rect 2556 6010 2612 6012
rect 2636 6010 2692 6012
rect 1516 5958 1554 6010
rect 1554 5958 1566 6010
rect 1566 5958 1572 6010
rect 1596 5958 1618 6010
rect 1618 5958 1630 6010
rect 1630 5958 1652 6010
rect 1676 5958 1682 6010
rect 1682 5958 1694 6010
rect 1694 5958 1732 6010
rect 1756 5958 1758 6010
rect 1758 5958 1810 6010
rect 1810 5958 1812 6010
rect 1836 5958 1874 6010
rect 1874 5958 1886 6010
rect 1886 5958 1892 6010
rect 1916 5958 1938 6010
rect 1938 5958 1950 6010
rect 1950 5958 1972 6010
rect 1996 5958 2002 6010
rect 2002 5958 2014 6010
rect 2014 5958 2052 6010
rect 2076 5958 2078 6010
rect 2078 5958 2130 6010
rect 2130 5958 2132 6010
rect 2156 5958 2194 6010
rect 2194 5958 2206 6010
rect 2206 5958 2212 6010
rect 2236 5958 2258 6010
rect 2258 5958 2270 6010
rect 2270 5958 2292 6010
rect 2316 5958 2322 6010
rect 2322 5958 2334 6010
rect 2334 5958 2372 6010
rect 2396 5958 2398 6010
rect 2398 5958 2450 6010
rect 2450 5958 2452 6010
rect 2476 5958 2514 6010
rect 2514 5958 2526 6010
rect 2526 5958 2532 6010
rect 2556 5958 2578 6010
rect 2578 5958 2590 6010
rect 2590 5958 2612 6010
rect 2636 5958 2642 6010
rect 2642 5958 2654 6010
rect 2654 5958 2692 6010
rect 1516 5956 1572 5958
rect 1596 5956 1652 5958
rect 1676 5956 1732 5958
rect 1756 5956 1812 5958
rect 1836 5956 1892 5958
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 2316 5956 2372 5958
rect 2396 5956 2452 5958
rect 2476 5956 2532 5958
rect 2556 5956 2612 5958
rect 2636 5956 2692 5958
rect 1516 4922 1572 4924
rect 1596 4922 1652 4924
rect 1676 4922 1732 4924
rect 1756 4922 1812 4924
rect 1836 4922 1892 4924
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 2316 4922 2372 4924
rect 2396 4922 2452 4924
rect 2476 4922 2532 4924
rect 2556 4922 2612 4924
rect 2636 4922 2692 4924
rect 1516 4870 1554 4922
rect 1554 4870 1566 4922
rect 1566 4870 1572 4922
rect 1596 4870 1618 4922
rect 1618 4870 1630 4922
rect 1630 4870 1652 4922
rect 1676 4870 1682 4922
rect 1682 4870 1694 4922
rect 1694 4870 1732 4922
rect 1756 4870 1758 4922
rect 1758 4870 1810 4922
rect 1810 4870 1812 4922
rect 1836 4870 1874 4922
rect 1874 4870 1886 4922
rect 1886 4870 1892 4922
rect 1916 4870 1938 4922
rect 1938 4870 1950 4922
rect 1950 4870 1972 4922
rect 1996 4870 2002 4922
rect 2002 4870 2014 4922
rect 2014 4870 2052 4922
rect 2076 4870 2078 4922
rect 2078 4870 2130 4922
rect 2130 4870 2132 4922
rect 2156 4870 2194 4922
rect 2194 4870 2206 4922
rect 2206 4870 2212 4922
rect 2236 4870 2258 4922
rect 2258 4870 2270 4922
rect 2270 4870 2292 4922
rect 2316 4870 2322 4922
rect 2322 4870 2334 4922
rect 2334 4870 2372 4922
rect 2396 4870 2398 4922
rect 2398 4870 2450 4922
rect 2450 4870 2452 4922
rect 2476 4870 2514 4922
rect 2514 4870 2526 4922
rect 2526 4870 2532 4922
rect 2556 4870 2578 4922
rect 2578 4870 2590 4922
rect 2590 4870 2612 4922
rect 2636 4870 2642 4922
rect 2642 4870 2654 4922
rect 2654 4870 2692 4922
rect 1516 4868 1572 4870
rect 1596 4868 1652 4870
rect 1676 4868 1732 4870
rect 1756 4868 1812 4870
rect 1836 4868 1892 4870
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 2316 4868 2372 4870
rect 2396 4868 2452 4870
rect 2476 4868 2532 4870
rect 2556 4868 2612 4870
rect 2636 4868 2692 4870
rect 1398 3984 1454 4040
rect 1516 3834 1572 3836
rect 1596 3834 1652 3836
rect 1676 3834 1732 3836
rect 1756 3834 1812 3836
rect 1836 3834 1892 3836
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 2316 3834 2372 3836
rect 2396 3834 2452 3836
rect 2476 3834 2532 3836
rect 2556 3834 2612 3836
rect 2636 3834 2692 3836
rect 1516 3782 1554 3834
rect 1554 3782 1566 3834
rect 1566 3782 1572 3834
rect 1596 3782 1618 3834
rect 1618 3782 1630 3834
rect 1630 3782 1652 3834
rect 1676 3782 1682 3834
rect 1682 3782 1694 3834
rect 1694 3782 1732 3834
rect 1756 3782 1758 3834
rect 1758 3782 1810 3834
rect 1810 3782 1812 3834
rect 1836 3782 1874 3834
rect 1874 3782 1886 3834
rect 1886 3782 1892 3834
rect 1916 3782 1938 3834
rect 1938 3782 1950 3834
rect 1950 3782 1972 3834
rect 1996 3782 2002 3834
rect 2002 3782 2014 3834
rect 2014 3782 2052 3834
rect 2076 3782 2078 3834
rect 2078 3782 2130 3834
rect 2130 3782 2132 3834
rect 2156 3782 2194 3834
rect 2194 3782 2206 3834
rect 2206 3782 2212 3834
rect 2236 3782 2258 3834
rect 2258 3782 2270 3834
rect 2270 3782 2292 3834
rect 2316 3782 2322 3834
rect 2322 3782 2334 3834
rect 2334 3782 2372 3834
rect 2396 3782 2398 3834
rect 2398 3782 2450 3834
rect 2450 3782 2452 3834
rect 2476 3782 2514 3834
rect 2514 3782 2526 3834
rect 2526 3782 2532 3834
rect 2556 3782 2578 3834
rect 2578 3782 2590 3834
rect 2590 3782 2612 3834
rect 2636 3782 2642 3834
rect 2642 3782 2654 3834
rect 2654 3782 2692 3834
rect 1516 3780 1572 3782
rect 1596 3780 1652 3782
rect 1676 3780 1732 3782
rect 1756 3780 1812 3782
rect 1836 3780 1892 3782
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 2316 3780 2372 3782
rect 2396 3780 2452 3782
rect 2476 3780 2532 3782
rect 2556 3780 2612 3782
rect 2636 3780 2692 3782
rect 1122 3440 1178 3496
rect 1030 3168 1086 3224
rect 938 2896 994 2952
rect 938 2352 994 2408
rect 1030 2080 1086 2136
rect 3882 12416 3938 12472
rect 4158 13368 4214 13424
rect 4526 14456 4582 14512
rect 4526 14184 4582 14240
rect 4526 14068 4582 14104
rect 4526 14048 4528 14068
rect 4528 14048 4580 14068
rect 4580 14048 4582 14068
rect 4434 13504 4490 13560
rect 4250 13232 4306 13288
rect 4066 12960 4122 13016
rect 4434 12280 4490 12336
rect 3790 11756 3846 11792
rect 3790 11736 3792 11756
rect 3792 11736 3844 11756
rect 3844 11736 3846 11756
rect 3974 11056 4030 11112
rect 4158 10784 4214 10840
rect 4066 10512 4122 10568
rect 1516 2746 1572 2748
rect 1596 2746 1652 2748
rect 1676 2746 1732 2748
rect 1756 2746 1812 2748
rect 1836 2746 1892 2748
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 2316 2746 2372 2748
rect 2396 2746 2452 2748
rect 2476 2746 2532 2748
rect 2556 2746 2612 2748
rect 2636 2746 2692 2748
rect 1516 2694 1554 2746
rect 1554 2694 1566 2746
rect 1566 2694 1572 2746
rect 1596 2694 1618 2746
rect 1618 2694 1630 2746
rect 1630 2694 1652 2746
rect 1676 2694 1682 2746
rect 1682 2694 1694 2746
rect 1694 2694 1732 2746
rect 1756 2694 1758 2746
rect 1758 2694 1810 2746
rect 1810 2694 1812 2746
rect 1836 2694 1874 2746
rect 1874 2694 1886 2746
rect 1886 2694 1892 2746
rect 1916 2694 1938 2746
rect 1938 2694 1950 2746
rect 1950 2694 1972 2746
rect 1996 2694 2002 2746
rect 2002 2694 2014 2746
rect 2014 2694 2052 2746
rect 2076 2694 2078 2746
rect 2078 2694 2130 2746
rect 2130 2694 2132 2746
rect 2156 2694 2194 2746
rect 2194 2694 2206 2746
rect 2206 2694 2212 2746
rect 2236 2694 2258 2746
rect 2258 2694 2270 2746
rect 2270 2694 2292 2746
rect 2316 2694 2322 2746
rect 2322 2694 2334 2746
rect 2334 2694 2372 2746
rect 2396 2694 2398 2746
rect 2398 2694 2450 2746
rect 2450 2694 2452 2746
rect 2476 2694 2514 2746
rect 2514 2694 2526 2746
rect 2526 2694 2532 2746
rect 2556 2694 2578 2746
rect 2578 2694 2590 2746
rect 2590 2694 2612 2746
rect 2636 2694 2642 2746
rect 2642 2694 2654 2746
rect 2654 2694 2692 2746
rect 1516 2692 1572 2694
rect 1596 2692 1652 2694
rect 1676 2692 1732 2694
rect 1756 2692 1812 2694
rect 1836 2692 1892 2694
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 2316 2692 2372 2694
rect 2396 2692 2452 2694
rect 2476 2692 2532 2694
rect 2556 2692 2612 2694
rect 2636 2692 2692 2694
rect 3698 2488 3754 2544
rect 3422 1828 3478 1864
rect 3422 1808 3424 1828
rect 3424 1808 3476 1828
rect 3476 1808 3478 1828
rect 3514 1536 3570 1592
rect 1122 1264 1178 1320
rect 3330 720 3386 776
rect 4158 9016 4214 9072
rect 4342 10784 4398 10840
rect 5446 16632 5502 16688
rect 5170 15428 5226 15464
rect 5170 15408 5172 15428
rect 5172 15408 5224 15428
rect 5224 15408 5226 15428
rect 4986 15000 5042 15056
rect 4894 14864 4950 14920
rect 5078 13776 5134 13832
rect 5516 16346 5572 16348
rect 5596 16346 5652 16348
rect 5676 16346 5732 16348
rect 5756 16346 5812 16348
rect 5836 16346 5892 16348
rect 5916 16346 5972 16348
rect 5996 16346 6052 16348
rect 6076 16346 6132 16348
rect 6156 16346 6212 16348
rect 6236 16346 6292 16348
rect 6316 16346 6372 16348
rect 6396 16346 6452 16348
rect 6476 16346 6532 16348
rect 6556 16346 6612 16348
rect 6636 16346 6692 16348
rect 5516 16294 5554 16346
rect 5554 16294 5566 16346
rect 5566 16294 5572 16346
rect 5596 16294 5618 16346
rect 5618 16294 5630 16346
rect 5630 16294 5652 16346
rect 5676 16294 5682 16346
rect 5682 16294 5694 16346
rect 5694 16294 5732 16346
rect 5756 16294 5758 16346
rect 5758 16294 5810 16346
rect 5810 16294 5812 16346
rect 5836 16294 5874 16346
rect 5874 16294 5886 16346
rect 5886 16294 5892 16346
rect 5916 16294 5938 16346
rect 5938 16294 5950 16346
rect 5950 16294 5972 16346
rect 5996 16294 6002 16346
rect 6002 16294 6014 16346
rect 6014 16294 6052 16346
rect 6076 16294 6078 16346
rect 6078 16294 6130 16346
rect 6130 16294 6132 16346
rect 6156 16294 6194 16346
rect 6194 16294 6206 16346
rect 6206 16294 6212 16346
rect 6236 16294 6258 16346
rect 6258 16294 6270 16346
rect 6270 16294 6292 16346
rect 6316 16294 6322 16346
rect 6322 16294 6334 16346
rect 6334 16294 6372 16346
rect 6396 16294 6398 16346
rect 6398 16294 6450 16346
rect 6450 16294 6452 16346
rect 6476 16294 6514 16346
rect 6514 16294 6526 16346
rect 6526 16294 6532 16346
rect 6556 16294 6578 16346
rect 6578 16294 6590 16346
rect 6590 16294 6612 16346
rect 6636 16294 6642 16346
rect 6642 16294 6654 16346
rect 6654 16294 6692 16346
rect 5516 16292 5572 16294
rect 5596 16292 5652 16294
rect 5676 16292 5732 16294
rect 5756 16292 5812 16294
rect 5836 16292 5892 16294
rect 5916 16292 5972 16294
rect 5996 16292 6052 16294
rect 6076 16292 6132 16294
rect 6156 16292 6212 16294
rect 6236 16292 6292 16294
rect 6316 16292 6372 16294
rect 6396 16292 6452 16294
rect 6476 16292 6532 16294
rect 6556 16292 6612 16294
rect 6636 16292 6692 16294
rect 6182 15700 6238 15736
rect 6182 15680 6184 15700
rect 6184 15680 6236 15700
rect 6236 15680 6238 15700
rect 5446 15544 5502 15600
rect 5516 15258 5572 15260
rect 5596 15258 5652 15260
rect 5676 15258 5732 15260
rect 5756 15258 5812 15260
rect 5836 15258 5892 15260
rect 5916 15258 5972 15260
rect 5996 15258 6052 15260
rect 6076 15258 6132 15260
rect 6156 15258 6212 15260
rect 6236 15258 6292 15260
rect 6316 15258 6372 15260
rect 6396 15258 6452 15260
rect 6476 15258 6532 15260
rect 6556 15258 6612 15260
rect 6636 15258 6692 15260
rect 5516 15206 5554 15258
rect 5554 15206 5566 15258
rect 5566 15206 5572 15258
rect 5596 15206 5618 15258
rect 5618 15206 5630 15258
rect 5630 15206 5652 15258
rect 5676 15206 5682 15258
rect 5682 15206 5694 15258
rect 5694 15206 5732 15258
rect 5756 15206 5758 15258
rect 5758 15206 5810 15258
rect 5810 15206 5812 15258
rect 5836 15206 5874 15258
rect 5874 15206 5886 15258
rect 5886 15206 5892 15258
rect 5916 15206 5938 15258
rect 5938 15206 5950 15258
rect 5950 15206 5972 15258
rect 5996 15206 6002 15258
rect 6002 15206 6014 15258
rect 6014 15206 6052 15258
rect 6076 15206 6078 15258
rect 6078 15206 6130 15258
rect 6130 15206 6132 15258
rect 6156 15206 6194 15258
rect 6194 15206 6206 15258
rect 6206 15206 6212 15258
rect 6236 15206 6258 15258
rect 6258 15206 6270 15258
rect 6270 15206 6292 15258
rect 6316 15206 6322 15258
rect 6322 15206 6334 15258
rect 6334 15206 6372 15258
rect 6396 15206 6398 15258
rect 6398 15206 6450 15258
rect 6450 15206 6452 15258
rect 6476 15206 6514 15258
rect 6514 15206 6526 15258
rect 6526 15206 6532 15258
rect 6556 15206 6578 15258
rect 6578 15206 6590 15258
rect 6590 15206 6612 15258
rect 6636 15206 6642 15258
rect 6642 15206 6654 15258
rect 6654 15206 6692 15258
rect 5516 15204 5572 15206
rect 5596 15204 5652 15206
rect 5676 15204 5732 15206
rect 5756 15204 5812 15206
rect 5836 15204 5892 15206
rect 5916 15204 5972 15206
rect 5996 15204 6052 15206
rect 6076 15204 6132 15206
rect 6156 15204 6212 15206
rect 6236 15204 6292 15206
rect 6316 15204 6372 15206
rect 6396 15204 6452 15206
rect 6476 15204 6532 15206
rect 6556 15204 6612 15206
rect 6636 15204 6692 15206
rect 5630 15000 5686 15056
rect 6550 15036 6552 15056
rect 6552 15036 6604 15056
rect 6604 15036 6606 15056
rect 6550 15000 6606 15036
rect 5446 14592 5502 14648
rect 5538 14456 5594 14512
rect 5722 14728 5778 14784
rect 5630 14320 5686 14376
rect 6458 14728 6514 14784
rect 6274 14476 6330 14512
rect 6274 14456 6276 14476
rect 6276 14456 6328 14476
rect 6328 14456 6330 14476
rect 6642 14592 6698 14648
rect 5516 14170 5572 14172
rect 5596 14170 5652 14172
rect 5676 14170 5732 14172
rect 5756 14170 5812 14172
rect 5836 14170 5892 14172
rect 5916 14170 5972 14172
rect 5996 14170 6052 14172
rect 6076 14170 6132 14172
rect 6156 14170 6212 14172
rect 6236 14170 6292 14172
rect 6316 14170 6372 14172
rect 6396 14170 6452 14172
rect 6476 14170 6532 14172
rect 6556 14170 6612 14172
rect 6636 14170 6692 14172
rect 5516 14118 5554 14170
rect 5554 14118 5566 14170
rect 5566 14118 5572 14170
rect 5596 14118 5618 14170
rect 5618 14118 5630 14170
rect 5630 14118 5652 14170
rect 5676 14118 5682 14170
rect 5682 14118 5694 14170
rect 5694 14118 5732 14170
rect 5756 14118 5758 14170
rect 5758 14118 5810 14170
rect 5810 14118 5812 14170
rect 5836 14118 5874 14170
rect 5874 14118 5886 14170
rect 5886 14118 5892 14170
rect 5916 14118 5938 14170
rect 5938 14118 5950 14170
rect 5950 14118 5972 14170
rect 5996 14118 6002 14170
rect 6002 14118 6014 14170
rect 6014 14118 6052 14170
rect 6076 14118 6078 14170
rect 6078 14118 6130 14170
rect 6130 14118 6132 14170
rect 6156 14118 6194 14170
rect 6194 14118 6206 14170
rect 6206 14118 6212 14170
rect 6236 14118 6258 14170
rect 6258 14118 6270 14170
rect 6270 14118 6292 14170
rect 6316 14118 6322 14170
rect 6322 14118 6334 14170
rect 6334 14118 6372 14170
rect 6396 14118 6398 14170
rect 6398 14118 6450 14170
rect 6450 14118 6452 14170
rect 6476 14118 6514 14170
rect 6514 14118 6526 14170
rect 6526 14118 6532 14170
rect 6556 14118 6578 14170
rect 6578 14118 6590 14170
rect 6590 14118 6612 14170
rect 6636 14118 6642 14170
rect 6642 14118 6654 14170
rect 6654 14118 6692 14170
rect 5516 14116 5572 14118
rect 5596 14116 5652 14118
rect 5676 14116 5732 14118
rect 5756 14116 5812 14118
rect 5836 14116 5892 14118
rect 5916 14116 5972 14118
rect 5996 14116 6052 14118
rect 6076 14116 6132 14118
rect 6156 14116 6212 14118
rect 6236 14116 6292 14118
rect 6316 14116 6372 14118
rect 6396 14116 6452 14118
rect 6476 14116 6532 14118
rect 6556 14116 6612 14118
rect 6636 14116 6692 14118
rect 5538 13524 5594 13560
rect 5538 13504 5540 13524
rect 5540 13504 5592 13524
rect 5592 13504 5594 13524
rect 5170 13232 5226 13288
rect 4986 12960 5042 13016
rect 4894 12824 4950 12880
rect 4894 12436 4950 12472
rect 4894 12416 4896 12436
rect 4896 12416 4948 12436
rect 4948 12416 4950 12436
rect 5906 13504 5962 13560
rect 5722 13232 5778 13288
rect 6642 13268 6644 13288
rect 6644 13268 6696 13288
rect 6696 13268 6698 13288
rect 6642 13232 6698 13268
rect 5170 12960 5226 13016
rect 5516 13082 5572 13084
rect 5596 13082 5652 13084
rect 5676 13082 5732 13084
rect 5756 13082 5812 13084
rect 5836 13082 5892 13084
rect 5916 13082 5972 13084
rect 5996 13082 6052 13084
rect 6076 13082 6132 13084
rect 6156 13082 6212 13084
rect 6236 13082 6292 13084
rect 6316 13082 6372 13084
rect 6396 13082 6452 13084
rect 6476 13082 6532 13084
rect 6556 13082 6612 13084
rect 6636 13082 6692 13084
rect 5516 13030 5554 13082
rect 5554 13030 5566 13082
rect 5566 13030 5572 13082
rect 5596 13030 5618 13082
rect 5618 13030 5630 13082
rect 5630 13030 5652 13082
rect 5676 13030 5682 13082
rect 5682 13030 5694 13082
rect 5694 13030 5732 13082
rect 5756 13030 5758 13082
rect 5758 13030 5810 13082
rect 5810 13030 5812 13082
rect 5836 13030 5874 13082
rect 5874 13030 5886 13082
rect 5886 13030 5892 13082
rect 5916 13030 5938 13082
rect 5938 13030 5950 13082
rect 5950 13030 5972 13082
rect 5996 13030 6002 13082
rect 6002 13030 6014 13082
rect 6014 13030 6052 13082
rect 6076 13030 6078 13082
rect 6078 13030 6130 13082
rect 6130 13030 6132 13082
rect 6156 13030 6194 13082
rect 6194 13030 6206 13082
rect 6206 13030 6212 13082
rect 6236 13030 6258 13082
rect 6258 13030 6270 13082
rect 6270 13030 6292 13082
rect 6316 13030 6322 13082
rect 6322 13030 6334 13082
rect 6334 13030 6372 13082
rect 6396 13030 6398 13082
rect 6398 13030 6450 13082
rect 6450 13030 6452 13082
rect 6476 13030 6514 13082
rect 6514 13030 6526 13082
rect 6526 13030 6532 13082
rect 6556 13030 6578 13082
rect 6578 13030 6590 13082
rect 6590 13030 6612 13082
rect 6636 13030 6642 13082
rect 6642 13030 6654 13082
rect 6654 13030 6692 13082
rect 5516 13028 5572 13030
rect 5596 13028 5652 13030
rect 5676 13028 5732 13030
rect 5756 13028 5812 13030
rect 5836 13028 5892 13030
rect 5916 13028 5972 13030
rect 5996 13028 6052 13030
rect 6076 13028 6132 13030
rect 6156 13028 6212 13030
rect 6236 13028 6292 13030
rect 6316 13028 6372 13030
rect 6396 13028 6452 13030
rect 6476 13028 6532 13030
rect 6556 13028 6612 13030
rect 6636 13028 6692 13030
rect 4894 11464 4950 11520
rect 4618 10920 4674 10976
rect 5262 12280 5318 12336
rect 4986 9968 5042 10024
rect 5814 12824 5870 12880
rect 5722 12688 5778 12744
rect 5446 12280 5502 12336
rect 5630 12316 5632 12336
rect 5632 12316 5684 12336
rect 5684 12316 5686 12336
rect 5630 12280 5686 12316
rect 5998 12416 6054 12472
rect 6550 12824 6606 12880
rect 7194 15680 7250 15736
rect 6918 14456 6974 14512
rect 6826 13640 6882 13696
rect 6826 12688 6882 12744
rect 6182 12280 6238 12336
rect 6458 12144 6514 12200
rect 6642 12144 6698 12200
rect 5262 11620 5318 11656
rect 5262 11600 5264 11620
rect 5264 11600 5316 11620
rect 5316 11600 5318 11620
rect 5078 9560 5134 9616
rect 5262 10648 5318 10704
rect 5516 11994 5572 11996
rect 5596 11994 5652 11996
rect 5676 11994 5732 11996
rect 5756 11994 5812 11996
rect 5836 11994 5892 11996
rect 5916 11994 5972 11996
rect 5996 11994 6052 11996
rect 6076 11994 6132 11996
rect 6156 11994 6212 11996
rect 6236 11994 6292 11996
rect 6316 11994 6372 11996
rect 6396 11994 6452 11996
rect 6476 11994 6532 11996
rect 6556 11994 6612 11996
rect 6636 11994 6692 11996
rect 5516 11942 5554 11994
rect 5554 11942 5566 11994
rect 5566 11942 5572 11994
rect 5596 11942 5618 11994
rect 5618 11942 5630 11994
rect 5630 11942 5652 11994
rect 5676 11942 5682 11994
rect 5682 11942 5694 11994
rect 5694 11942 5732 11994
rect 5756 11942 5758 11994
rect 5758 11942 5810 11994
rect 5810 11942 5812 11994
rect 5836 11942 5874 11994
rect 5874 11942 5886 11994
rect 5886 11942 5892 11994
rect 5916 11942 5938 11994
rect 5938 11942 5950 11994
rect 5950 11942 5972 11994
rect 5996 11942 6002 11994
rect 6002 11942 6014 11994
rect 6014 11942 6052 11994
rect 6076 11942 6078 11994
rect 6078 11942 6130 11994
rect 6130 11942 6132 11994
rect 6156 11942 6194 11994
rect 6194 11942 6206 11994
rect 6206 11942 6212 11994
rect 6236 11942 6258 11994
rect 6258 11942 6270 11994
rect 6270 11942 6292 11994
rect 6316 11942 6322 11994
rect 6322 11942 6334 11994
rect 6334 11942 6372 11994
rect 6396 11942 6398 11994
rect 6398 11942 6450 11994
rect 6450 11942 6452 11994
rect 6476 11942 6514 11994
rect 6514 11942 6526 11994
rect 6526 11942 6532 11994
rect 6556 11942 6578 11994
rect 6578 11942 6590 11994
rect 6590 11942 6612 11994
rect 6636 11942 6642 11994
rect 6642 11942 6654 11994
rect 6654 11942 6692 11994
rect 5516 11940 5572 11942
rect 5596 11940 5652 11942
rect 5676 11940 5732 11942
rect 5756 11940 5812 11942
rect 5836 11940 5892 11942
rect 5916 11940 5972 11942
rect 5996 11940 6052 11942
rect 6076 11940 6132 11942
rect 6156 11940 6212 11942
rect 6236 11940 6292 11942
rect 6316 11940 6372 11942
rect 6396 11940 6452 11942
rect 6476 11940 6532 11942
rect 6556 11940 6612 11942
rect 6636 11940 6692 11942
rect 5630 11756 5686 11792
rect 5630 11736 5632 11756
rect 5632 11736 5684 11756
rect 5684 11736 5686 11756
rect 5814 11464 5870 11520
rect 5998 11328 6054 11384
rect 6550 11464 6606 11520
rect 6918 12280 6974 12336
rect 6826 11736 6882 11792
rect 7010 12008 7066 12064
rect 5516 10906 5572 10908
rect 5596 10906 5652 10908
rect 5676 10906 5732 10908
rect 5756 10906 5812 10908
rect 5836 10906 5892 10908
rect 5916 10906 5972 10908
rect 5996 10906 6052 10908
rect 6076 10906 6132 10908
rect 6156 10906 6212 10908
rect 6236 10906 6292 10908
rect 6316 10906 6372 10908
rect 6396 10906 6452 10908
rect 6476 10906 6532 10908
rect 6556 10906 6612 10908
rect 6636 10906 6692 10908
rect 5516 10854 5554 10906
rect 5554 10854 5566 10906
rect 5566 10854 5572 10906
rect 5596 10854 5618 10906
rect 5618 10854 5630 10906
rect 5630 10854 5652 10906
rect 5676 10854 5682 10906
rect 5682 10854 5694 10906
rect 5694 10854 5732 10906
rect 5756 10854 5758 10906
rect 5758 10854 5810 10906
rect 5810 10854 5812 10906
rect 5836 10854 5874 10906
rect 5874 10854 5886 10906
rect 5886 10854 5892 10906
rect 5916 10854 5938 10906
rect 5938 10854 5950 10906
rect 5950 10854 5972 10906
rect 5996 10854 6002 10906
rect 6002 10854 6014 10906
rect 6014 10854 6052 10906
rect 6076 10854 6078 10906
rect 6078 10854 6130 10906
rect 6130 10854 6132 10906
rect 6156 10854 6194 10906
rect 6194 10854 6206 10906
rect 6206 10854 6212 10906
rect 6236 10854 6258 10906
rect 6258 10854 6270 10906
rect 6270 10854 6292 10906
rect 6316 10854 6322 10906
rect 6322 10854 6334 10906
rect 6334 10854 6372 10906
rect 6396 10854 6398 10906
rect 6398 10854 6450 10906
rect 6450 10854 6452 10906
rect 6476 10854 6514 10906
rect 6514 10854 6526 10906
rect 6526 10854 6532 10906
rect 6556 10854 6578 10906
rect 6578 10854 6590 10906
rect 6590 10854 6612 10906
rect 6636 10854 6642 10906
rect 6642 10854 6654 10906
rect 6654 10854 6692 10906
rect 5516 10852 5572 10854
rect 5596 10852 5652 10854
rect 5676 10852 5732 10854
rect 5756 10852 5812 10854
rect 5836 10852 5892 10854
rect 5916 10852 5972 10854
rect 5996 10852 6052 10854
rect 6076 10852 6132 10854
rect 6156 10852 6212 10854
rect 6236 10852 6292 10854
rect 6316 10852 6372 10854
rect 6396 10852 6452 10854
rect 6476 10852 6532 10854
rect 6556 10852 6612 10854
rect 6636 10852 6692 10854
rect 5538 10548 5540 10568
rect 5540 10548 5592 10568
rect 5592 10548 5594 10568
rect 5538 10512 5594 10548
rect 6550 10240 6606 10296
rect 6642 9968 6698 10024
rect 5516 9818 5572 9820
rect 5596 9818 5652 9820
rect 5676 9818 5732 9820
rect 5756 9818 5812 9820
rect 5836 9818 5892 9820
rect 5916 9818 5972 9820
rect 5996 9818 6052 9820
rect 6076 9818 6132 9820
rect 6156 9818 6212 9820
rect 6236 9818 6292 9820
rect 6316 9818 6372 9820
rect 6396 9818 6452 9820
rect 6476 9818 6532 9820
rect 6556 9818 6612 9820
rect 6636 9818 6692 9820
rect 5516 9766 5554 9818
rect 5554 9766 5566 9818
rect 5566 9766 5572 9818
rect 5596 9766 5618 9818
rect 5618 9766 5630 9818
rect 5630 9766 5652 9818
rect 5676 9766 5682 9818
rect 5682 9766 5694 9818
rect 5694 9766 5732 9818
rect 5756 9766 5758 9818
rect 5758 9766 5810 9818
rect 5810 9766 5812 9818
rect 5836 9766 5874 9818
rect 5874 9766 5886 9818
rect 5886 9766 5892 9818
rect 5916 9766 5938 9818
rect 5938 9766 5950 9818
rect 5950 9766 5972 9818
rect 5996 9766 6002 9818
rect 6002 9766 6014 9818
rect 6014 9766 6052 9818
rect 6076 9766 6078 9818
rect 6078 9766 6130 9818
rect 6130 9766 6132 9818
rect 6156 9766 6194 9818
rect 6194 9766 6206 9818
rect 6206 9766 6212 9818
rect 6236 9766 6258 9818
rect 6258 9766 6270 9818
rect 6270 9766 6292 9818
rect 6316 9766 6322 9818
rect 6322 9766 6334 9818
rect 6334 9766 6372 9818
rect 6396 9766 6398 9818
rect 6398 9766 6450 9818
rect 6450 9766 6452 9818
rect 6476 9766 6514 9818
rect 6514 9766 6526 9818
rect 6526 9766 6532 9818
rect 6556 9766 6578 9818
rect 6578 9766 6590 9818
rect 6590 9766 6612 9818
rect 6636 9766 6642 9818
rect 6642 9766 6654 9818
rect 6654 9766 6692 9818
rect 5516 9764 5572 9766
rect 5596 9764 5652 9766
rect 5676 9764 5732 9766
rect 5756 9764 5812 9766
rect 5836 9764 5892 9766
rect 5916 9764 5972 9766
rect 5996 9764 6052 9766
rect 6076 9764 6132 9766
rect 6156 9764 6212 9766
rect 6236 9764 6292 9766
rect 6316 9764 6372 9766
rect 6396 9764 6452 9766
rect 6476 9764 6532 9766
rect 6556 9764 6612 9766
rect 6636 9764 6692 9766
rect 5516 8730 5572 8732
rect 5596 8730 5652 8732
rect 5676 8730 5732 8732
rect 5756 8730 5812 8732
rect 5836 8730 5892 8732
rect 5916 8730 5972 8732
rect 5996 8730 6052 8732
rect 6076 8730 6132 8732
rect 6156 8730 6212 8732
rect 6236 8730 6292 8732
rect 6316 8730 6372 8732
rect 6396 8730 6452 8732
rect 6476 8730 6532 8732
rect 6556 8730 6612 8732
rect 6636 8730 6692 8732
rect 5516 8678 5554 8730
rect 5554 8678 5566 8730
rect 5566 8678 5572 8730
rect 5596 8678 5618 8730
rect 5618 8678 5630 8730
rect 5630 8678 5652 8730
rect 5676 8678 5682 8730
rect 5682 8678 5694 8730
rect 5694 8678 5732 8730
rect 5756 8678 5758 8730
rect 5758 8678 5810 8730
rect 5810 8678 5812 8730
rect 5836 8678 5874 8730
rect 5874 8678 5886 8730
rect 5886 8678 5892 8730
rect 5916 8678 5938 8730
rect 5938 8678 5950 8730
rect 5950 8678 5972 8730
rect 5996 8678 6002 8730
rect 6002 8678 6014 8730
rect 6014 8678 6052 8730
rect 6076 8678 6078 8730
rect 6078 8678 6130 8730
rect 6130 8678 6132 8730
rect 6156 8678 6194 8730
rect 6194 8678 6206 8730
rect 6206 8678 6212 8730
rect 6236 8678 6258 8730
rect 6258 8678 6270 8730
rect 6270 8678 6292 8730
rect 6316 8678 6322 8730
rect 6322 8678 6334 8730
rect 6334 8678 6372 8730
rect 6396 8678 6398 8730
rect 6398 8678 6450 8730
rect 6450 8678 6452 8730
rect 6476 8678 6514 8730
rect 6514 8678 6526 8730
rect 6526 8678 6532 8730
rect 6556 8678 6578 8730
rect 6578 8678 6590 8730
rect 6590 8678 6612 8730
rect 6636 8678 6642 8730
rect 6642 8678 6654 8730
rect 6654 8678 6692 8730
rect 5516 8676 5572 8678
rect 5596 8676 5652 8678
rect 5676 8676 5732 8678
rect 5756 8676 5812 8678
rect 5836 8676 5892 8678
rect 5916 8676 5972 8678
rect 5996 8676 6052 8678
rect 6076 8676 6132 8678
rect 6156 8676 6212 8678
rect 6236 8676 6292 8678
rect 6316 8676 6372 8678
rect 6396 8676 6452 8678
rect 6476 8676 6532 8678
rect 6556 8676 6612 8678
rect 6636 8676 6692 8678
rect 5446 8336 5502 8392
rect 5516 7642 5572 7644
rect 5596 7642 5652 7644
rect 5676 7642 5732 7644
rect 5756 7642 5812 7644
rect 5836 7642 5892 7644
rect 5916 7642 5972 7644
rect 5996 7642 6052 7644
rect 6076 7642 6132 7644
rect 6156 7642 6212 7644
rect 6236 7642 6292 7644
rect 6316 7642 6372 7644
rect 6396 7642 6452 7644
rect 6476 7642 6532 7644
rect 6556 7642 6612 7644
rect 6636 7642 6692 7644
rect 5516 7590 5554 7642
rect 5554 7590 5566 7642
rect 5566 7590 5572 7642
rect 5596 7590 5618 7642
rect 5618 7590 5630 7642
rect 5630 7590 5652 7642
rect 5676 7590 5682 7642
rect 5682 7590 5694 7642
rect 5694 7590 5732 7642
rect 5756 7590 5758 7642
rect 5758 7590 5810 7642
rect 5810 7590 5812 7642
rect 5836 7590 5874 7642
rect 5874 7590 5886 7642
rect 5886 7590 5892 7642
rect 5916 7590 5938 7642
rect 5938 7590 5950 7642
rect 5950 7590 5972 7642
rect 5996 7590 6002 7642
rect 6002 7590 6014 7642
rect 6014 7590 6052 7642
rect 6076 7590 6078 7642
rect 6078 7590 6130 7642
rect 6130 7590 6132 7642
rect 6156 7590 6194 7642
rect 6194 7590 6206 7642
rect 6206 7590 6212 7642
rect 6236 7590 6258 7642
rect 6258 7590 6270 7642
rect 6270 7590 6292 7642
rect 6316 7590 6322 7642
rect 6322 7590 6334 7642
rect 6334 7590 6372 7642
rect 6396 7590 6398 7642
rect 6398 7590 6450 7642
rect 6450 7590 6452 7642
rect 6476 7590 6514 7642
rect 6514 7590 6526 7642
rect 6526 7590 6532 7642
rect 6556 7590 6578 7642
rect 6578 7590 6590 7642
rect 6590 7590 6612 7642
rect 6636 7590 6642 7642
rect 6642 7590 6654 7642
rect 6654 7590 6692 7642
rect 5516 7588 5572 7590
rect 5596 7588 5652 7590
rect 5676 7588 5732 7590
rect 5756 7588 5812 7590
rect 5836 7588 5892 7590
rect 5916 7588 5972 7590
rect 5996 7588 6052 7590
rect 6076 7588 6132 7590
rect 6156 7588 6212 7590
rect 6236 7588 6292 7590
rect 6316 7588 6372 7590
rect 6396 7588 6452 7590
rect 6476 7588 6532 7590
rect 6556 7588 6612 7590
rect 6636 7588 6692 7590
rect 5722 7384 5778 7440
rect 5538 7284 5540 7304
rect 5540 7284 5592 7304
rect 5592 7284 5594 7304
rect 5538 7248 5594 7284
rect 5516 6554 5572 6556
rect 5596 6554 5652 6556
rect 5676 6554 5732 6556
rect 5756 6554 5812 6556
rect 5836 6554 5892 6556
rect 5916 6554 5972 6556
rect 5996 6554 6052 6556
rect 6076 6554 6132 6556
rect 6156 6554 6212 6556
rect 6236 6554 6292 6556
rect 6316 6554 6372 6556
rect 6396 6554 6452 6556
rect 6476 6554 6532 6556
rect 6556 6554 6612 6556
rect 6636 6554 6692 6556
rect 5516 6502 5554 6554
rect 5554 6502 5566 6554
rect 5566 6502 5572 6554
rect 5596 6502 5618 6554
rect 5618 6502 5630 6554
rect 5630 6502 5652 6554
rect 5676 6502 5682 6554
rect 5682 6502 5694 6554
rect 5694 6502 5732 6554
rect 5756 6502 5758 6554
rect 5758 6502 5810 6554
rect 5810 6502 5812 6554
rect 5836 6502 5874 6554
rect 5874 6502 5886 6554
rect 5886 6502 5892 6554
rect 5916 6502 5938 6554
rect 5938 6502 5950 6554
rect 5950 6502 5972 6554
rect 5996 6502 6002 6554
rect 6002 6502 6014 6554
rect 6014 6502 6052 6554
rect 6076 6502 6078 6554
rect 6078 6502 6130 6554
rect 6130 6502 6132 6554
rect 6156 6502 6194 6554
rect 6194 6502 6206 6554
rect 6206 6502 6212 6554
rect 6236 6502 6258 6554
rect 6258 6502 6270 6554
rect 6270 6502 6292 6554
rect 6316 6502 6322 6554
rect 6322 6502 6334 6554
rect 6334 6502 6372 6554
rect 6396 6502 6398 6554
rect 6398 6502 6450 6554
rect 6450 6502 6452 6554
rect 6476 6502 6514 6554
rect 6514 6502 6526 6554
rect 6526 6502 6532 6554
rect 6556 6502 6578 6554
rect 6578 6502 6590 6554
rect 6590 6502 6612 6554
rect 6636 6502 6642 6554
rect 6642 6502 6654 6554
rect 6654 6502 6692 6554
rect 5516 6500 5572 6502
rect 5596 6500 5652 6502
rect 5676 6500 5732 6502
rect 5756 6500 5812 6502
rect 5836 6500 5892 6502
rect 5916 6500 5972 6502
rect 5996 6500 6052 6502
rect 6076 6500 6132 6502
rect 6156 6500 6212 6502
rect 6236 6500 6292 6502
rect 6316 6500 6372 6502
rect 6396 6500 6452 6502
rect 6476 6500 6532 6502
rect 6556 6500 6612 6502
rect 6636 6500 6692 6502
rect 5354 6160 5410 6216
rect 5516 5466 5572 5468
rect 5596 5466 5652 5468
rect 5676 5466 5732 5468
rect 5756 5466 5812 5468
rect 5836 5466 5892 5468
rect 5916 5466 5972 5468
rect 5996 5466 6052 5468
rect 6076 5466 6132 5468
rect 6156 5466 6212 5468
rect 6236 5466 6292 5468
rect 6316 5466 6372 5468
rect 6396 5466 6452 5468
rect 6476 5466 6532 5468
rect 6556 5466 6612 5468
rect 6636 5466 6692 5468
rect 5516 5414 5554 5466
rect 5554 5414 5566 5466
rect 5566 5414 5572 5466
rect 5596 5414 5618 5466
rect 5618 5414 5630 5466
rect 5630 5414 5652 5466
rect 5676 5414 5682 5466
rect 5682 5414 5694 5466
rect 5694 5414 5732 5466
rect 5756 5414 5758 5466
rect 5758 5414 5810 5466
rect 5810 5414 5812 5466
rect 5836 5414 5874 5466
rect 5874 5414 5886 5466
rect 5886 5414 5892 5466
rect 5916 5414 5938 5466
rect 5938 5414 5950 5466
rect 5950 5414 5972 5466
rect 5996 5414 6002 5466
rect 6002 5414 6014 5466
rect 6014 5414 6052 5466
rect 6076 5414 6078 5466
rect 6078 5414 6130 5466
rect 6130 5414 6132 5466
rect 6156 5414 6194 5466
rect 6194 5414 6206 5466
rect 6206 5414 6212 5466
rect 6236 5414 6258 5466
rect 6258 5414 6270 5466
rect 6270 5414 6292 5466
rect 6316 5414 6322 5466
rect 6322 5414 6334 5466
rect 6334 5414 6372 5466
rect 6396 5414 6398 5466
rect 6398 5414 6450 5466
rect 6450 5414 6452 5466
rect 6476 5414 6514 5466
rect 6514 5414 6526 5466
rect 6526 5414 6532 5466
rect 6556 5414 6578 5466
rect 6578 5414 6590 5466
rect 6590 5414 6612 5466
rect 6636 5414 6642 5466
rect 6642 5414 6654 5466
rect 6654 5414 6692 5466
rect 5516 5412 5572 5414
rect 5596 5412 5652 5414
rect 5676 5412 5732 5414
rect 5756 5412 5812 5414
rect 5836 5412 5892 5414
rect 5916 5412 5972 5414
rect 5996 5412 6052 5414
rect 6076 5412 6132 5414
rect 6156 5412 6212 5414
rect 6236 5412 6292 5414
rect 6316 5412 6372 5414
rect 6396 5412 6452 5414
rect 6476 5412 6532 5414
rect 6556 5412 6612 5414
rect 6636 5412 6692 5414
rect 6458 5228 6514 5264
rect 6458 5208 6460 5228
rect 6460 5208 6512 5228
rect 6512 5208 6514 5228
rect 7286 15136 7342 15192
rect 7654 15952 7710 16008
rect 7470 15272 7526 15328
rect 7378 14728 7434 14784
rect 7746 15408 7802 15464
rect 7654 14320 7710 14376
rect 7378 13232 7434 13288
rect 7194 12960 7250 13016
rect 7562 13096 7618 13152
rect 7286 12198 7342 12200
rect 7286 12146 7288 12198
rect 7288 12146 7340 12198
rect 7340 12146 7342 12198
rect 7286 12144 7342 12146
rect 7286 10920 7342 10976
rect 6826 6840 6882 6896
rect 5516 4378 5572 4380
rect 5596 4378 5652 4380
rect 5676 4378 5732 4380
rect 5756 4378 5812 4380
rect 5836 4378 5892 4380
rect 5916 4378 5972 4380
rect 5996 4378 6052 4380
rect 6076 4378 6132 4380
rect 6156 4378 6212 4380
rect 6236 4378 6292 4380
rect 6316 4378 6372 4380
rect 6396 4378 6452 4380
rect 6476 4378 6532 4380
rect 6556 4378 6612 4380
rect 6636 4378 6692 4380
rect 5516 4326 5554 4378
rect 5554 4326 5566 4378
rect 5566 4326 5572 4378
rect 5596 4326 5618 4378
rect 5618 4326 5630 4378
rect 5630 4326 5652 4378
rect 5676 4326 5682 4378
rect 5682 4326 5694 4378
rect 5694 4326 5732 4378
rect 5756 4326 5758 4378
rect 5758 4326 5810 4378
rect 5810 4326 5812 4378
rect 5836 4326 5874 4378
rect 5874 4326 5886 4378
rect 5886 4326 5892 4378
rect 5916 4326 5938 4378
rect 5938 4326 5950 4378
rect 5950 4326 5972 4378
rect 5996 4326 6002 4378
rect 6002 4326 6014 4378
rect 6014 4326 6052 4378
rect 6076 4326 6078 4378
rect 6078 4326 6130 4378
rect 6130 4326 6132 4378
rect 6156 4326 6194 4378
rect 6194 4326 6206 4378
rect 6206 4326 6212 4378
rect 6236 4326 6258 4378
rect 6258 4326 6270 4378
rect 6270 4326 6292 4378
rect 6316 4326 6322 4378
rect 6322 4326 6334 4378
rect 6334 4326 6372 4378
rect 6396 4326 6398 4378
rect 6398 4326 6450 4378
rect 6450 4326 6452 4378
rect 6476 4326 6514 4378
rect 6514 4326 6526 4378
rect 6526 4326 6532 4378
rect 6556 4326 6578 4378
rect 6578 4326 6590 4378
rect 6590 4326 6612 4378
rect 6636 4326 6642 4378
rect 6642 4326 6654 4378
rect 6654 4326 6692 4378
rect 5516 4324 5572 4326
rect 5596 4324 5652 4326
rect 5676 4324 5732 4326
rect 5756 4324 5812 4326
rect 5836 4324 5892 4326
rect 5916 4324 5972 4326
rect 5996 4324 6052 4326
rect 6076 4324 6132 4326
rect 6156 4324 6212 4326
rect 6236 4324 6292 4326
rect 6316 4324 6372 4326
rect 6396 4324 6452 4326
rect 6476 4324 6532 4326
rect 6556 4324 6612 4326
rect 6636 4324 6692 4326
rect 5722 3576 5778 3632
rect 3514 1028 3516 1048
rect 3516 1028 3568 1048
rect 3568 1028 3570 1048
rect 3514 992 3570 1028
rect 3422 448 3478 504
rect 4066 176 4122 232
rect 5516 3290 5572 3292
rect 5596 3290 5652 3292
rect 5676 3290 5732 3292
rect 5756 3290 5812 3292
rect 5836 3290 5892 3292
rect 5916 3290 5972 3292
rect 5996 3290 6052 3292
rect 6076 3290 6132 3292
rect 6156 3290 6212 3292
rect 6236 3290 6292 3292
rect 6316 3290 6372 3292
rect 6396 3290 6452 3292
rect 6476 3290 6532 3292
rect 6556 3290 6612 3292
rect 6636 3290 6692 3292
rect 5516 3238 5554 3290
rect 5554 3238 5566 3290
rect 5566 3238 5572 3290
rect 5596 3238 5618 3290
rect 5618 3238 5630 3290
rect 5630 3238 5652 3290
rect 5676 3238 5682 3290
rect 5682 3238 5694 3290
rect 5694 3238 5732 3290
rect 5756 3238 5758 3290
rect 5758 3238 5810 3290
rect 5810 3238 5812 3290
rect 5836 3238 5874 3290
rect 5874 3238 5886 3290
rect 5886 3238 5892 3290
rect 5916 3238 5938 3290
rect 5938 3238 5950 3290
rect 5950 3238 5972 3290
rect 5996 3238 6002 3290
rect 6002 3238 6014 3290
rect 6014 3238 6052 3290
rect 6076 3238 6078 3290
rect 6078 3238 6130 3290
rect 6130 3238 6132 3290
rect 6156 3238 6194 3290
rect 6194 3238 6206 3290
rect 6206 3238 6212 3290
rect 6236 3238 6258 3290
rect 6258 3238 6270 3290
rect 6270 3238 6292 3290
rect 6316 3238 6322 3290
rect 6322 3238 6334 3290
rect 6334 3238 6372 3290
rect 6396 3238 6398 3290
rect 6398 3238 6450 3290
rect 6450 3238 6452 3290
rect 6476 3238 6514 3290
rect 6514 3238 6526 3290
rect 6526 3238 6532 3290
rect 6556 3238 6578 3290
rect 6578 3238 6590 3290
rect 6590 3238 6612 3290
rect 6636 3238 6642 3290
rect 6642 3238 6654 3290
rect 6654 3238 6692 3290
rect 5516 3236 5572 3238
rect 5596 3236 5652 3238
rect 5676 3236 5732 3238
rect 5756 3236 5812 3238
rect 5836 3236 5892 3238
rect 5916 3236 5972 3238
rect 5996 3236 6052 3238
rect 6076 3236 6132 3238
rect 6156 3236 6212 3238
rect 6236 3236 6292 3238
rect 6316 3236 6372 3238
rect 6396 3236 6452 3238
rect 6476 3236 6532 3238
rect 6556 3236 6612 3238
rect 6636 3236 6692 3238
rect 7102 10240 7158 10296
rect 7102 8608 7158 8664
rect 13516 17434 13572 17436
rect 13596 17434 13652 17436
rect 13676 17434 13732 17436
rect 13756 17434 13812 17436
rect 13836 17434 13892 17436
rect 13916 17434 13972 17436
rect 13996 17434 14052 17436
rect 14076 17434 14132 17436
rect 14156 17434 14212 17436
rect 14236 17434 14292 17436
rect 14316 17434 14372 17436
rect 14396 17434 14452 17436
rect 14476 17434 14532 17436
rect 14556 17434 14612 17436
rect 14636 17434 14692 17436
rect 13516 17382 13554 17434
rect 13554 17382 13566 17434
rect 13566 17382 13572 17434
rect 13596 17382 13618 17434
rect 13618 17382 13630 17434
rect 13630 17382 13652 17434
rect 13676 17382 13682 17434
rect 13682 17382 13694 17434
rect 13694 17382 13732 17434
rect 13756 17382 13758 17434
rect 13758 17382 13810 17434
rect 13810 17382 13812 17434
rect 13836 17382 13874 17434
rect 13874 17382 13886 17434
rect 13886 17382 13892 17434
rect 13916 17382 13938 17434
rect 13938 17382 13950 17434
rect 13950 17382 13972 17434
rect 13996 17382 14002 17434
rect 14002 17382 14014 17434
rect 14014 17382 14052 17434
rect 14076 17382 14078 17434
rect 14078 17382 14130 17434
rect 14130 17382 14132 17434
rect 14156 17382 14194 17434
rect 14194 17382 14206 17434
rect 14206 17382 14212 17434
rect 14236 17382 14258 17434
rect 14258 17382 14270 17434
rect 14270 17382 14292 17434
rect 14316 17382 14322 17434
rect 14322 17382 14334 17434
rect 14334 17382 14372 17434
rect 14396 17382 14398 17434
rect 14398 17382 14450 17434
rect 14450 17382 14452 17434
rect 14476 17382 14514 17434
rect 14514 17382 14526 17434
rect 14526 17382 14532 17434
rect 14556 17382 14578 17434
rect 14578 17382 14590 17434
rect 14590 17382 14612 17434
rect 14636 17382 14642 17434
rect 14642 17382 14654 17434
rect 14654 17382 14692 17434
rect 13516 17380 13572 17382
rect 13596 17380 13652 17382
rect 13676 17380 13732 17382
rect 13756 17380 13812 17382
rect 13836 17380 13892 17382
rect 13916 17380 13972 17382
rect 13996 17380 14052 17382
rect 14076 17380 14132 17382
rect 14156 17380 14212 17382
rect 14236 17380 14292 17382
rect 14316 17380 14372 17382
rect 14396 17380 14452 17382
rect 14476 17380 14532 17382
rect 14556 17380 14612 17382
rect 14636 17380 14692 17382
rect 10874 17176 10930 17232
rect 7746 12280 7802 12336
rect 7654 11872 7710 11928
rect 8022 13504 8078 13560
rect 8206 13776 8262 13832
rect 8206 13232 8262 13288
rect 8114 12688 8170 12744
rect 7930 12144 7986 12200
rect 7654 11600 7710 11656
rect 8114 11872 8170 11928
rect 7378 8472 7434 8528
rect 7562 10240 7618 10296
rect 7470 7384 7526 7440
rect 7838 10920 7894 10976
rect 8482 11600 8538 11656
rect 8758 13504 8814 13560
rect 8666 12688 8722 12744
rect 8666 12280 8722 12336
rect 8206 11192 8262 11248
rect 8114 11056 8170 11112
rect 8022 10920 8078 10976
rect 7930 10784 7986 10840
rect 7838 10376 7894 10432
rect 7746 10240 7802 10296
rect 7746 10104 7802 10160
rect 7838 9424 7894 9480
rect 7746 8472 7802 8528
rect 8206 10376 8262 10432
rect 8114 10104 8170 10160
rect 8022 9560 8078 9616
rect 8390 11328 8446 11384
rect 7746 3984 7802 4040
rect 5516 2202 5572 2204
rect 5596 2202 5652 2204
rect 5676 2202 5732 2204
rect 5756 2202 5812 2204
rect 5836 2202 5892 2204
rect 5916 2202 5972 2204
rect 5996 2202 6052 2204
rect 6076 2202 6132 2204
rect 6156 2202 6212 2204
rect 6236 2202 6292 2204
rect 6316 2202 6372 2204
rect 6396 2202 6452 2204
rect 6476 2202 6532 2204
rect 6556 2202 6612 2204
rect 6636 2202 6692 2204
rect 5516 2150 5554 2202
rect 5554 2150 5566 2202
rect 5566 2150 5572 2202
rect 5596 2150 5618 2202
rect 5618 2150 5630 2202
rect 5630 2150 5652 2202
rect 5676 2150 5682 2202
rect 5682 2150 5694 2202
rect 5694 2150 5732 2202
rect 5756 2150 5758 2202
rect 5758 2150 5810 2202
rect 5810 2150 5812 2202
rect 5836 2150 5874 2202
rect 5874 2150 5886 2202
rect 5886 2150 5892 2202
rect 5916 2150 5938 2202
rect 5938 2150 5950 2202
rect 5950 2150 5972 2202
rect 5996 2150 6002 2202
rect 6002 2150 6014 2202
rect 6014 2150 6052 2202
rect 6076 2150 6078 2202
rect 6078 2150 6130 2202
rect 6130 2150 6132 2202
rect 6156 2150 6194 2202
rect 6194 2150 6206 2202
rect 6206 2150 6212 2202
rect 6236 2150 6258 2202
rect 6258 2150 6270 2202
rect 6270 2150 6292 2202
rect 6316 2150 6322 2202
rect 6322 2150 6334 2202
rect 6334 2150 6372 2202
rect 6396 2150 6398 2202
rect 6398 2150 6450 2202
rect 6450 2150 6452 2202
rect 6476 2150 6514 2202
rect 6514 2150 6526 2202
rect 6526 2150 6532 2202
rect 6556 2150 6578 2202
rect 6578 2150 6590 2202
rect 6590 2150 6612 2202
rect 6636 2150 6642 2202
rect 6642 2150 6654 2202
rect 6654 2150 6692 2202
rect 5516 2148 5572 2150
rect 5596 2148 5652 2150
rect 5676 2148 5732 2150
rect 5756 2148 5812 2150
rect 5836 2148 5892 2150
rect 5916 2148 5972 2150
rect 5996 2148 6052 2150
rect 6076 2148 6132 2150
rect 6156 2148 6212 2150
rect 6236 2148 6292 2150
rect 6316 2148 6372 2150
rect 6396 2148 6452 2150
rect 6476 2148 6532 2150
rect 6556 2148 6612 2150
rect 6636 2148 6692 2150
rect 8574 11212 8630 11248
rect 8574 11192 8576 11212
rect 8576 11192 8628 11212
rect 8628 11192 8630 11212
rect 8482 11056 8538 11112
rect 9516 16890 9572 16892
rect 9596 16890 9652 16892
rect 9676 16890 9732 16892
rect 9756 16890 9812 16892
rect 9836 16890 9892 16892
rect 9916 16890 9972 16892
rect 9996 16890 10052 16892
rect 10076 16890 10132 16892
rect 10156 16890 10212 16892
rect 10236 16890 10292 16892
rect 10316 16890 10372 16892
rect 10396 16890 10452 16892
rect 10476 16890 10532 16892
rect 10556 16890 10612 16892
rect 10636 16890 10692 16892
rect 9516 16838 9554 16890
rect 9554 16838 9566 16890
rect 9566 16838 9572 16890
rect 9596 16838 9618 16890
rect 9618 16838 9630 16890
rect 9630 16838 9652 16890
rect 9676 16838 9682 16890
rect 9682 16838 9694 16890
rect 9694 16838 9732 16890
rect 9756 16838 9758 16890
rect 9758 16838 9810 16890
rect 9810 16838 9812 16890
rect 9836 16838 9874 16890
rect 9874 16838 9886 16890
rect 9886 16838 9892 16890
rect 9916 16838 9938 16890
rect 9938 16838 9950 16890
rect 9950 16838 9972 16890
rect 9996 16838 10002 16890
rect 10002 16838 10014 16890
rect 10014 16838 10052 16890
rect 10076 16838 10078 16890
rect 10078 16838 10130 16890
rect 10130 16838 10132 16890
rect 10156 16838 10194 16890
rect 10194 16838 10206 16890
rect 10206 16838 10212 16890
rect 10236 16838 10258 16890
rect 10258 16838 10270 16890
rect 10270 16838 10292 16890
rect 10316 16838 10322 16890
rect 10322 16838 10334 16890
rect 10334 16838 10372 16890
rect 10396 16838 10398 16890
rect 10398 16838 10450 16890
rect 10450 16838 10452 16890
rect 10476 16838 10514 16890
rect 10514 16838 10526 16890
rect 10526 16838 10532 16890
rect 10556 16838 10578 16890
rect 10578 16838 10590 16890
rect 10590 16838 10612 16890
rect 10636 16838 10642 16890
rect 10642 16838 10654 16890
rect 10654 16838 10692 16890
rect 9516 16836 9572 16838
rect 9596 16836 9652 16838
rect 9676 16836 9732 16838
rect 9756 16836 9812 16838
rect 9836 16836 9892 16838
rect 9916 16836 9972 16838
rect 9996 16836 10052 16838
rect 10076 16836 10132 16838
rect 10156 16836 10212 16838
rect 10236 16836 10292 16838
rect 10316 16836 10372 16838
rect 10396 16836 10452 16838
rect 10476 16836 10532 16838
rect 10556 16836 10612 16838
rect 10636 16836 10692 16838
rect 9516 15802 9572 15804
rect 9596 15802 9652 15804
rect 9676 15802 9732 15804
rect 9756 15802 9812 15804
rect 9836 15802 9892 15804
rect 9916 15802 9972 15804
rect 9996 15802 10052 15804
rect 10076 15802 10132 15804
rect 10156 15802 10212 15804
rect 10236 15802 10292 15804
rect 10316 15802 10372 15804
rect 10396 15802 10452 15804
rect 10476 15802 10532 15804
rect 10556 15802 10612 15804
rect 10636 15802 10692 15804
rect 9516 15750 9554 15802
rect 9554 15750 9566 15802
rect 9566 15750 9572 15802
rect 9596 15750 9618 15802
rect 9618 15750 9630 15802
rect 9630 15750 9652 15802
rect 9676 15750 9682 15802
rect 9682 15750 9694 15802
rect 9694 15750 9732 15802
rect 9756 15750 9758 15802
rect 9758 15750 9810 15802
rect 9810 15750 9812 15802
rect 9836 15750 9874 15802
rect 9874 15750 9886 15802
rect 9886 15750 9892 15802
rect 9916 15750 9938 15802
rect 9938 15750 9950 15802
rect 9950 15750 9972 15802
rect 9996 15750 10002 15802
rect 10002 15750 10014 15802
rect 10014 15750 10052 15802
rect 10076 15750 10078 15802
rect 10078 15750 10130 15802
rect 10130 15750 10132 15802
rect 10156 15750 10194 15802
rect 10194 15750 10206 15802
rect 10206 15750 10212 15802
rect 10236 15750 10258 15802
rect 10258 15750 10270 15802
rect 10270 15750 10292 15802
rect 10316 15750 10322 15802
rect 10322 15750 10334 15802
rect 10334 15750 10372 15802
rect 10396 15750 10398 15802
rect 10398 15750 10450 15802
rect 10450 15750 10452 15802
rect 10476 15750 10514 15802
rect 10514 15750 10526 15802
rect 10526 15750 10532 15802
rect 10556 15750 10578 15802
rect 10578 15750 10590 15802
rect 10590 15750 10612 15802
rect 10636 15750 10642 15802
rect 10642 15750 10654 15802
rect 10654 15750 10692 15802
rect 9516 15748 9572 15750
rect 9596 15748 9652 15750
rect 9676 15748 9732 15750
rect 9756 15748 9812 15750
rect 9836 15748 9892 15750
rect 9916 15748 9972 15750
rect 9996 15748 10052 15750
rect 10076 15748 10132 15750
rect 10156 15748 10212 15750
rect 10236 15748 10292 15750
rect 10316 15748 10372 15750
rect 10396 15748 10452 15750
rect 10476 15748 10532 15750
rect 10556 15748 10612 15750
rect 10636 15748 10692 15750
rect 9034 14048 9090 14104
rect 9034 12144 9090 12200
rect 9126 11872 9182 11928
rect 9402 14884 9458 14920
rect 9402 14864 9404 14884
rect 9404 14864 9456 14884
rect 9456 14864 9458 14884
rect 9516 14714 9572 14716
rect 9596 14714 9652 14716
rect 9676 14714 9732 14716
rect 9756 14714 9812 14716
rect 9836 14714 9892 14716
rect 9916 14714 9972 14716
rect 9996 14714 10052 14716
rect 10076 14714 10132 14716
rect 10156 14714 10212 14716
rect 10236 14714 10292 14716
rect 10316 14714 10372 14716
rect 10396 14714 10452 14716
rect 10476 14714 10532 14716
rect 10556 14714 10612 14716
rect 10636 14714 10692 14716
rect 9516 14662 9554 14714
rect 9554 14662 9566 14714
rect 9566 14662 9572 14714
rect 9596 14662 9618 14714
rect 9618 14662 9630 14714
rect 9630 14662 9652 14714
rect 9676 14662 9682 14714
rect 9682 14662 9694 14714
rect 9694 14662 9732 14714
rect 9756 14662 9758 14714
rect 9758 14662 9810 14714
rect 9810 14662 9812 14714
rect 9836 14662 9874 14714
rect 9874 14662 9886 14714
rect 9886 14662 9892 14714
rect 9916 14662 9938 14714
rect 9938 14662 9950 14714
rect 9950 14662 9972 14714
rect 9996 14662 10002 14714
rect 10002 14662 10014 14714
rect 10014 14662 10052 14714
rect 10076 14662 10078 14714
rect 10078 14662 10130 14714
rect 10130 14662 10132 14714
rect 10156 14662 10194 14714
rect 10194 14662 10206 14714
rect 10206 14662 10212 14714
rect 10236 14662 10258 14714
rect 10258 14662 10270 14714
rect 10270 14662 10292 14714
rect 10316 14662 10322 14714
rect 10322 14662 10334 14714
rect 10334 14662 10372 14714
rect 10396 14662 10398 14714
rect 10398 14662 10450 14714
rect 10450 14662 10452 14714
rect 10476 14662 10514 14714
rect 10514 14662 10526 14714
rect 10526 14662 10532 14714
rect 10556 14662 10578 14714
rect 10578 14662 10590 14714
rect 10590 14662 10612 14714
rect 10636 14662 10642 14714
rect 10642 14662 10654 14714
rect 10654 14662 10692 14714
rect 9516 14660 9572 14662
rect 9596 14660 9652 14662
rect 9676 14660 9732 14662
rect 9756 14660 9812 14662
rect 9836 14660 9892 14662
rect 9916 14660 9972 14662
rect 9996 14660 10052 14662
rect 10076 14660 10132 14662
rect 10156 14660 10212 14662
rect 10236 14660 10292 14662
rect 10316 14660 10372 14662
rect 10396 14660 10452 14662
rect 10476 14660 10532 14662
rect 10556 14660 10612 14662
rect 10636 14660 10692 14662
rect 10322 14048 10378 14104
rect 9516 13626 9572 13628
rect 9596 13626 9652 13628
rect 9676 13626 9732 13628
rect 9756 13626 9812 13628
rect 9836 13626 9892 13628
rect 9916 13626 9972 13628
rect 9996 13626 10052 13628
rect 10076 13626 10132 13628
rect 10156 13626 10212 13628
rect 10236 13626 10292 13628
rect 10316 13626 10372 13628
rect 10396 13626 10452 13628
rect 10476 13626 10532 13628
rect 10556 13626 10612 13628
rect 10636 13626 10692 13628
rect 9516 13574 9554 13626
rect 9554 13574 9566 13626
rect 9566 13574 9572 13626
rect 9596 13574 9618 13626
rect 9618 13574 9630 13626
rect 9630 13574 9652 13626
rect 9676 13574 9682 13626
rect 9682 13574 9694 13626
rect 9694 13574 9732 13626
rect 9756 13574 9758 13626
rect 9758 13574 9810 13626
rect 9810 13574 9812 13626
rect 9836 13574 9874 13626
rect 9874 13574 9886 13626
rect 9886 13574 9892 13626
rect 9916 13574 9938 13626
rect 9938 13574 9950 13626
rect 9950 13574 9972 13626
rect 9996 13574 10002 13626
rect 10002 13574 10014 13626
rect 10014 13574 10052 13626
rect 10076 13574 10078 13626
rect 10078 13574 10130 13626
rect 10130 13574 10132 13626
rect 10156 13574 10194 13626
rect 10194 13574 10206 13626
rect 10206 13574 10212 13626
rect 10236 13574 10258 13626
rect 10258 13574 10270 13626
rect 10270 13574 10292 13626
rect 10316 13574 10322 13626
rect 10322 13574 10334 13626
rect 10334 13574 10372 13626
rect 10396 13574 10398 13626
rect 10398 13574 10450 13626
rect 10450 13574 10452 13626
rect 10476 13574 10514 13626
rect 10514 13574 10526 13626
rect 10526 13574 10532 13626
rect 10556 13574 10578 13626
rect 10578 13574 10590 13626
rect 10590 13574 10612 13626
rect 10636 13574 10642 13626
rect 10642 13574 10654 13626
rect 10654 13574 10692 13626
rect 9516 13572 9572 13574
rect 9596 13572 9652 13574
rect 9676 13572 9732 13574
rect 9756 13572 9812 13574
rect 9836 13572 9892 13574
rect 9916 13572 9972 13574
rect 9996 13572 10052 13574
rect 10076 13572 10132 13574
rect 10156 13572 10212 13574
rect 10236 13572 10292 13574
rect 10316 13572 10372 13574
rect 10396 13572 10452 13574
rect 10476 13572 10532 13574
rect 10556 13572 10612 13574
rect 10636 13572 10692 13574
rect 9402 12688 9458 12744
rect 10138 12688 10194 12744
rect 10782 13232 10838 13288
rect 10874 12824 10930 12880
rect 9516 12538 9572 12540
rect 9596 12538 9652 12540
rect 9676 12538 9732 12540
rect 9756 12538 9812 12540
rect 9836 12538 9892 12540
rect 9916 12538 9972 12540
rect 9996 12538 10052 12540
rect 10076 12538 10132 12540
rect 10156 12538 10212 12540
rect 10236 12538 10292 12540
rect 10316 12538 10372 12540
rect 10396 12538 10452 12540
rect 10476 12538 10532 12540
rect 10556 12538 10612 12540
rect 10636 12538 10692 12540
rect 9516 12486 9554 12538
rect 9554 12486 9566 12538
rect 9566 12486 9572 12538
rect 9596 12486 9618 12538
rect 9618 12486 9630 12538
rect 9630 12486 9652 12538
rect 9676 12486 9682 12538
rect 9682 12486 9694 12538
rect 9694 12486 9732 12538
rect 9756 12486 9758 12538
rect 9758 12486 9810 12538
rect 9810 12486 9812 12538
rect 9836 12486 9874 12538
rect 9874 12486 9886 12538
rect 9886 12486 9892 12538
rect 9916 12486 9938 12538
rect 9938 12486 9950 12538
rect 9950 12486 9972 12538
rect 9996 12486 10002 12538
rect 10002 12486 10014 12538
rect 10014 12486 10052 12538
rect 10076 12486 10078 12538
rect 10078 12486 10130 12538
rect 10130 12486 10132 12538
rect 10156 12486 10194 12538
rect 10194 12486 10206 12538
rect 10206 12486 10212 12538
rect 10236 12486 10258 12538
rect 10258 12486 10270 12538
rect 10270 12486 10292 12538
rect 10316 12486 10322 12538
rect 10322 12486 10334 12538
rect 10334 12486 10372 12538
rect 10396 12486 10398 12538
rect 10398 12486 10450 12538
rect 10450 12486 10452 12538
rect 10476 12486 10514 12538
rect 10514 12486 10526 12538
rect 10526 12486 10532 12538
rect 10556 12486 10578 12538
rect 10578 12486 10590 12538
rect 10590 12486 10612 12538
rect 10636 12486 10642 12538
rect 10642 12486 10654 12538
rect 10654 12486 10692 12538
rect 9516 12484 9572 12486
rect 9596 12484 9652 12486
rect 9676 12484 9732 12486
rect 9756 12484 9812 12486
rect 9836 12484 9892 12486
rect 9916 12484 9972 12486
rect 9996 12484 10052 12486
rect 10076 12484 10132 12486
rect 10156 12484 10212 12486
rect 10236 12484 10292 12486
rect 10316 12484 10372 12486
rect 10396 12484 10452 12486
rect 10476 12484 10532 12486
rect 10556 12484 10612 12486
rect 10636 12484 10692 12486
rect 9402 12300 9458 12336
rect 9402 12280 9404 12300
rect 9404 12280 9456 12300
rect 9456 12280 9458 12300
rect 9310 11872 9366 11928
rect 9218 11736 9274 11792
rect 9402 11756 9458 11792
rect 9402 11736 9404 11756
rect 9404 11736 9456 11756
rect 9456 11736 9458 11756
rect 8574 10512 8630 10568
rect 8942 11464 8998 11520
rect 9034 11328 9090 11384
rect 8850 10920 8906 10976
rect 8850 7792 8906 7848
rect 9034 10240 9090 10296
rect 9770 12144 9826 12200
rect 10322 12280 10378 12336
rect 9862 11736 9918 11792
rect 10690 12280 10746 12336
rect 10046 11600 10102 11656
rect 10230 11600 10286 11656
rect 10782 12144 10838 12200
rect 17516 16890 17572 16892
rect 17596 16890 17652 16892
rect 17676 16890 17732 16892
rect 17756 16890 17812 16892
rect 17836 16890 17892 16892
rect 17916 16890 17972 16892
rect 17996 16890 18052 16892
rect 18076 16890 18132 16892
rect 18156 16890 18212 16892
rect 18236 16890 18292 16892
rect 18316 16890 18372 16892
rect 18396 16890 18452 16892
rect 18476 16890 18532 16892
rect 18556 16890 18612 16892
rect 18636 16890 18692 16892
rect 17516 16838 17554 16890
rect 17554 16838 17566 16890
rect 17566 16838 17572 16890
rect 17596 16838 17618 16890
rect 17618 16838 17630 16890
rect 17630 16838 17652 16890
rect 17676 16838 17682 16890
rect 17682 16838 17694 16890
rect 17694 16838 17732 16890
rect 17756 16838 17758 16890
rect 17758 16838 17810 16890
rect 17810 16838 17812 16890
rect 17836 16838 17874 16890
rect 17874 16838 17886 16890
rect 17886 16838 17892 16890
rect 17916 16838 17938 16890
rect 17938 16838 17950 16890
rect 17950 16838 17972 16890
rect 17996 16838 18002 16890
rect 18002 16838 18014 16890
rect 18014 16838 18052 16890
rect 18076 16838 18078 16890
rect 18078 16838 18130 16890
rect 18130 16838 18132 16890
rect 18156 16838 18194 16890
rect 18194 16838 18206 16890
rect 18206 16838 18212 16890
rect 18236 16838 18258 16890
rect 18258 16838 18270 16890
rect 18270 16838 18292 16890
rect 18316 16838 18322 16890
rect 18322 16838 18334 16890
rect 18334 16838 18372 16890
rect 18396 16838 18398 16890
rect 18398 16838 18450 16890
rect 18450 16838 18452 16890
rect 18476 16838 18514 16890
rect 18514 16838 18526 16890
rect 18526 16838 18532 16890
rect 18556 16838 18578 16890
rect 18578 16838 18590 16890
rect 18590 16838 18612 16890
rect 18636 16838 18642 16890
rect 18642 16838 18654 16890
rect 18654 16838 18692 16890
rect 17516 16836 17572 16838
rect 17596 16836 17652 16838
rect 17676 16836 17732 16838
rect 17756 16836 17812 16838
rect 17836 16836 17892 16838
rect 17916 16836 17972 16838
rect 17996 16836 18052 16838
rect 18076 16836 18132 16838
rect 18156 16836 18212 16838
rect 18236 16836 18292 16838
rect 18316 16836 18372 16838
rect 18396 16836 18452 16838
rect 18476 16836 18532 16838
rect 18556 16836 18612 16838
rect 18636 16836 18692 16838
rect 18786 16632 18842 16688
rect 11426 15544 11482 15600
rect 11150 12552 11206 12608
rect 11518 15272 11574 15328
rect 10782 11772 10784 11792
rect 10784 11772 10836 11792
rect 10836 11772 10838 11792
rect 10782 11736 10838 11772
rect 9516 11450 9572 11452
rect 9596 11450 9652 11452
rect 9676 11450 9732 11452
rect 9756 11450 9812 11452
rect 9836 11450 9892 11452
rect 9916 11450 9972 11452
rect 9996 11450 10052 11452
rect 10076 11450 10132 11452
rect 10156 11450 10212 11452
rect 10236 11450 10292 11452
rect 10316 11450 10372 11452
rect 10396 11450 10452 11452
rect 10476 11450 10532 11452
rect 10556 11450 10612 11452
rect 10636 11450 10692 11452
rect 9516 11398 9554 11450
rect 9554 11398 9566 11450
rect 9566 11398 9572 11450
rect 9596 11398 9618 11450
rect 9618 11398 9630 11450
rect 9630 11398 9652 11450
rect 9676 11398 9682 11450
rect 9682 11398 9694 11450
rect 9694 11398 9732 11450
rect 9756 11398 9758 11450
rect 9758 11398 9810 11450
rect 9810 11398 9812 11450
rect 9836 11398 9874 11450
rect 9874 11398 9886 11450
rect 9886 11398 9892 11450
rect 9916 11398 9938 11450
rect 9938 11398 9950 11450
rect 9950 11398 9972 11450
rect 9996 11398 10002 11450
rect 10002 11398 10014 11450
rect 10014 11398 10052 11450
rect 10076 11398 10078 11450
rect 10078 11398 10130 11450
rect 10130 11398 10132 11450
rect 10156 11398 10194 11450
rect 10194 11398 10206 11450
rect 10206 11398 10212 11450
rect 10236 11398 10258 11450
rect 10258 11398 10270 11450
rect 10270 11398 10292 11450
rect 10316 11398 10322 11450
rect 10322 11398 10334 11450
rect 10334 11398 10372 11450
rect 10396 11398 10398 11450
rect 10398 11398 10450 11450
rect 10450 11398 10452 11450
rect 10476 11398 10514 11450
rect 10514 11398 10526 11450
rect 10526 11398 10532 11450
rect 10556 11398 10578 11450
rect 10578 11398 10590 11450
rect 10590 11398 10612 11450
rect 10636 11398 10642 11450
rect 10642 11398 10654 11450
rect 10654 11398 10692 11450
rect 9516 11396 9572 11398
rect 9596 11396 9652 11398
rect 9676 11396 9732 11398
rect 9756 11396 9812 11398
rect 9836 11396 9892 11398
rect 9916 11396 9972 11398
rect 9996 11396 10052 11398
rect 10076 11396 10132 11398
rect 10156 11396 10212 11398
rect 10236 11396 10292 11398
rect 10316 11396 10372 11398
rect 10396 11396 10452 11398
rect 10476 11396 10532 11398
rect 10556 11396 10612 11398
rect 10636 11396 10692 11398
rect 9954 11212 10010 11248
rect 9954 11192 9956 11212
rect 9956 11192 10008 11212
rect 10008 11192 10010 11212
rect 10598 11192 10654 11248
rect 9678 11056 9734 11112
rect 9402 10512 9458 10568
rect 9586 10512 9642 10568
rect 9862 10920 9918 10976
rect 10138 10512 10194 10568
rect 11058 12008 11114 12064
rect 10966 10920 11022 10976
rect 10690 10512 10746 10568
rect 10782 10376 10838 10432
rect 9516 10362 9572 10364
rect 9596 10362 9652 10364
rect 9676 10362 9732 10364
rect 9756 10362 9812 10364
rect 9836 10362 9892 10364
rect 9916 10362 9972 10364
rect 9996 10362 10052 10364
rect 10076 10362 10132 10364
rect 10156 10362 10212 10364
rect 10236 10362 10292 10364
rect 10316 10362 10372 10364
rect 10396 10362 10452 10364
rect 10476 10362 10532 10364
rect 10556 10362 10612 10364
rect 10636 10362 10692 10364
rect 9516 10310 9554 10362
rect 9554 10310 9566 10362
rect 9566 10310 9572 10362
rect 9596 10310 9618 10362
rect 9618 10310 9630 10362
rect 9630 10310 9652 10362
rect 9676 10310 9682 10362
rect 9682 10310 9694 10362
rect 9694 10310 9732 10362
rect 9756 10310 9758 10362
rect 9758 10310 9810 10362
rect 9810 10310 9812 10362
rect 9836 10310 9874 10362
rect 9874 10310 9886 10362
rect 9886 10310 9892 10362
rect 9916 10310 9938 10362
rect 9938 10310 9950 10362
rect 9950 10310 9972 10362
rect 9996 10310 10002 10362
rect 10002 10310 10014 10362
rect 10014 10310 10052 10362
rect 10076 10310 10078 10362
rect 10078 10310 10130 10362
rect 10130 10310 10132 10362
rect 10156 10310 10194 10362
rect 10194 10310 10206 10362
rect 10206 10310 10212 10362
rect 10236 10310 10258 10362
rect 10258 10310 10270 10362
rect 10270 10310 10292 10362
rect 10316 10310 10322 10362
rect 10322 10310 10334 10362
rect 10334 10310 10372 10362
rect 10396 10310 10398 10362
rect 10398 10310 10450 10362
rect 10450 10310 10452 10362
rect 10476 10310 10514 10362
rect 10514 10310 10526 10362
rect 10526 10310 10532 10362
rect 10556 10310 10578 10362
rect 10578 10310 10590 10362
rect 10590 10310 10612 10362
rect 10636 10310 10642 10362
rect 10642 10310 10654 10362
rect 10654 10310 10692 10362
rect 9516 10308 9572 10310
rect 9596 10308 9652 10310
rect 9676 10308 9732 10310
rect 9756 10308 9812 10310
rect 9836 10308 9892 10310
rect 9916 10308 9972 10310
rect 9996 10308 10052 10310
rect 10076 10308 10132 10310
rect 10156 10308 10212 10310
rect 10236 10308 10292 10310
rect 10316 10308 10372 10310
rect 10396 10308 10452 10310
rect 10476 10308 10532 10310
rect 10556 10308 10612 10310
rect 10636 10308 10692 10310
rect 9402 10104 9458 10160
rect 9770 10104 9826 10160
rect 10690 9444 10746 9480
rect 10690 9424 10692 9444
rect 10692 9424 10744 9444
rect 10744 9424 10746 9444
rect 9516 9274 9572 9276
rect 9596 9274 9652 9276
rect 9676 9274 9732 9276
rect 9756 9274 9812 9276
rect 9836 9274 9892 9276
rect 9916 9274 9972 9276
rect 9996 9274 10052 9276
rect 10076 9274 10132 9276
rect 10156 9274 10212 9276
rect 10236 9274 10292 9276
rect 10316 9274 10372 9276
rect 10396 9274 10452 9276
rect 10476 9274 10532 9276
rect 10556 9274 10612 9276
rect 10636 9274 10692 9276
rect 9516 9222 9554 9274
rect 9554 9222 9566 9274
rect 9566 9222 9572 9274
rect 9596 9222 9618 9274
rect 9618 9222 9630 9274
rect 9630 9222 9652 9274
rect 9676 9222 9682 9274
rect 9682 9222 9694 9274
rect 9694 9222 9732 9274
rect 9756 9222 9758 9274
rect 9758 9222 9810 9274
rect 9810 9222 9812 9274
rect 9836 9222 9874 9274
rect 9874 9222 9886 9274
rect 9886 9222 9892 9274
rect 9916 9222 9938 9274
rect 9938 9222 9950 9274
rect 9950 9222 9972 9274
rect 9996 9222 10002 9274
rect 10002 9222 10014 9274
rect 10014 9222 10052 9274
rect 10076 9222 10078 9274
rect 10078 9222 10130 9274
rect 10130 9222 10132 9274
rect 10156 9222 10194 9274
rect 10194 9222 10206 9274
rect 10206 9222 10212 9274
rect 10236 9222 10258 9274
rect 10258 9222 10270 9274
rect 10270 9222 10292 9274
rect 10316 9222 10322 9274
rect 10322 9222 10334 9274
rect 10334 9222 10372 9274
rect 10396 9222 10398 9274
rect 10398 9222 10450 9274
rect 10450 9222 10452 9274
rect 10476 9222 10514 9274
rect 10514 9222 10526 9274
rect 10526 9222 10532 9274
rect 10556 9222 10578 9274
rect 10578 9222 10590 9274
rect 10590 9222 10612 9274
rect 10636 9222 10642 9274
rect 10642 9222 10654 9274
rect 10654 9222 10692 9274
rect 9516 9220 9572 9222
rect 9596 9220 9652 9222
rect 9676 9220 9732 9222
rect 9756 9220 9812 9222
rect 9836 9220 9892 9222
rect 9916 9220 9972 9222
rect 9996 9220 10052 9222
rect 10076 9220 10132 9222
rect 10156 9220 10212 9222
rect 10236 9220 10292 9222
rect 10316 9220 10372 9222
rect 10396 9220 10452 9222
rect 10476 9220 10532 9222
rect 10556 9220 10612 9222
rect 10636 9220 10692 9222
rect 9126 3576 9182 3632
rect 8942 3440 8998 3496
rect 9516 8186 9572 8188
rect 9596 8186 9652 8188
rect 9676 8186 9732 8188
rect 9756 8186 9812 8188
rect 9836 8186 9892 8188
rect 9916 8186 9972 8188
rect 9996 8186 10052 8188
rect 10076 8186 10132 8188
rect 10156 8186 10212 8188
rect 10236 8186 10292 8188
rect 10316 8186 10372 8188
rect 10396 8186 10452 8188
rect 10476 8186 10532 8188
rect 10556 8186 10612 8188
rect 10636 8186 10692 8188
rect 9516 8134 9554 8186
rect 9554 8134 9566 8186
rect 9566 8134 9572 8186
rect 9596 8134 9618 8186
rect 9618 8134 9630 8186
rect 9630 8134 9652 8186
rect 9676 8134 9682 8186
rect 9682 8134 9694 8186
rect 9694 8134 9732 8186
rect 9756 8134 9758 8186
rect 9758 8134 9810 8186
rect 9810 8134 9812 8186
rect 9836 8134 9874 8186
rect 9874 8134 9886 8186
rect 9886 8134 9892 8186
rect 9916 8134 9938 8186
rect 9938 8134 9950 8186
rect 9950 8134 9972 8186
rect 9996 8134 10002 8186
rect 10002 8134 10014 8186
rect 10014 8134 10052 8186
rect 10076 8134 10078 8186
rect 10078 8134 10130 8186
rect 10130 8134 10132 8186
rect 10156 8134 10194 8186
rect 10194 8134 10206 8186
rect 10206 8134 10212 8186
rect 10236 8134 10258 8186
rect 10258 8134 10270 8186
rect 10270 8134 10292 8186
rect 10316 8134 10322 8186
rect 10322 8134 10334 8186
rect 10334 8134 10372 8186
rect 10396 8134 10398 8186
rect 10398 8134 10450 8186
rect 10450 8134 10452 8186
rect 10476 8134 10514 8186
rect 10514 8134 10526 8186
rect 10526 8134 10532 8186
rect 10556 8134 10578 8186
rect 10578 8134 10590 8186
rect 10590 8134 10612 8186
rect 10636 8134 10642 8186
rect 10642 8134 10654 8186
rect 10654 8134 10692 8186
rect 9516 8132 9572 8134
rect 9596 8132 9652 8134
rect 9676 8132 9732 8134
rect 9756 8132 9812 8134
rect 9836 8132 9892 8134
rect 9916 8132 9972 8134
rect 9996 8132 10052 8134
rect 10076 8132 10132 8134
rect 10156 8132 10212 8134
rect 10236 8132 10292 8134
rect 10316 8132 10372 8134
rect 10396 8132 10452 8134
rect 10476 8132 10532 8134
rect 10556 8132 10612 8134
rect 10636 8132 10692 8134
rect 9516 7098 9572 7100
rect 9596 7098 9652 7100
rect 9676 7098 9732 7100
rect 9756 7098 9812 7100
rect 9836 7098 9892 7100
rect 9916 7098 9972 7100
rect 9996 7098 10052 7100
rect 10076 7098 10132 7100
rect 10156 7098 10212 7100
rect 10236 7098 10292 7100
rect 10316 7098 10372 7100
rect 10396 7098 10452 7100
rect 10476 7098 10532 7100
rect 10556 7098 10612 7100
rect 10636 7098 10692 7100
rect 9516 7046 9554 7098
rect 9554 7046 9566 7098
rect 9566 7046 9572 7098
rect 9596 7046 9618 7098
rect 9618 7046 9630 7098
rect 9630 7046 9652 7098
rect 9676 7046 9682 7098
rect 9682 7046 9694 7098
rect 9694 7046 9732 7098
rect 9756 7046 9758 7098
rect 9758 7046 9810 7098
rect 9810 7046 9812 7098
rect 9836 7046 9874 7098
rect 9874 7046 9886 7098
rect 9886 7046 9892 7098
rect 9916 7046 9938 7098
rect 9938 7046 9950 7098
rect 9950 7046 9972 7098
rect 9996 7046 10002 7098
rect 10002 7046 10014 7098
rect 10014 7046 10052 7098
rect 10076 7046 10078 7098
rect 10078 7046 10130 7098
rect 10130 7046 10132 7098
rect 10156 7046 10194 7098
rect 10194 7046 10206 7098
rect 10206 7046 10212 7098
rect 10236 7046 10258 7098
rect 10258 7046 10270 7098
rect 10270 7046 10292 7098
rect 10316 7046 10322 7098
rect 10322 7046 10334 7098
rect 10334 7046 10372 7098
rect 10396 7046 10398 7098
rect 10398 7046 10450 7098
rect 10450 7046 10452 7098
rect 10476 7046 10514 7098
rect 10514 7046 10526 7098
rect 10526 7046 10532 7098
rect 10556 7046 10578 7098
rect 10578 7046 10590 7098
rect 10590 7046 10612 7098
rect 10636 7046 10642 7098
rect 10642 7046 10654 7098
rect 10654 7046 10692 7098
rect 9516 7044 9572 7046
rect 9596 7044 9652 7046
rect 9676 7044 9732 7046
rect 9756 7044 9812 7046
rect 9836 7044 9892 7046
rect 9916 7044 9972 7046
rect 9996 7044 10052 7046
rect 10076 7044 10132 7046
rect 10156 7044 10212 7046
rect 10236 7044 10292 7046
rect 10316 7044 10372 7046
rect 10396 7044 10452 7046
rect 10476 7044 10532 7046
rect 10556 7044 10612 7046
rect 10636 7044 10692 7046
rect 9516 6010 9572 6012
rect 9596 6010 9652 6012
rect 9676 6010 9732 6012
rect 9756 6010 9812 6012
rect 9836 6010 9892 6012
rect 9916 6010 9972 6012
rect 9996 6010 10052 6012
rect 10076 6010 10132 6012
rect 10156 6010 10212 6012
rect 10236 6010 10292 6012
rect 10316 6010 10372 6012
rect 10396 6010 10452 6012
rect 10476 6010 10532 6012
rect 10556 6010 10612 6012
rect 10636 6010 10692 6012
rect 9516 5958 9554 6010
rect 9554 5958 9566 6010
rect 9566 5958 9572 6010
rect 9596 5958 9618 6010
rect 9618 5958 9630 6010
rect 9630 5958 9652 6010
rect 9676 5958 9682 6010
rect 9682 5958 9694 6010
rect 9694 5958 9732 6010
rect 9756 5958 9758 6010
rect 9758 5958 9810 6010
rect 9810 5958 9812 6010
rect 9836 5958 9874 6010
rect 9874 5958 9886 6010
rect 9886 5958 9892 6010
rect 9916 5958 9938 6010
rect 9938 5958 9950 6010
rect 9950 5958 9972 6010
rect 9996 5958 10002 6010
rect 10002 5958 10014 6010
rect 10014 5958 10052 6010
rect 10076 5958 10078 6010
rect 10078 5958 10130 6010
rect 10130 5958 10132 6010
rect 10156 5958 10194 6010
rect 10194 5958 10206 6010
rect 10206 5958 10212 6010
rect 10236 5958 10258 6010
rect 10258 5958 10270 6010
rect 10270 5958 10292 6010
rect 10316 5958 10322 6010
rect 10322 5958 10334 6010
rect 10334 5958 10372 6010
rect 10396 5958 10398 6010
rect 10398 5958 10450 6010
rect 10450 5958 10452 6010
rect 10476 5958 10514 6010
rect 10514 5958 10526 6010
rect 10526 5958 10532 6010
rect 10556 5958 10578 6010
rect 10578 5958 10590 6010
rect 10590 5958 10612 6010
rect 10636 5958 10642 6010
rect 10642 5958 10654 6010
rect 10654 5958 10692 6010
rect 9516 5956 9572 5958
rect 9596 5956 9652 5958
rect 9676 5956 9732 5958
rect 9756 5956 9812 5958
rect 9836 5956 9892 5958
rect 9916 5956 9972 5958
rect 9996 5956 10052 5958
rect 10076 5956 10132 5958
rect 10156 5956 10212 5958
rect 10236 5956 10292 5958
rect 10316 5956 10372 5958
rect 10396 5956 10452 5958
rect 10476 5956 10532 5958
rect 10556 5956 10612 5958
rect 10636 5956 10692 5958
rect 9516 4922 9572 4924
rect 9596 4922 9652 4924
rect 9676 4922 9732 4924
rect 9756 4922 9812 4924
rect 9836 4922 9892 4924
rect 9916 4922 9972 4924
rect 9996 4922 10052 4924
rect 10076 4922 10132 4924
rect 10156 4922 10212 4924
rect 10236 4922 10292 4924
rect 10316 4922 10372 4924
rect 10396 4922 10452 4924
rect 10476 4922 10532 4924
rect 10556 4922 10612 4924
rect 10636 4922 10692 4924
rect 9516 4870 9554 4922
rect 9554 4870 9566 4922
rect 9566 4870 9572 4922
rect 9596 4870 9618 4922
rect 9618 4870 9630 4922
rect 9630 4870 9652 4922
rect 9676 4870 9682 4922
rect 9682 4870 9694 4922
rect 9694 4870 9732 4922
rect 9756 4870 9758 4922
rect 9758 4870 9810 4922
rect 9810 4870 9812 4922
rect 9836 4870 9874 4922
rect 9874 4870 9886 4922
rect 9886 4870 9892 4922
rect 9916 4870 9938 4922
rect 9938 4870 9950 4922
rect 9950 4870 9972 4922
rect 9996 4870 10002 4922
rect 10002 4870 10014 4922
rect 10014 4870 10052 4922
rect 10076 4870 10078 4922
rect 10078 4870 10130 4922
rect 10130 4870 10132 4922
rect 10156 4870 10194 4922
rect 10194 4870 10206 4922
rect 10206 4870 10212 4922
rect 10236 4870 10258 4922
rect 10258 4870 10270 4922
rect 10270 4870 10292 4922
rect 10316 4870 10322 4922
rect 10322 4870 10334 4922
rect 10334 4870 10372 4922
rect 10396 4870 10398 4922
rect 10398 4870 10450 4922
rect 10450 4870 10452 4922
rect 10476 4870 10514 4922
rect 10514 4870 10526 4922
rect 10526 4870 10532 4922
rect 10556 4870 10578 4922
rect 10578 4870 10590 4922
rect 10590 4870 10612 4922
rect 10636 4870 10642 4922
rect 10642 4870 10654 4922
rect 10654 4870 10692 4922
rect 9516 4868 9572 4870
rect 9596 4868 9652 4870
rect 9676 4868 9732 4870
rect 9756 4868 9812 4870
rect 9836 4868 9892 4870
rect 9916 4868 9972 4870
rect 9996 4868 10052 4870
rect 10076 4868 10132 4870
rect 10156 4868 10212 4870
rect 10236 4868 10292 4870
rect 10316 4868 10372 4870
rect 10396 4868 10452 4870
rect 10476 4868 10532 4870
rect 10556 4868 10612 4870
rect 10636 4868 10692 4870
rect 10690 4548 10746 4584
rect 10690 4528 10692 4548
rect 10692 4528 10744 4548
rect 10744 4528 10746 4548
rect 9516 3834 9572 3836
rect 9596 3834 9652 3836
rect 9676 3834 9732 3836
rect 9756 3834 9812 3836
rect 9836 3834 9892 3836
rect 9916 3834 9972 3836
rect 9996 3834 10052 3836
rect 10076 3834 10132 3836
rect 10156 3834 10212 3836
rect 10236 3834 10292 3836
rect 10316 3834 10372 3836
rect 10396 3834 10452 3836
rect 10476 3834 10532 3836
rect 10556 3834 10612 3836
rect 10636 3834 10692 3836
rect 9516 3782 9554 3834
rect 9554 3782 9566 3834
rect 9566 3782 9572 3834
rect 9596 3782 9618 3834
rect 9618 3782 9630 3834
rect 9630 3782 9652 3834
rect 9676 3782 9682 3834
rect 9682 3782 9694 3834
rect 9694 3782 9732 3834
rect 9756 3782 9758 3834
rect 9758 3782 9810 3834
rect 9810 3782 9812 3834
rect 9836 3782 9874 3834
rect 9874 3782 9886 3834
rect 9886 3782 9892 3834
rect 9916 3782 9938 3834
rect 9938 3782 9950 3834
rect 9950 3782 9972 3834
rect 9996 3782 10002 3834
rect 10002 3782 10014 3834
rect 10014 3782 10052 3834
rect 10076 3782 10078 3834
rect 10078 3782 10130 3834
rect 10130 3782 10132 3834
rect 10156 3782 10194 3834
rect 10194 3782 10206 3834
rect 10206 3782 10212 3834
rect 10236 3782 10258 3834
rect 10258 3782 10270 3834
rect 10270 3782 10292 3834
rect 10316 3782 10322 3834
rect 10322 3782 10334 3834
rect 10334 3782 10372 3834
rect 10396 3782 10398 3834
rect 10398 3782 10450 3834
rect 10450 3782 10452 3834
rect 10476 3782 10514 3834
rect 10514 3782 10526 3834
rect 10526 3782 10532 3834
rect 10556 3782 10578 3834
rect 10578 3782 10590 3834
rect 10590 3782 10612 3834
rect 10636 3782 10642 3834
rect 10642 3782 10654 3834
rect 10654 3782 10692 3834
rect 9516 3780 9572 3782
rect 9596 3780 9652 3782
rect 9676 3780 9732 3782
rect 9756 3780 9812 3782
rect 9836 3780 9892 3782
rect 9916 3780 9972 3782
rect 9996 3780 10052 3782
rect 10076 3780 10132 3782
rect 10156 3780 10212 3782
rect 10236 3780 10292 3782
rect 10316 3780 10372 3782
rect 10396 3780 10452 3782
rect 10476 3780 10532 3782
rect 10556 3780 10612 3782
rect 10636 3780 10692 3782
rect 9586 3576 9642 3632
rect 10414 3304 10470 3360
rect 10598 3168 10654 3224
rect 11058 9152 11114 9208
rect 11058 9016 11114 9072
rect 9516 2746 9572 2748
rect 9596 2746 9652 2748
rect 9676 2746 9732 2748
rect 9756 2746 9812 2748
rect 9836 2746 9892 2748
rect 9916 2746 9972 2748
rect 9996 2746 10052 2748
rect 10076 2746 10132 2748
rect 10156 2746 10212 2748
rect 10236 2746 10292 2748
rect 10316 2746 10372 2748
rect 10396 2746 10452 2748
rect 10476 2746 10532 2748
rect 10556 2746 10612 2748
rect 10636 2746 10692 2748
rect 9516 2694 9554 2746
rect 9554 2694 9566 2746
rect 9566 2694 9572 2746
rect 9596 2694 9618 2746
rect 9618 2694 9630 2746
rect 9630 2694 9652 2746
rect 9676 2694 9682 2746
rect 9682 2694 9694 2746
rect 9694 2694 9732 2746
rect 9756 2694 9758 2746
rect 9758 2694 9810 2746
rect 9810 2694 9812 2746
rect 9836 2694 9874 2746
rect 9874 2694 9886 2746
rect 9886 2694 9892 2746
rect 9916 2694 9938 2746
rect 9938 2694 9950 2746
rect 9950 2694 9972 2746
rect 9996 2694 10002 2746
rect 10002 2694 10014 2746
rect 10014 2694 10052 2746
rect 10076 2694 10078 2746
rect 10078 2694 10130 2746
rect 10130 2694 10132 2746
rect 10156 2694 10194 2746
rect 10194 2694 10206 2746
rect 10206 2694 10212 2746
rect 10236 2694 10258 2746
rect 10258 2694 10270 2746
rect 10270 2694 10292 2746
rect 10316 2694 10322 2746
rect 10322 2694 10334 2746
rect 10334 2694 10372 2746
rect 10396 2694 10398 2746
rect 10398 2694 10450 2746
rect 10450 2694 10452 2746
rect 10476 2694 10514 2746
rect 10514 2694 10526 2746
rect 10526 2694 10532 2746
rect 10556 2694 10578 2746
rect 10578 2694 10590 2746
rect 10590 2694 10612 2746
rect 10636 2694 10642 2746
rect 10642 2694 10654 2746
rect 10654 2694 10692 2746
rect 9516 2692 9572 2694
rect 9596 2692 9652 2694
rect 9676 2692 9732 2694
rect 9756 2692 9812 2694
rect 9836 2692 9892 2694
rect 9916 2692 9972 2694
rect 9996 2692 10052 2694
rect 10076 2692 10132 2694
rect 10156 2692 10212 2694
rect 10236 2692 10292 2694
rect 10316 2692 10372 2694
rect 10396 2692 10452 2694
rect 10476 2692 10532 2694
rect 10556 2692 10612 2694
rect 10636 2692 10692 2694
rect 10874 2760 10930 2816
rect 11702 14864 11758 14920
rect 11794 12960 11850 13016
rect 11794 12552 11850 12608
rect 11702 11736 11758 11792
rect 11794 11294 11850 11350
rect 11702 11056 11758 11112
rect 11426 10920 11482 10976
rect 11242 9832 11298 9888
rect 11334 9560 11390 9616
rect 11242 7656 11298 7712
rect 11058 6840 11114 6896
rect 11058 3984 11114 4040
rect 11058 3576 11114 3632
rect 11058 3304 11114 3360
rect 11426 7656 11482 7712
rect 12070 11192 12126 11248
rect 11978 11056 12034 11112
rect 11794 10648 11850 10704
rect 11794 10512 11850 10568
rect 11702 10104 11758 10160
rect 11702 6976 11758 7032
rect 11242 3848 11298 3904
rect 13516 16346 13572 16348
rect 13596 16346 13652 16348
rect 13676 16346 13732 16348
rect 13756 16346 13812 16348
rect 13836 16346 13892 16348
rect 13916 16346 13972 16348
rect 13996 16346 14052 16348
rect 14076 16346 14132 16348
rect 14156 16346 14212 16348
rect 14236 16346 14292 16348
rect 14316 16346 14372 16348
rect 14396 16346 14452 16348
rect 14476 16346 14532 16348
rect 14556 16346 14612 16348
rect 14636 16346 14692 16348
rect 13516 16294 13554 16346
rect 13554 16294 13566 16346
rect 13566 16294 13572 16346
rect 13596 16294 13618 16346
rect 13618 16294 13630 16346
rect 13630 16294 13652 16346
rect 13676 16294 13682 16346
rect 13682 16294 13694 16346
rect 13694 16294 13732 16346
rect 13756 16294 13758 16346
rect 13758 16294 13810 16346
rect 13810 16294 13812 16346
rect 13836 16294 13874 16346
rect 13874 16294 13886 16346
rect 13886 16294 13892 16346
rect 13916 16294 13938 16346
rect 13938 16294 13950 16346
rect 13950 16294 13972 16346
rect 13996 16294 14002 16346
rect 14002 16294 14014 16346
rect 14014 16294 14052 16346
rect 14076 16294 14078 16346
rect 14078 16294 14130 16346
rect 14130 16294 14132 16346
rect 14156 16294 14194 16346
rect 14194 16294 14206 16346
rect 14206 16294 14212 16346
rect 14236 16294 14258 16346
rect 14258 16294 14270 16346
rect 14270 16294 14292 16346
rect 14316 16294 14322 16346
rect 14322 16294 14334 16346
rect 14334 16294 14372 16346
rect 14396 16294 14398 16346
rect 14398 16294 14450 16346
rect 14450 16294 14452 16346
rect 14476 16294 14514 16346
rect 14514 16294 14526 16346
rect 14526 16294 14532 16346
rect 14556 16294 14578 16346
rect 14578 16294 14590 16346
rect 14590 16294 14612 16346
rect 14636 16294 14642 16346
rect 14642 16294 14654 16346
rect 14654 16294 14692 16346
rect 13516 16292 13572 16294
rect 13596 16292 13652 16294
rect 13676 16292 13732 16294
rect 13756 16292 13812 16294
rect 13836 16292 13892 16294
rect 13916 16292 13972 16294
rect 13996 16292 14052 16294
rect 14076 16292 14132 16294
rect 14156 16292 14212 16294
rect 14236 16292 14292 16294
rect 14316 16292 14372 16294
rect 14396 16292 14452 16294
rect 14476 16292 14532 16294
rect 14556 16292 14612 16294
rect 14636 16292 14692 16294
rect 16578 15952 16634 16008
rect 12254 12552 12310 12608
rect 12346 12416 12402 12472
rect 12346 12144 12402 12200
rect 12254 12008 12310 12064
rect 12162 10104 12218 10160
rect 12346 11328 12402 11384
rect 12438 10512 12494 10568
rect 12438 10376 12494 10432
rect 13516 15258 13572 15260
rect 13596 15258 13652 15260
rect 13676 15258 13732 15260
rect 13756 15258 13812 15260
rect 13836 15258 13892 15260
rect 13916 15258 13972 15260
rect 13996 15258 14052 15260
rect 14076 15258 14132 15260
rect 14156 15258 14212 15260
rect 14236 15258 14292 15260
rect 14316 15258 14372 15260
rect 14396 15258 14452 15260
rect 14476 15258 14532 15260
rect 14556 15258 14612 15260
rect 14636 15258 14692 15260
rect 13516 15206 13554 15258
rect 13554 15206 13566 15258
rect 13566 15206 13572 15258
rect 13596 15206 13618 15258
rect 13618 15206 13630 15258
rect 13630 15206 13652 15258
rect 13676 15206 13682 15258
rect 13682 15206 13694 15258
rect 13694 15206 13732 15258
rect 13756 15206 13758 15258
rect 13758 15206 13810 15258
rect 13810 15206 13812 15258
rect 13836 15206 13874 15258
rect 13874 15206 13886 15258
rect 13886 15206 13892 15258
rect 13916 15206 13938 15258
rect 13938 15206 13950 15258
rect 13950 15206 13972 15258
rect 13996 15206 14002 15258
rect 14002 15206 14014 15258
rect 14014 15206 14052 15258
rect 14076 15206 14078 15258
rect 14078 15206 14130 15258
rect 14130 15206 14132 15258
rect 14156 15206 14194 15258
rect 14194 15206 14206 15258
rect 14206 15206 14212 15258
rect 14236 15206 14258 15258
rect 14258 15206 14270 15258
rect 14270 15206 14292 15258
rect 14316 15206 14322 15258
rect 14322 15206 14334 15258
rect 14334 15206 14372 15258
rect 14396 15206 14398 15258
rect 14398 15206 14450 15258
rect 14450 15206 14452 15258
rect 14476 15206 14514 15258
rect 14514 15206 14526 15258
rect 14526 15206 14532 15258
rect 14556 15206 14578 15258
rect 14578 15206 14590 15258
rect 14590 15206 14612 15258
rect 14636 15206 14642 15258
rect 14642 15206 14654 15258
rect 14654 15206 14692 15258
rect 13516 15204 13572 15206
rect 13596 15204 13652 15206
rect 13676 15204 13732 15206
rect 13756 15204 13812 15206
rect 13836 15204 13892 15206
rect 13916 15204 13972 15206
rect 13996 15204 14052 15206
rect 14076 15204 14132 15206
rect 14156 15204 14212 15206
rect 14236 15204 14292 15206
rect 14316 15204 14372 15206
rect 14396 15204 14452 15206
rect 14476 15204 14532 15206
rect 14556 15204 14612 15206
rect 14636 15204 14692 15206
rect 12806 11736 12862 11792
rect 12438 8064 12494 8120
rect 12714 8608 12770 8664
rect 12622 7112 12678 7168
rect 12438 6740 12440 6760
rect 12440 6740 12492 6760
rect 12492 6740 12494 6760
rect 12438 6704 12494 6740
rect 12530 6316 12586 6352
rect 12530 6296 12532 6316
rect 12532 6296 12584 6316
rect 12584 6296 12586 6316
rect 11702 2760 11758 2816
rect 12346 3848 12402 3904
rect 13516 14170 13572 14172
rect 13596 14170 13652 14172
rect 13676 14170 13732 14172
rect 13756 14170 13812 14172
rect 13836 14170 13892 14172
rect 13916 14170 13972 14172
rect 13996 14170 14052 14172
rect 14076 14170 14132 14172
rect 14156 14170 14212 14172
rect 14236 14170 14292 14172
rect 14316 14170 14372 14172
rect 14396 14170 14452 14172
rect 14476 14170 14532 14172
rect 14556 14170 14612 14172
rect 14636 14170 14692 14172
rect 13516 14118 13554 14170
rect 13554 14118 13566 14170
rect 13566 14118 13572 14170
rect 13596 14118 13618 14170
rect 13618 14118 13630 14170
rect 13630 14118 13652 14170
rect 13676 14118 13682 14170
rect 13682 14118 13694 14170
rect 13694 14118 13732 14170
rect 13756 14118 13758 14170
rect 13758 14118 13810 14170
rect 13810 14118 13812 14170
rect 13836 14118 13874 14170
rect 13874 14118 13886 14170
rect 13886 14118 13892 14170
rect 13916 14118 13938 14170
rect 13938 14118 13950 14170
rect 13950 14118 13972 14170
rect 13996 14118 14002 14170
rect 14002 14118 14014 14170
rect 14014 14118 14052 14170
rect 14076 14118 14078 14170
rect 14078 14118 14130 14170
rect 14130 14118 14132 14170
rect 14156 14118 14194 14170
rect 14194 14118 14206 14170
rect 14206 14118 14212 14170
rect 14236 14118 14258 14170
rect 14258 14118 14270 14170
rect 14270 14118 14292 14170
rect 14316 14118 14322 14170
rect 14322 14118 14334 14170
rect 14334 14118 14372 14170
rect 14396 14118 14398 14170
rect 14398 14118 14450 14170
rect 14450 14118 14452 14170
rect 14476 14118 14514 14170
rect 14514 14118 14526 14170
rect 14526 14118 14532 14170
rect 14556 14118 14578 14170
rect 14578 14118 14590 14170
rect 14590 14118 14612 14170
rect 14636 14118 14642 14170
rect 14642 14118 14654 14170
rect 14654 14118 14692 14170
rect 13516 14116 13572 14118
rect 13596 14116 13652 14118
rect 13676 14116 13732 14118
rect 13756 14116 13812 14118
rect 13836 14116 13892 14118
rect 13916 14116 13972 14118
rect 13996 14116 14052 14118
rect 14076 14116 14132 14118
rect 14156 14116 14212 14118
rect 14236 14116 14292 14118
rect 14316 14116 14372 14118
rect 14396 14116 14452 14118
rect 14476 14116 14532 14118
rect 14556 14116 14612 14118
rect 14636 14116 14692 14118
rect 15750 14456 15806 14512
rect 13516 13082 13572 13084
rect 13596 13082 13652 13084
rect 13676 13082 13732 13084
rect 13756 13082 13812 13084
rect 13836 13082 13892 13084
rect 13916 13082 13972 13084
rect 13996 13082 14052 13084
rect 14076 13082 14132 13084
rect 14156 13082 14212 13084
rect 14236 13082 14292 13084
rect 14316 13082 14372 13084
rect 14396 13082 14452 13084
rect 14476 13082 14532 13084
rect 14556 13082 14612 13084
rect 14636 13082 14692 13084
rect 13516 13030 13554 13082
rect 13554 13030 13566 13082
rect 13566 13030 13572 13082
rect 13596 13030 13618 13082
rect 13618 13030 13630 13082
rect 13630 13030 13652 13082
rect 13676 13030 13682 13082
rect 13682 13030 13694 13082
rect 13694 13030 13732 13082
rect 13756 13030 13758 13082
rect 13758 13030 13810 13082
rect 13810 13030 13812 13082
rect 13836 13030 13874 13082
rect 13874 13030 13886 13082
rect 13886 13030 13892 13082
rect 13916 13030 13938 13082
rect 13938 13030 13950 13082
rect 13950 13030 13972 13082
rect 13996 13030 14002 13082
rect 14002 13030 14014 13082
rect 14014 13030 14052 13082
rect 14076 13030 14078 13082
rect 14078 13030 14130 13082
rect 14130 13030 14132 13082
rect 14156 13030 14194 13082
rect 14194 13030 14206 13082
rect 14206 13030 14212 13082
rect 14236 13030 14258 13082
rect 14258 13030 14270 13082
rect 14270 13030 14292 13082
rect 14316 13030 14322 13082
rect 14322 13030 14334 13082
rect 14334 13030 14372 13082
rect 14396 13030 14398 13082
rect 14398 13030 14450 13082
rect 14450 13030 14452 13082
rect 14476 13030 14514 13082
rect 14514 13030 14526 13082
rect 14526 13030 14532 13082
rect 14556 13030 14578 13082
rect 14578 13030 14590 13082
rect 14590 13030 14612 13082
rect 14636 13030 14642 13082
rect 14642 13030 14654 13082
rect 14654 13030 14692 13082
rect 13516 13028 13572 13030
rect 13596 13028 13652 13030
rect 13676 13028 13732 13030
rect 13756 13028 13812 13030
rect 13836 13028 13892 13030
rect 13916 13028 13972 13030
rect 13996 13028 14052 13030
rect 14076 13028 14132 13030
rect 14156 13028 14212 13030
rect 14236 13028 14292 13030
rect 14316 13028 14372 13030
rect 14396 13028 14452 13030
rect 14476 13028 14532 13030
rect 14556 13028 14612 13030
rect 14636 13028 14692 13030
rect 13516 11994 13572 11996
rect 13596 11994 13652 11996
rect 13676 11994 13732 11996
rect 13756 11994 13812 11996
rect 13836 11994 13892 11996
rect 13916 11994 13972 11996
rect 13996 11994 14052 11996
rect 14076 11994 14132 11996
rect 14156 11994 14212 11996
rect 14236 11994 14292 11996
rect 14316 11994 14372 11996
rect 14396 11994 14452 11996
rect 14476 11994 14532 11996
rect 14556 11994 14612 11996
rect 14636 11994 14692 11996
rect 13516 11942 13554 11994
rect 13554 11942 13566 11994
rect 13566 11942 13572 11994
rect 13596 11942 13618 11994
rect 13618 11942 13630 11994
rect 13630 11942 13652 11994
rect 13676 11942 13682 11994
rect 13682 11942 13694 11994
rect 13694 11942 13732 11994
rect 13756 11942 13758 11994
rect 13758 11942 13810 11994
rect 13810 11942 13812 11994
rect 13836 11942 13874 11994
rect 13874 11942 13886 11994
rect 13886 11942 13892 11994
rect 13916 11942 13938 11994
rect 13938 11942 13950 11994
rect 13950 11942 13972 11994
rect 13996 11942 14002 11994
rect 14002 11942 14014 11994
rect 14014 11942 14052 11994
rect 14076 11942 14078 11994
rect 14078 11942 14130 11994
rect 14130 11942 14132 11994
rect 14156 11942 14194 11994
rect 14194 11942 14206 11994
rect 14206 11942 14212 11994
rect 14236 11942 14258 11994
rect 14258 11942 14270 11994
rect 14270 11942 14292 11994
rect 14316 11942 14322 11994
rect 14322 11942 14334 11994
rect 14334 11942 14372 11994
rect 14396 11942 14398 11994
rect 14398 11942 14450 11994
rect 14450 11942 14452 11994
rect 14476 11942 14514 11994
rect 14514 11942 14526 11994
rect 14526 11942 14532 11994
rect 14556 11942 14578 11994
rect 14578 11942 14590 11994
rect 14590 11942 14612 11994
rect 14636 11942 14642 11994
rect 14642 11942 14654 11994
rect 14654 11942 14692 11994
rect 13516 11940 13572 11942
rect 13596 11940 13652 11942
rect 13676 11940 13732 11942
rect 13756 11940 13812 11942
rect 13836 11940 13892 11942
rect 13916 11940 13972 11942
rect 13996 11940 14052 11942
rect 14076 11940 14132 11942
rect 14156 11940 14212 11942
rect 14236 11940 14292 11942
rect 14316 11940 14372 11942
rect 14396 11940 14452 11942
rect 14476 11940 14532 11942
rect 14556 11940 14612 11942
rect 14636 11940 14692 11942
rect 14462 11212 14518 11248
rect 14462 11192 14464 11212
rect 14464 11192 14516 11212
rect 14516 11192 14518 11212
rect 14646 11736 14702 11792
rect 13516 10906 13572 10908
rect 13596 10906 13652 10908
rect 13676 10906 13732 10908
rect 13756 10906 13812 10908
rect 13836 10906 13892 10908
rect 13916 10906 13972 10908
rect 13996 10906 14052 10908
rect 14076 10906 14132 10908
rect 14156 10906 14212 10908
rect 14236 10906 14292 10908
rect 14316 10906 14372 10908
rect 14396 10906 14452 10908
rect 14476 10906 14532 10908
rect 14556 10906 14612 10908
rect 14636 10906 14692 10908
rect 13516 10854 13554 10906
rect 13554 10854 13566 10906
rect 13566 10854 13572 10906
rect 13596 10854 13618 10906
rect 13618 10854 13630 10906
rect 13630 10854 13652 10906
rect 13676 10854 13682 10906
rect 13682 10854 13694 10906
rect 13694 10854 13732 10906
rect 13756 10854 13758 10906
rect 13758 10854 13810 10906
rect 13810 10854 13812 10906
rect 13836 10854 13874 10906
rect 13874 10854 13886 10906
rect 13886 10854 13892 10906
rect 13916 10854 13938 10906
rect 13938 10854 13950 10906
rect 13950 10854 13972 10906
rect 13996 10854 14002 10906
rect 14002 10854 14014 10906
rect 14014 10854 14052 10906
rect 14076 10854 14078 10906
rect 14078 10854 14130 10906
rect 14130 10854 14132 10906
rect 14156 10854 14194 10906
rect 14194 10854 14206 10906
rect 14206 10854 14212 10906
rect 14236 10854 14258 10906
rect 14258 10854 14270 10906
rect 14270 10854 14292 10906
rect 14316 10854 14322 10906
rect 14322 10854 14334 10906
rect 14334 10854 14372 10906
rect 14396 10854 14398 10906
rect 14398 10854 14450 10906
rect 14450 10854 14452 10906
rect 14476 10854 14514 10906
rect 14514 10854 14526 10906
rect 14526 10854 14532 10906
rect 14556 10854 14578 10906
rect 14578 10854 14590 10906
rect 14590 10854 14612 10906
rect 14636 10854 14642 10906
rect 14642 10854 14654 10906
rect 14654 10854 14692 10906
rect 13516 10852 13572 10854
rect 13596 10852 13652 10854
rect 13676 10852 13732 10854
rect 13756 10852 13812 10854
rect 13836 10852 13892 10854
rect 13916 10852 13972 10854
rect 13996 10852 14052 10854
rect 14076 10852 14132 10854
rect 14156 10852 14212 10854
rect 14236 10852 14292 10854
rect 14316 10852 14372 10854
rect 14396 10852 14452 10854
rect 14476 10852 14532 10854
rect 14556 10852 14612 10854
rect 14636 10852 14692 10854
rect 13266 9868 13268 9888
rect 13268 9868 13320 9888
rect 13320 9868 13322 9888
rect 13266 9832 13322 9868
rect 14738 10512 14794 10568
rect 14462 10104 14518 10160
rect 14278 9968 14334 10024
rect 13516 9818 13572 9820
rect 13596 9818 13652 9820
rect 13676 9818 13732 9820
rect 13756 9818 13812 9820
rect 13836 9818 13892 9820
rect 13916 9818 13972 9820
rect 13996 9818 14052 9820
rect 14076 9818 14132 9820
rect 14156 9818 14212 9820
rect 14236 9818 14292 9820
rect 14316 9818 14372 9820
rect 14396 9818 14452 9820
rect 14476 9818 14532 9820
rect 14556 9818 14612 9820
rect 14636 9818 14692 9820
rect 13516 9766 13554 9818
rect 13554 9766 13566 9818
rect 13566 9766 13572 9818
rect 13596 9766 13618 9818
rect 13618 9766 13630 9818
rect 13630 9766 13652 9818
rect 13676 9766 13682 9818
rect 13682 9766 13694 9818
rect 13694 9766 13732 9818
rect 13756 9766 13758 9818
rect 13758 9766 13810 9818
rect 13810 9766 13812 9818
rect 13836 9766 13874 9818
rect 13874 9766 13886 9818
rect 13886 9766 13892 9818
rect 13916 9766 13938 9818
rect 13938 9766 13950 9818
rect 13950 9766 13972 9818
rect 13996 9766 14002 9818
rect 14002 9766 14014 9818
rect 14014 9766 14052 9818
rect 14076 9766 14078 9818
rect 14078 9766 14130 9818
rect 14130 9766 14132 9818
rect 14156 9766 14194 9818
rect 14194 9766 14206 9818
rect 14206 9766 14212 9818
rect 14236 9766 14258 9818
rect 14258 9766 14270 9818
rect 14270 9766 14292 9818
rect 14316 9766 14322 9818
rect 14322 9766 14334 9818
rect 14334 9766 14372 9818
rect 14396 9766 14398 9818
rect 14398 9766 14450 9818
rect 14450 9766 14452 9818
rect 14476 9766 14514 9818
rect 14514 9766 14526 9818
rect 14526 9766 14532 9818
rect 14556 9766 14578 9818
rect 14578 9766 14590 9818
rect 14590 9766 14612 9818
rect 14636 9766 14642 9818
rect 14642 9766 14654 9818
rect 14654 9766 14692 9818
rect 13516 9764 13572 9766
rect 13596 9764 13652 9766
rect 13676 9764 13732 9766
rect 13756 9764 13812 9766
rect 13836 9764 13892 9766
rect 13916 9764 13972 9766
rect 13996 9764 14052 9766
rect 14076 9764 14132 9766
rect 14156 9764 14212 9766
rect 14236 9764 14292 9766
rect 14316 9764 14372 9766
rect 14396 9764 14452 9766
rect 14476 9764 14532 9766
rect 14556 9764 14612 9766
rect 14636 9764 14692 9766
rect 13174 8900 13230 8936
rect 13174 8880 13176 8900
rect 13176 8880 13228 8900
rect 13228 8880 13230 8900
rect 13174 8744 13230 8800
rect 12714 3712 12770 3768
rect 12990 3168 13046 3224
rect 12714 2932 12716 2952
rect 12716 2932 12768 2952
rect 12768 2932 12770 2952
rect 12714 2896 12770 2932
rect 13358 9560 13414 9616
rect 13818 9424 13874 9480
rect 13542 9152 13598 9208
rect 13818 8880 13874 8936
rect 14646 9560 14702 9616
rect 14554 8880 14610 8936
rect 13516 8730 13572 8732
rect 13596 8730 13652 8732
rect 13676 8730 13732 8732
rect 13756 8730 13812 8732
rect 13836 8730 13892 8732
rect 13916 8730 13972 8732
rect 13996 8730 14052 8732
rect 14076 8730 14132 8732
rect 14156 8730 14212 8732
rect 14236 8730 14292 8732
rect 14316 8730 14372 8732
rect 14396 8730 14452 8732
rect 14476 8730 14532 8732
rect 14556 8730 14612 8732
rect 14636 8730 14692 8732
rect 13516 8678 13554 8730
rect 13554 8678 13566 8730
rect 13566 8678 13572 8730
rect 13596 8678 13618 8730
rect 13618 8678 13630 8730
rect 13630 8678 13652 8730
rect 13676 8678 13682 8730
rect 13682 8678 13694 8730
rect 13694 8678 13732 8730
rect 13756 8678 13758 8730
rect 13758 8678 13810 8730
rect 13810 8678 13812 8730
rect 13836 8678 13874 8730
rect 13874 8678 13886 8730
rect 13886 8678 13892 8730
rect 13916 8678 13938 8730
rect 13938 8678 13950 8730
rect 13950 8678 13972 8730
rect 13996 8678 14002 8730
rect 14002 8678 14014 8730
rect 14014 8678 14052 8730
rect 14076 8678 14078 8730
rect 14078 8678 14130 8730
rect 14130 8678 14132 8730
rect 14156 8678 14194 8730
rect 14194 8678 14206 8730
rect 14206 8678 14212 8730
rect 14236 8678 14258 8730
rect 14258 8678 14270 8730
rect 14270 8678 14292 8730
rect 14316 8678 14322 8730
rect 14322 8678 14334 8730
rect 14334 8678 14372 8730
rect 14396 8678 14398 8730
rect 14398 8678 14450 8730
rect 14450 8678 14452 8730
rect 14476 8678 14514 8730
rect 14514 8678 14526 8730
rect 14526 8678 14532 8730
rect 14556 8678 14578 8730
rect 14578 8678 14590 8730
rect 14590 8678 14612 8730
rect 14636 8678 14642 8730
rect 14642 8678 14654 8730
rect 14654 8678 14692 8730
rect 13516 8676 13572 8678
rect 13596 8676 13652 8678
rect 13676 8676 13732 8678
rect 13756 8676 13812 8678
rect 13836 8676 13892 8678
rect 13916 8676 13972 8678
rect 13996 8676 14052 8678
rect 14076 8676 14132 8678
rect 14156 8676 14212 8678
rect 14236 8676 14292 8678
rect 14316 8676 14372 8678
rect 14396 8676 14452 8678
rect 14476 8676 14532 8678
rect 14556 8676 14612 8678
rect 14636 8676 14692 8678
rect 14094 8472 14150 8528
rect 14554 7828 14556 7848
rect 14556 7828 14608 7848
rect 14608 7828 14610 7848
rect 14554 7792 14610 7828
rect 13516 7642 13572 7644
rect 13596 7642 13652 7644
rect 13676 7642 13732 7644
rect 13756 7642 13812 7644
rect 13836 7642 13892 7644
rect 13916 7642 13972 7644
rect 13996 7642 14052 7644
rect 14076 7642 14132 7644
rect 14156 7642 14212 7644
rect 14236 7642 14292 7644
rect 14316 7642 14372 7644
rect 14396 7642 14452 7644
rect 14476 7642 14532 7644
rect 14556 7642 14612 7644
rect 14636 7642 14692 7644
rect 13516 7590 13554 7642
rect 13554 7590 13566 7642
rect 13566 7590 13572 7642
rect 13596 7590 13618 7642
rect 13618 7590 13630 7642
rect 13630 7590 13652 7642
rect 13676 7590 13682 7642
rect 13682 7590 13694 7642
rect 13694 7590 13732 7642
rect 13756 7590 13758 7642
rect 13758 7590 13810 7642
rect 13810 7590 13812 7642
rect 13836 7590 13874 7642
rect 13874 7590 13886 7642
rect 13886 7590 13892 7642
rect 13916 7590 13938 7642
rect 13938 7590 13950 7642
rect 13950 7590 13972 7642
rect 13996 7590 14002 7642
rect 14002 7590 14014 7642
rect 14014 7590 14052 7642
rect 14076 7590 14078 7642
rect 14078 7590 14130 7642
rect 14130 7590 14132 7642
rect 14156 7590 14194 7642
rect 14194 7590 14206 7642
rect 14206 7590 14212 7642
rect 14236 7590 14258 7642
rect 14258 7590 14270 7642
rect 14270 7590 14292 7642
rect 14316 7590 14322 7642
rect 14322 7590 14334 7642
rect 14334 7590 14372 7642
rect 14396 7590 14398 7642
rect 14398 7590 14450 7642
rect 14450 7590 14452 7642
rect 14476 7590 14514 7642
rect 14514 7590 14526 7642
rect 14526 7590 14532 7642
rect 14556 7590 14578 7642
rect 14578 7590 14590 7642
rect 14590 7590 14612 7642
rect 14636 7590 14642 7642
rect 14642 7590 14654 7642
rect 14654 7590 14692 7642
rect 13516 7588 13572 7590
rect 13596 7588 13652 7590
rect 13676 7588 13732 7590
rect 13756 7588 13812 7590
rect 13836 7588 13892 7590
rect 13916 7588 13972 7590
rect 13996 7588 14052 7590
rect 14076 7588 14132 7590
rect 14156 7588 14212 7590
rect 14236 7588 14292 7590
rect 14316 7588 14372 7590
rect 14396 7588 14452 7590
rect 14476 7588 14532 7590
rect 14556 7588 14612 7590
rect 14636 7588 14692 7590
rect 14830 8336 14886 8392
rect 13516 6554 13572 6556
rect 13596 6554 13652 6556
rect 13676 6554 13732 6556
rect 13756 6554 13812 6556
rect 13836 6554 13892 6556
rect 13916 6554 13972 6556
rect 13996 6554 14052 6556
rect 14076 6554 14132 6556
rect 14156 6554 14212 6556
rect 14236 6554 14292 6556
rect 14316 6554 14372 6556
rect 14396 6554 14452 6556
rect 14476 6554 14532 6556
rect 14556 6554 14612 6556
rect 14636 6554 14692 6556
rect 13516 6502 13554 6554
rect 13554 6502 13566 6554
rect 13566 6502 13572 6554
rect 13596 6502 13618 6554
rect 13618 6502 13630 6554
rect 13630 6502 13652 6554
rect 13676 6502 13682 6554
rect 13682 6502 13694 6554
rect 13694 6502 13732 6554
rect 13756 6502 13758 6554
rect 13758 6502 13810 6554
rect 13810 6502 13812 6554
rect 13836 6502 13874 6554
rect 13874 6502 13886 6554
rect 13886 6502 13892 6554
rect 13916 6502 13938 6554
rect 13938 6502 13950 6554
rect 13950 6502 13972 6554
rect 13996 6502 14002 6554
rect 14002 6502 14014 6554
rect 14014 6502 14052 6554
rect 14076 6502 14078 6554
rect 14078 6502 14130 6554
rect 14130 6502 14132 6554
rect 14156 6502 14194 6554
rect 14194 6502 14206 6554
rect 14206 6502 14212 6554
rect 14236 6502 14258 6554
rect 14258 6502 14270 6554
rect 14270 6502 14292 6554
rect 14316 6502 14322 6554
rect 14322 6502 14334 6554
rect 14334 6502 14372 6554
rect 14396 6502 14398 6554
rect 14398 6502 14450 6554
rect 14450 6502 14452 6554
rect 14476 6502 14514 6554
rect 14514 6502 14526 6554
rect 14526 6502 14532 6554
rect 14556 6502 14578 6554
rect 14578 6502 14590 6554
rect 14590 6502 14612 6554
rect 14636 6502 14642 6554
rect 14642 6502 14654 6554
rect 14654 6502 14692 6554
rect 13516 6500 13572 6502
rect 13596 6500 13652 6502
rect 13676 6500 13732 6502
rect 13756 6500 13812 6502
rect 13836 6500 13892 6502
rect 13916 6500 13972 6502
rect 13996 6500 14052 6502
rect 14076 6500 14132 6502
rect 14156 6500 14212 6502
rect 14236 6500 14292 6502
rect 14316 6500 14372 6502
rect 14396 6500 14452 6502
rect 14476 6500 14532 6502
rect 14556 6500 14612 6502
rect 14636 6500 14692 6502
rect 14554 6332 14556 6352
rect 14556 6332 14608 6352
rect 14608 6332 14610 6352
rect 14554 6296 14610 6332
rect 14554 6024 14610 6080
rect 13516 5466 13572 5468
rect 13596 5466 13652 5468
rect 13676 5466 13732 5468
rect 13756 5466 13812 5468
rect 13836 5466 13892 5468
rect 13916 5466 13972 5468
rect 13996 5466 14052 5468
rect 14076 5466 14132 5468
rect 14156 5466 14212 5468
rect 14236 5466 14292 5468
rect 14316 5466 14372 5468
rect 14396 5466 14452 5468
rect 14476 5466 14532 5468
rect 14556 5466 14612 5468
rect 14636 5466 14692 5468
rect 13516 5414 13554 5466
rect 13554 5414 13566 5466
rect 13566 5414 13572 5466
rect 13596 5414 13618 5466
rect 13618 5414 13630 5466
rect 13630 5414 13652 5466
rect 13676 5414 13682 5466
rect 13682 5414 13694 5466
rect 13694 5414 13732 5466
rect 13756 5414 13758 5466
rect 13758 5414 13810 5466
rect 13810 5414 13812 5466
rect 13836 5414 13874 5466
rect 13874 5414 13886 5466
rect 13886 5414 13892 5466
rect 13916 5414 13938 5466
rect 13938 5414 13950 5466
rect 13950 5414 13972 5466
rect 13996 5414 14002 5466
rect 14002 5414 14014 5466
rect 14014 5414 14052 5466
rect 14076 5414 14078 5466
rect 14078 5414 14130 5466
rect 14130 5414 14132 5466
rect 14156 5414 14194 5466
rect 14194 5414 14206 5466
rect 14206 5414 14212 5466
rect 14236 5414 14258 5466
rect 14258 5414 14270 5466
rect 14270 5414 14292 5466
rect 14316 5414 14322 5466
rect 14322 5414 14334 5466
rect 14334 5414 14372 5466
rect 14396 5414 14398 5466
rect 14398 5414 14450 5466
rect 14450 5414 14452 5466
rect 14476 5414 14514 5466
rect 14514 5414 14526 5466
rect 14526 5414 14532 5466
rect 14556 5414 14578 5466
rect 14578 5414 14590 5466
rect 14590 5414 14612 5466
rect 14636 5414 14642 5466
rect 14642 5414 14654 5466
rect 14654 5414 14692 5466
rect 13516 5412 13572 5414
rect 13596 5412 13652 5414
rect 13676 5412 13732 5414
rect 13756 5412 13812 5414
rect 13836 5412 13892 5414
rect 13916 5412 13972 5414
rect 13996 5412 14052 5414
rect 14076 5412 14132 5414
rect 14156 5412 14212 5414
rect 14236 5412 14292 5414
rect 14316 5412 14372 5414
rect 14396 5412 14452 5414
rect 14476 5412 14532 5414
rect 14556 5412 14612 5414
rect 14636 5412 14692 5414
rect 13516 4378 13572 4380
rect 13596 4378 13652 4380
rect 13676 4378 13732 4380
rect 13756 4378 13812 4380
rect 13836 4378 13892 4380
rect 13916 4378 13972 4380
rect 13996 4378 14052 4380
rect 14076 4378 14132 4380
rect 14156 4378 14212 4380
rect 14236 4378 14292 4380
rect 14316 4378 14372 4380
rect 14396 4378 14452 4380
rect 14476 4378 14532 4380
rect 14556 4378 14612 4380
rect 14636 4378 14692 4380
rect 13516 4326 13554 4378
rect 13554 4326 13566 4378
rect 13566 4326 13572 4378
rect 13596 4326 13618 4378
rect 13618 4326 13630 4378
rect 13630 4326 13652 4378
rect 13676 4326 13682 4378
rect 13682 4326 13694 4378
rect 13694 4326 13732 4378
rect 13756 4326 13758 4378
rect 13758 4326 13810 4378
rect 13810 4326 13812 4378
rect 13836 4326 13874 4378
rect 13874 4326 13886 4378
rect 13886 4326 13892 4378
rect 13916 4326 13938 4378
rect 13938 4326 13950 4378
rect 13950 4326 13972 4378
rect 13996 4326 14002 4378
rect 14002 4326 14014 4378
rect 14014 4326 14052 4378
rect 14076 4326 14078 4378
rect 14078 4326 14130 4378
rect 14130 4326 14132 4378
rect 14156 4326 14194 4378
rect 14194 4326 14206 4378
rect 14206 4326 14212 4378
rect 14236 4326 14258 4378
rect 14258 4326 14270 4378
rect 14270 4326 14292 4378
rect 14316 4326 14322 4378
rect 14322 4326 14334 4378
rect 14334 4326 14372 4378
rect 14396 4326 14398 4378
rect 14398 4326 14450 4378
rect 14450 4326 14452 4378
rect 14476 4326 14514 4378
rect 14514 4326 14526 4378
rect 14526 4326 14532 4378
rect 14556 4326 14578 4378
rect 14578 4326 14590 4378
rect 14590 4326 14612 4378
rect 14636 4326 14642 4378
rect 14642 4326 14654 4378
rect 14654 4326 14692 4378
rect 13516 4324 13572 4326
rect 13596 4324 13652 4326
rect 13676 4324 13732 4326
rect 13756 4324 13812 4326
rect 13836 4324 13892 4326
rect 13916 4324 13972 4326
rect 13996 4324 14052 4326
rect 14076 4324 14132 4326
rect 14156 4324 14212 4326
rect 14236 4324 14292 4326
rect 14316 4324 14372 4326
rect 14396 4324 14452 4326
rect 14476 4324 14532 4326
rect 14556 4324 14612 4326
rect 14636 4324 14692 4326
rect 14186 3984 14242 4040
rect 14646 3712 14702 3768
rect 14278 3460 14334 3496
rect 14278 3440 14280 3460
rect 14280 3440 14332 3460
rect 14332 3440 14334 3460
rect 14462 3476 14464 3496
rect 14464 3476 14516 3496
rect 14516 3476 14518 3496
rect 14462 3440 14518 3476
rect 13516 3290 13572 3292
rect 13596 3290 13652 3292
rect 13676 3290 13732 3292
rect 13756 3290 13812 3292
rect 13836 3290 13892 3292
rect 13916 3290 13972 3292
rect 13996 3290 14052 3292
rect 14076 3290 14132 3292
rect 14156 3290 14212 3292
rect 14236 3290 14292 3292
rect 14316 3290 14372 3292
rect 14396 3290 14452 3292
rect 14476 3290 14532 3292
rect 14556 3290 14612 3292
rect 14636 3290 14692 3292
rect 13516 3238 13554 3290
rect 13554 3238 13566 3290
rect 13566 3238 13572 3290
rect 13596 3238 13618 3290
rect 13618 3238 13630 3290
rect 13630 3238 13652 3290
rect 13676 3238 13682 3290
rect 13682 3238 13694 3290
rect 13694 3238 13732 3290
rect 13756 3238 13758 3290
rect 13758 3238 13810 3290
rect 13810 3238 13812 3290
rect 13836 3238 13874 3290
rect 13874 3238 13886 3290
rect 13886 3238 13892 3290
rect 13916 3238 13938 3290
rect 13938 3238 13950 3290
rect 13950 3238 13972 3290
rect 13996 3238 14002 3290
rect 14002 3238 14014 3290
rect 14014 3238 14052 3290
rect 14076 3238 14078 3290
rect 14078 3238 14130 3290
rect 14130 3238 14132 3290
rect 14156 3238 14194 3290
rect 14194 3238 14206 3290
rect 14206 3238 14212 3290
rect 14236 3238 14258 3290
rect 14258 3238 14270 3290
rect 14270 3238 14292 3290
rect 14316 3238 14322 3290
rect 14322 3238 14334 3290
rect 14334 3238 14372 3290
rect 14396 3238 14398 3290
rect 14398 3238 14450 3290
rect 14450 3238 14452 3290
rect 14476 3238 14514 3290
rect 14514 3238 14526 3290
rect 14526 3238 14532 3290
rect 14556 3238 14578 3290
rect 14578 3238 14590 3290
rect 14590 3238 14612 3290
rect 14636 3238 14642 3290
rect 14642 3238 14654 3290
rect 14654 3238 14692 3290
rect 13516 3236 13572 3238
rect 13596 3236 13652 3238
rect 13676 3236 13732 3238
rect 13756 3236 13812 3238
rect 13836 3236 13892 3238
rect 13916 3236 13972 3238
rect 13996 3236 14052 3238
rect 14076 3236 14132 3238
rect 14156 3236 14212 3238
rect 14236 3236 14292 3238
rect 14316 3236 14372 3238
rect 14396 3236 14452 3238
rect 14476 3236 14532 3238
rect 14556 3236 14612 3238
rect 14636 3236 14692 3238
rect 13082 2508 13138 2544
rect 13082 2488 13084 2508
rect 13084 2488 13136 2508
rect 13136 2488 13138 2508
rect 13516 2202 13572 2204
rect 13596 2202 13652 2204
rect 13676 2202 13732 2204
rect 13756 2202 13812 2204
rect 13836 2202 13892 2204
rect 13916 2202 13972 2204
rect 13996 2202 14052 2204
rect 14076 2202 14132 2204
rect 14156 2202 14212 2204
rect 14236 2202 14292 2204
rect 14316 2202 14372 2204
rect 14396 2202 14452 2204
rect 14476 2202 14532 2204
rect 14556 2202 14612 2204
rect 14636 2202 14692 2204
rect 13516 2150 13554 2202
rect 13554 2150 13566 2202
rect 13566 2150 13572 2202
rect 13596 2150 13618 2202
rect 13618 2150 13630 2202
rect 13630 2150 13652 2202
rect 13676 2150 13682 2202
rect 13682 2150 13694 2202
rect 13694 2150 13732 2202
rect 13756 2150 13758 2202
rect 13758 2150 13810 2202
rect 13810 2150 13812 2202
rect 13836 2150 13874 2202
rect 13874 2150 13886 2202
rect 13886 2150 13892 2202
rect 13916 2150 13938 2202
rect 13938 2150 13950 2202
rect 13950 2150 13972 2202
rect 13996 2150 14002 2202
rect 14002 2150 14014 2202
rect 14014 2150 14052 2202
rect 14076 2150 14078 2202
rect 14078 2150 14130 2202
rect 14130 2150 14132 2202
rect 14156 2150 14194 2202
rect 14194 2150 14206 2202
rect 14206 2150 14212 2202
rect 14236 2150 14258 2202
rect 14258 2150 14270 2202
rect 14270 2150 14292 2202
rect 14316 2150 14322 2202
rect 14322 2150 14334 2202
rect 14334 2150 14372 2202
rect 14396 2150 14398 2202
rect 14398 2150 14450 2202
rect 14450 2150 14452 2202
rect 14476 2150 14514 2202
rect 14514 2150 14526 2202
rect 14526 2150 14532 2202
rect 14556 2150 14578 2202
rect 14578 2150 14590 2202
rect 14590 2150 14612 2202
rect 14636 2150 14642 2202
rect 14642 2150 14654 2202
rect 14654 2150 14692 2202
rect 13516 2148 13572 2150
rect 13596 2148 13652 2150
rect 13676 2148 13732 2150
rect 13756 2148 13812 2150
rect 13836 2148 13892 2150
rect 13916 2148 13972 2150
rect 13996 2148 14052 2150
rect 14076 2148 14132 2150
rect 14156 2148 14212 2150
rect 14236 2148 14292 2150
rect 14316 2148 14372 2150
rect 14396 2148 14452 2150
rect 14476 2148 14532 2150
rect 14556 2148 14612 2150
rect 14636 2148 14692 2150
rect 15106 11192 15162 11248
rect 15290 11192 15346 11248
rect 15382 8064 15438 8120
rect 15198 6704 15254 6760
rect 15474 6976 15530 7032
rect 15750 9560 15806 9616
rect 15750 9460 15752 9480
rect 15752 9460 15804 9480
rect 15804 9460 15806 9480
rect 15750 9424 15806 9460
rect 15566 6296 15622 6352
rect 15382 6024 15438 6080
rect 16026 10512 16082 10568
rect 16026 6704 16082 6760
rect 17516 15802 17572 15804
rect 17596 15802 17652 15804
rect 17676 15802 17732 15804
rect 17756 15802 17812 15804
rect 17836 15802 17892 15804
rect 17916 15802 17972 15804
rect 17996 15802 18052 15804
rect 18076 15802 18132 15804
rect 18156 15802 18212 15804
rect 18236 15802 18292 15804
rect 18316 15802 18372 15804
rect 18396 15802 18452 15804
rect 18476 15802 18532 15804
rect 18556 15802 18612 15804
rect 18636 15802 18692 15804
rect 17516 15750 17554 15802
rect 17554 15750 17566 15802
rect 17566 15750 17572 15802
rect 17596 15750 17618 15802
rect 17618 15750 17630 15802
rect 17630 15750 17652 15802
rect 17676 15750 17682 15802
rect 17682 15750 17694 15802
rect 17694 15750 17732 15802
rect 17756 15750 17758 15802
rect 17758 15750 17810 15802
rect 17810 15750 17812 15802
rect 17836 15750 17874 15802
rect 17874 15750 17886 15802
rect 17886 15750 17892 15802
rect 17916 15750 17938 15802
rect 17938 15750 17950 15802
rect 17950 15750 17972 15802
rect 17996 15750 18002 15802
rect 18002 15750 18014 15802
rect 18014 15750 18052 15802
rect 18076 15750 18078 15802
rect 18078 15750 18130 15802
rect 18130 15750 18132 15802
rect 18156 15750 18194 15802
rect 18194 15750 18206 15802
rect 18206 15750 18212 15802
rect 18236 15750 18258 15802
rect 18258 15750 18270 15802
rect 18270 15750 18292 15802
rect 18316 15750 18322 15802
rect 18322 15750 18334 15802
rect 18334 15750 18372 15802
rect 18396 15750 18398 15802
rect 18398 15750 18450 15802
rect 18450 15750 18452 15802
rect 18476 15750 18514 15802
rect 18514 15750 18526 15802
rect 18526 15750 18532 15802
rect 18556 15750 18578 15802
rect 18578 15750 18590 15802
rect 18590 15750 18612 15802
rect 18636 15750 18642 15802
rect 18642 15750 18654 15802
rect 18654 15750 18692 15802
rect 17516 15748 17572 15750
rect 17596 15748 17652 15750
rect 17676 15748 17732 15750
rect 17756 15748 17812 15750
rect 17836 15748 17892 15750
rect 17916 15748 17972 15750
rect 17996 15748 18052 15750
rect 18076 15748 18132 15750
rect 18156 15748 18212 15750
rect 18236 15748 18292 15750
rect 18316 15748 18372 15750
rect 18396 15748 18452 15750
rect 18476 15748 18532 15750
rect 18556 15748 18612 15750
rect 18636 15748 18692 15750
rect 17516 14714 17572 14716
rect 17596 14714 17652 14716
rect 17676 14714 17732 14716
rect 17756 14714 17812 14716
rect 17836 14714 17892 14716
rect 17916 14714 17972 14716
rect 17996 14714 18052 14716
rect 18076 14714 18132 14716
rect 18156 14714 18212 14716
rect 18236 14714 18292 14716
rect 18316 14714 18372 14716
rect 18396 14714 18452 14716
rect 18476 14714 18532 14716
rect 18556 14714 18612 14716
rect 18636 14714 18692 14716
rect 17516 14662 17554 14714
rect 17554 14662 17566 14714
rect 17566 14662 17572 14714
rect 17596 14662 17618 14714
rect 17618 14662 17630 14714
rect 17630 14662 17652 14714
rect 17676 14662 17682 14714
rect 17682 14662 17694 14714
rect 17694 14662 17732 14714
rect 17756 14662 17758 14714
rect 17758 14662 17810 14714
rect 17810 14662 17812 14714
rect 17836 14662 17874 14714
rect 17874 14662 17886 14714
rect 17886 14662 17892 14714
rect 17916 14662 17938 14714
rect 17938 14662 17950 14714
rect 17950 14662 17972 14714
rect 17996 14662 18002 14714
rect 18002 14662 18014 14714
rect 18014 14662 18052 14714
rect 18076 14662 18078 14714
rect 18078 14662 18130 14714
rect 18130 14662 18132 14714
rect 18156 14662 18194 14714
rect 18194 14662 18206 14714
rect 18206 14662 18212 14714
rect 18236 14662 18258 14714
rect 18258 14662 18270 14714
rect 18270 14662 18292 14714
rect 18316 14662 18322 14714
rect 18322 14662 18334 14714
rect 18334 14662 18372 14714
rect 18396 14662 18398 14714
rect 18398 14662 18450 14714
rect 18450 14662 18452 14714
rect 18476 14662 18514 14714
rect 18514 14662 18526 14714
rect 18526 14662 18532 14714
rect 18556 14662 18578 14714
rect 18578 14662 18590 14714
rect 18590 14662 18612 14714
rect 18636 14662 18642 14714
rect 18642 14662 18654 14714
rect 18654 14662 18692 14714
rect 17516 14660 17572 14662
rect 17596 14660 17652 14662
rect 17676 14660 17732 14662
rect 17756 14660 17812 14662
rect 17836 14660 17892 14662
rect 17916 14660 17972 14662
rect 17996 14660 18052 14662
rect 18076 14660 18132 14662
rect 18156 14660 18212 14662
rect 18236 14660 18292 14662
rect 18316 14660 18372 14662
rect 18396 14660 18452 14662
rect 18476 14660 18532 14662
rect 18556 14660 18612 14662
rect 18636 14660 18692 14662
rect 17516 13626 17572 13628
rect 17596 13626 17652 13628
rect 17676 13626 17732 13628
rect 17756 13626 17812 13628
rect 17836 13626 17892 13628
rect 17916 13626 17972 13628
rect 17996 13626 18052 13628
rect 18076 13626 18132 13628
rect 18156 13626 18212 13628
rect 18236 13626 18292 13628
rect 18316 13626 18372 13628
rect 18396 13626 18452 13628
rect 18476 13626 18532 13628
rect 18556 13626 18612 13628
rect 18636 13626 18692 13628
rect 17516 13574 17554 13626
rect 17554 13574 17566 13626
rect 17566 13574 17572 13626
rect 17596 13574 17618 13626
rect 17618 13574 17630 13626
rect 17630 13574 17652 13626
rect 17676 13574 17682 13626
rect 17682 13574 17694 13626
rect 17694 13574 17732 13626
rect 17756 13574 17758 13626
rect 17758 13574 17810 13626
rect 17810 13574 17812 13626
rect 17836 13574 17874 13626
rect 17874 13574 17886 13626
rect 17886 13574 17892 13626
rect 17916 13574 17938 13626
rect 17938 13574 17950 13626
rect 17950 13574 17972 13626
rect 17996 13574 18002 13626
rect 18002 13574 18014 13626
rect 18014 13574 18052 13626
rect 18076 13574 18078 13626
rect 18078 13574 18130 13626
rect 18130 13574 18132 13626
rect 18156 13574 18194 13626
rect 18194 13574 18206 13626
rect 18206 13574 18212 13626
rect 18236 13574 18258 13626
rect 18258 13574 18270 13626
rect 18270 13574 18292 13626
rect 18316 13574 18322 13626
rect 18322 13574 18334 13626
rect 18334 13574 18372 13626
rect 18396 13574 18398 13626
rect 18398 13574 18450 13626
rect 18450 13574 18452 13626
rect 18476 13574 18514 13626
rect 18514 13574 18526 13626
rect 18526 13574 18532 13626
rect 18556 13574 18578 13626
rect 18578 13574 18590 13626
rect 18590 13574 18612 13626
rect 18636 13574 18642 13626
rect 18642 13574 18654 13626
rect 18654 13574 18692 13626
rect 17516 13572 17572 13574
rect 17596 13572 17652 13574
rect 17676 13572 17732 13574
rect 17756 13572 17812 13574
rect 17836 13572 17892 13574
rect 17916 13572 17972 13574
rect 17996 13572 18052 13574
rect 18076 13572 18132 13574
rect 18156 13572 18212 13574
rect 18236 13572 18292 13574
rect 18316 13572 18372 13574
rect 18396 13572 18452 13574
rect 18476 13572 18532 13574
rect 18556 13572 18612 13574
rect 18636 13572 18692 13574
rect 16210 9288 16266 9344
rect 16210 7112 16266 7168
rect 15106 2760 15162 2816
rect 16486 6704 16542 6760
rect 16394 5480 16450 5536
rect 16670 10920 16726 10976
rect 17516 12538 17572 12540
rect 17596 12538 17652 12540
rect 17676 12538 17732 12540
rect 17756 12538 17812 12540
rect 17836 12538 17892 12540
rect 17916 12538 17972 12540
rect 17996 12538 18052 12540
rect 18076 12538 18132 12540
rect 18156 12538 18212 12540
rect 18236 12538 18292 12540
rect 18316 12538 18372 12540
rect 18396 12538 18452 12540
rect 18476 12538 18532 12540
rect 18556 12538 18612 12540
rect 18636 12538 18692 12540
rect 17516 12486 17554 12538
rect 17554 12486 17566 12538
rect 17566 12486 17572 12538
rect 17596 12486 17618 12538
rect 17618 12486 17630 12538
rect 17630 12486 17652 12538
rect 17676 12486 17682 12538
rect 17682 12486 17694 12538
rect 17694 12486 17732 12538
rect 17756 12486 17758 12538
rect 17758 12486 17810 12538
rect 17810 12486 17812 12538
rect 17836 12486 17874 12538
rect 17874 12486 17886 12538
rect 17886 12486 17892 12538
rect 17916 12486 17938 12538
rect 17938 12486 17950 12538
rect 17950 12486 17972 12538
rect 17996 12486 18002 12538
rect 18002 12486 18014 12538
rect 18014 12486 18052 12538
rect 18076 12486 18078 12538
rect 18078 12486 18130 12538
rect 18130 12486 18132 12538
rect 18156 12486 18194 12538
rect 18194 12486 18206 12538
rect 18206 12486 18212 12538
rect 18236 12486 18258 12538
rect 18258 12486 18270 12538
rect 18270 12486 18292 12538
rect 18316 12486 18322 12538
rect 18322 12486 18334 12538
rect 18334 12486 18372 12538
rect 18396 12486 18398 12538
rect 18398 12486 18450 12538
rect 18450 12486 18452 12538
rect 18476 12486 18514 12538
rect 18514 12486 18526 12538
rect 18526 12486 18532 12538
rect 18556 12486 18578 12538
rect 18578 12486 18590 12538
rect 18590 12486 18612 12538
rect 18636 12486 18642 12538
rect 18642 12486 18654 12538
rect 18654 12486 18692 12538
rect 17516 12484 17572 12486
rect 17596 12484 17652 12486
rect 17676 12484 17732 12486
rect 17756 12484 17812 12486
rect 17836 12484 17892 12486
rect 17916 12484 17972 12486
rect 17996 12484 18052 12486
rect 18076 12484 18132 12486
rect 18156 12484 18212 12486
rect 18236 12484 18292 12486
rect 18316 12484 18372 12486
rect 18396 12484 18452 12486
rect 18476 12484 18532 12486
rect 18556 12484 18612 12486
rect 18636 12484 18692 12486
rect 16854 11192 16910 11248
rect 18694 11600 18750 11656
rect 17516 11450 17572 11452
rect 17596 11450 17652 11452
rect 17676 11450 17732 11452
rect 17756 11450 17812 11452
rect 17836 11450 17892 11452
rect 17916 11450 17972 11452
rect 17996 11450 18052 11452
rect 18076 11450 18132 11452
rect 18156 11450 18212 11452
rect 18236 11450 18292 11452
rect 18316 11450 18372 11452
rect 18396 11450 18452 11452
rect 18476 11450 18532 11452
rect 18556 11450 18612 11452
rect 18636 11450 18692 11452
rect 17516 11398 17554 11450
rect 17554 11398 17566 11450
rect 17566 11398 17572 11450
rect 17596 11398 17618 11450
rect 17618 11398 17630 11450
rect 17630 11398 17652 11450
rect 17676 11398 17682 11450
rect 17682 11398 17694 11450
rect 17694 11398 17732 11450
rect 17756 11398 17758 11450
rect 17758 11398 17810 11450
rect 17810 11398 17812 11450
rect 17836 11398 17874 11450
rect 17874 11398 17886 11450
rect 17886 11398 17892 11450
rect 17916 11398 17938 11450
rect 17938 11398 17950 11450
rect 17950 11398 17972 11450
rect 17996 11398 18002 11450
rect 18002 11398 18014 11450
rect 18014 11398 18052 11450
rect 18076 11398 18078 11450
rect 18078 11398 18130 11450
rect 18130 11398 18132 11450
rect 18156 11398 18194 11450
rect 18194 11398 18206 11450
rect 18206 11398 18212 11450
rect 18236 11398 18258 11450
rect 18258 11398 18270 11450
rect 18270 11398 18292 11450
rect 18316 11398 18322 11450
rect 18322 11398 18334 11450
rect 18334 11398 18372 11450
rect 18396 11398 18398 11450
rect 18398 11398 18450 11450
rect 18450 11398 18452 11450
rect 18476 11398 18514 11450
rect 18514 11398 18526 11450
rect 18526 11398 18532 11450
rect 18556 11398 18578 11450
rect 18578 11398 18590 11450
rect 18590 11398 18612 11450
rect 18636 11398 18642 11450
rect 18642 11398 18654 11450
rect 18654 11398 18692 11450
rect 17516 11396 17572 11398
rect 17596 11396 17652 11398
rect 17676 11396 17732 11398
rect 17756 11396 17812 11398
rect 17836 11396 17892 11398
rect 17916 11396 17972 11398
rect 17996 11396 18052 11398
rect 18076 11396 18132 11398
rect 18156 11396 18212 11398
rect 18236 11396 18292 11398
rect 18316 11396 18372 11398
rect 18396 11396 18452 11398
rect 18476 11396 18532 11398
rect 18556 11396 18612 11398
rect 18636 11396 18692 11398
rect 17516 10362 17572 10364
rect 17596 10362 17652 10364
rect 17676 10362 17732 10364
rect 17756 10362 17812 10364
rect 17836 10362 17892 10364
rect 17916 10362 17972 10364
rect 17996 10362 18052 10364
rect 18076 10362 18132 10364
rect 18156 10362 18212 10364
rect 18236 10362 18292 10364
rect 18316 10362 18372 10364
rect 18396 10362 18452 10364
rect 18476 10362 18532 10364
rect 18556 10362 18612 10364
rect 18636 10362 18692 10364
rect 17516 10310 17554 10362
rect 17554 10310 17566 10362
rect 17566 10310 17572 10362
rect 17596 10310 17618 10362
rect 17618 10310 17630 10362
rect 17630 10310 17652 10362
rect 17676 10310 17682 10362
rect 17682 10310 17694 10362
rect 17694 10310 17732 10362
rect 17756 10310 17758 10362
rect 17758 10310 17810 10362
rect 17810 10310 17812 10362
rect 17836 10310 17874 10362
rect 17874 10310 17886 10362
rect 17886 10310 17892 10362
rect 17916 10310 17938 10362
rect 17938 10310 17950 10362
rect 17950 10310 17972 10362
rect 17996 10310 18002 10362
rect 18002 10310 18014 10362
rect 18014 10310 18052 10362
rect 18076 10310 18078 10362
rect 18078 10310 18130 10362
rect 18130 10310 18132 10362
rect 18156 10310 18194 10362
rect 18194 10310 18206 10362
rect 18206 10310 18212 10362
rect 18236 10310 18258 10362
rect 18258 10310 18270 10362
rect 18270 10310 18292 10362
rect 18316 10310 18322 10362
rect 18322 10310 18334 10362
rect 18334 10310 18372 10362
rect 18396 10310 18398 10362
rect 18398 10310 18450 10362
rect 18450 10310 18452 10362
rect 18476 10310 18514 10362
rect 18514 10310 18526 10362
rect 18526 10310 18532 10362
rect 18556 10310 18578 10362
rect 18578 10310 18590 10362
rect 18590 10310 18612 10362
rect 18636 10310 18642 10362
rect 18642 10310 18654 10362
rect 18654 10310 18692 10362
rect 17516 10308 17572 10310
rect 17596 10308 17652 10310
rect 17676 10308 17732 10310
rect 17756 10308 17812 10310
rect 17836 10308 17892 10310
rect 17916 10308 17972 10310
rect 17996 10308 18052 10310
rect 18076 10308 18132 10310
rect 18156 10308 18212 10310
rect 18236 10308 18292 10310
rect 18316 10308 18372 10310
rect 18396 10308 18452 10310
rect 18476 10308 18532 10310
rect 18556 10308 18612 10310
rect 18636 10308 18692 10310
rect 17958 9444 18014 9480
rect 17958 9424 17960 9444
rect 17960 9424 18012 9444
rect 18012 9424 18014 9444
rect 18878 10648 18934 10704
rect 18694 9424 18750 9480
rect 17516 9274 17572 9276
rect 17596 9274 17652 9276
rect 17676 9274 17732 9276
rect 17756 9274 17812 9276
rect 17836 9274 17892 9276
rect 17916 9274 17972 9276
rect 17996 9274 18052 9276
rect 18076 9274 18132 9276
rect 18156 9274 18212 9276
rect 18236 9274 18292 9276
rect 18316 9274 18372 9276
rect 18396 9274 18452 9276
rect 18476 9274 18532 9276
rect 18556 9274 18612 9276
rect 18636 9274 18692 9276
rect 17516 9222 17554 9274
rect 17554 9222 17566 9274
rect 17566 9222 17572 9274
rect 17596 9222 17618 9274
rect 17618 9222 17630 9274
rect 17630 9222 17652 9274
rect 17676 9222 17682 9274
rect 17682 9222 17694 9274
rect 17694 9222 17732 9274
rect 17756 9222 17758 9274
rect 17758 9222 17810 9274
rect 17810 9222 17812 9274
rect 17836 9222 17874 9274
rect 17874 9222 17886 9274
rect 17886 9222 17892 9274
rect 17916 9222 17938 9274
rect 17938 9222 17950 9274
rect 17950 9222 17972 9274
rect 17996 9222 18002 9274
rect 18002 9222 18014 9274
rect 18014 9222 18052 9274
rect 18076 9222 18078 9274
rect 18078 9222 18130 9274
rect 18130 9222 18132 9274
rect 18156 9222 18194 9274
rect 18194 9222 18206 9274
rect 18206 9222 18212 9274
rect 18236 9222 18258 9274
rect 18258 9222 18270 9274
rect 18270 9222 18292 9274
rect 18316 9222 18322 9274
rect 18322 9222 18334 9274
rect 18334 9222 18372 9274
rect 18396 9222 18398 9274
rect 18398 9222 18450 9274
rect 18450 9222 18452 9274
rect 18476 9222 18514 9274
rect 18514 9222 18526 9274
rect 18526 9222 18532 9274
rect 18556 9222 18578 9274
rect 18578 9222 18590 9274
rect 18590 9222 18612 9274
rect 18636 9222 18642 9274
rect 18642 9222 18654 9274
rect 18654 9222 18692 9274
rect 17516 9220 17572 9222
rect 17596 9220 17652 9222
rect 17676 9220 17732 9222
rect 17756 9220 17812 9222
rect 17836 9220 17892 9222
rect 17916 9220 17972 9222
rect 17996 9220 18052 9222
rect 18076 9220 18132 9222
rect 18156 9220 18212 9222
rect 18236 9220 18292 9222
rect 18316 9220 18372 9222
rect 18396 9220 18452 9222
rect 18476 9220 18532 9222
rect 18556 9220 18612 9222
rect 18636 9220 18692 9222
rect 16854 6024 16910 6080
rect 16670 3576 16726 3632
rect 18142 9016 18198 9072
rect 17516 8186 17572 8188
rect 17596 8186 17652 8188
rect 17676 8186 17732 8188
rect 17756 8186 17812 8188
rect 17836 8186 17892 8188
rect 17916 8186 17972 8188
rect 17996 8186 18052 8188
rect 18076 8186 18132 8188
rect 18156 8186 18212 8188
rect 18236 8186 18292 8188
rect 18316 8186 18372 8188
rect 18396 8186 18452 8188
rect 18476 8186 18532 8188
rect 18556 8186 18612 8188
rect 18636 8186 18692 8188
rect 17516 8134 17554 8186
rect 17554 8134 17566 8186
rect 17566 8134 17572 8186
rect 17596 8134 17618 8186
rect 17618 8134 17630 8186
rect 17630 8134 17652 8186
rect 17676 8134 17682 8186
rect 17682 8134 17694 8186
rect 17694 8134 17732 8186
rect 17756 8134 17758 8186
rect 17758 8134 17810 8186
rect 17810 8134 17812 8186
rect 17836 8134 17874 8186
rect 17874 8134 17886 8186
rect 17886 8134 17892 8186
rect 17916 8134 17938 8186
rect 17938 8134 17950 8186
rect 17950 8134 17972 8186
rect 17996 8134 18002 8186
rect 18002 8134 18014 8186
rect 18014 8134 18052 8186
rect 18076 8134 18078 8186
rect 18078 8134 18130 8186
rect 18130 8134 18132 8186
rect 18156 8134 18194 8186
rect 18194 8134 18206 8186
rect 18206 8134 18212 8186
rect 18236 8134 18258 8186
rect 18258 8134 18270 8186
rect 18270 8134 18292 8186
rect 18316 8134 18322 8186
rect 18322 8134 18334 8186
rect 18334 8134 18372 8186
rect 18396 8134 18398 8186
rect 18398 8134 18450 8186
rect 18450 8134 18452 8186
rect 18476 8134 18514 8186
rect 18514 8134 18526 8186
rect 18526 8134 18532 8186
rect 18556 8134 18578 8186
rect 18578 8134 18590 8186
rect 18590 8134 18612 8186
rect 18636 8134 18642 8186
rect 18642 8134 18654 8186
rect 18654 8134 18692 8186
rect 17516 8132 17572 8134
rect 17596 8132 17652 8134
rect 17676 8132 17732 8134
rect 17756 8132 17812 8134
rect 17836 8132 17892 8134
rect 17916 8132 17972 8134
rect 17996 8132 18052 8134
rect 18076 8132 18132 8134
rect 18156 8132 18212 8134
rect 18236 8132 18292 8134
rect 18316 8132 18372 8134
rect 18396 8132 18452 8134
rect 18476 8132 18532 8134
rect 18556 8132 18612 8134
rect 18636 8132 18692 8134
rect 17516 7098 17572 7100
rect 17596 7098 17652 7100
rect 17676 7098 17732 7100
rect 17756 7098 17812 7100
rect 17836 7098 17892 7100
rect 17916 7098 17972 7100
rect 17996 7098 18052 7100
rect 18076 7098 18132 7100
rect 18156 7098 18212 7100
rect 18236 7098 18292 7100
rect 18316 7098 18372 7100
rect 18396 7098 18452 7100
rect 18476 7098 18532 7100
rect 18556 7098 18612 7100
rect 18636 7098 18692 7100
rect 17516 7046 17554 7098
rect 17554 7046 17566 7098
rect 17566 7046 17572 7098
rect 17596 7046 17618 7098
rect 17618 7046 17630 7098
rect 17630 7046 17652 7098
rect 17676 7046 17682 7098
rect 17682 7046 17694 7098
rect 17694 7046 17732 7098
rect 17756 7046 17758 7098
rect 17758 7046 17810 7098
rect 17810 7046 17812 7098
rect 17836 7046 17874 7098
rect 17874 7046 17886 7098
rect 17886 7046 17892 7098
rect 17916 7046 17938 7098
rect 17938 7046 17950 7098
rect 17950 7046 17972 7098
rect 17996 7046 18002 7098
rect 18002 7046 18014 7098
rect 18014 7046 18052 7098
rect 18076 7046 18078 7098
rect 18078 7046 18130 7098
rect 18130 7046 18132 7098
rect 18156 7046 18194 7098
rect 18194 7046 18206 7098
rect 18206 7046 18212 7098
rect 18236 7046 18258 7098
rect 18258 7046 18270 7098
rect 18270 7046 18292 7098
rect 18316 7046 18322 7098
rect 18322 7046 18334 7098
rect 18334 7046 18372 7098
rect 18396 7046 18398 7098
rect 18398 7046 18450 7098
rect 18450 7046 18452 7098
rect 18476 7046 18514 7098
rect 18514 7046 18526 7098
rect 18526 7046 18532 7098
rect 18556 7046 18578 7098
rect 18578 7046 18590 7098
rect 18590 7046 18612 7098
rect 18636 7046 18642 7098
rect 18642 7046 18654 7098
rect 18654 7046 18692 7098
rect 17516 7044 17572 7046
rect 17596 7044 17652 7046
rect 17676 7044 17732 7046
rect 17756 7044 17812 7046
rect 17836 7044 17892 7046
rect 17916 7044 17972 7046
rect 17996 7044 18052 7046
rect 18076 7044 18132 7046
rect 18156 7044 18212 7046
rect 18236 7044 18292 7046
rect 18316 7044 18372 7046
rect 18396 7044 18452 7046
rect 18476 7044 18532 7046
rect 18556 7044 18612 7046
rect 18636 7044 18692 7046
rect 18786 6160 18842 6216
rect 17516 6010 17572 6012
rect 17596 6010 17652 6012
rect 17676 6010 17732 6012
rect 17756 6010 17812 6012
rect 17836 6010 17892 6012
rect 17916 6010 17972 6012
rect 17996 6010 18052 6012
rect 18076 6010 18132 6012
rect 18156 6010 18212 6012
rect 18236 6010 18292 6012
rect 18316 6010 18372 6012
rect 18396 6010 18452 6012
rect 18476 6010 18532 6012
rect 18556 6010 18612 6012
rect 18636 6010 18692 6012
rect 17516 5958 17554 6010
rect 17554 5958 17566 6010
rect 17566 5958 17572 6010
rect 17596 5958 17618 6010
rect 17618 5958 17630 6010
rect 17630 5958 17652 6010
rect 17676 5958 17682 6010
rect 17682 5958 17694 6010
rect 17694 5958 17732 6010
rect 17756 5958 17758 6010
rect 17758 5958 17810 6010
rect 17810 5958 17812 6010
rect 17836 5958 17874 6010
rect 17874 5958 17886 6010
rect 17886 5958 17892 6010
rect 17916 5958 17938 6010
rect 17938 5958 17950 6010
rect 17950 5958 17972 6010
rect 17996 5958 18002 6010
rect 18002 5958 18014 6010
rect 18014 5958 18052 6010
rect 18076 5958 18078 6010
rect 18078 5958 18130 6010
rect 18130 5958 18132 6010
rect 18156 5958 18194 6010
rect 18194 5958 18206 6010
rect 18206 5958 18212 6010
rect 18236 5958 18258 6010
rect 18258 5958 18270 6010
rect 18270 5958 18292 6010
rect 18316 5958 18322 6010
rect 18322 5958 18334 6010
rect 18334 5958 18372 6010
rect 18396 5958 18398 6010
rect 18398 5958 18450 6010
rect 18450 5958 18452 6010
rect 18476 5958 18514 6010
rect 18514 5958 18526 6010
rect 18526 5958 18532 6010
rect 18556 5958 18578 6010
rect 18578 5958 18590 6010
rect 18590 5958 18612 6010
rect 18636 5958 18642 6010
rect 18642 5958 18654 6010
rect 18654 5958 18692 6010
rect 17516 5956 17572 5958
rect 17596 5956 17652 5958
rect 17676 5956 17732 5958
rect 17756 5956 17812 5958
rect 17836 5956 17892 5958
rect 17916 5956 17972 5958
rect 17996 5956 18052 5958
rect 18076 5956 18132 5958
rect 18156 5956 18212 5958
rect 18236 5956 18292 5958
rect 18316 5956 18372 5958
rect 18396 5956 18452 5958
rect 18476 5956 18532 5958
rect 18556 5956 18612 5958
rect 18636 5956 18692 5958
rect 18050 5752 18106 5808
rect 17516 4922 17572 4924
rect 17596 4922 17652 4924
rect 17676 4922 17732 4924
rect 17756 4922 17812 4924
rect 17836 4922 17892 4924
rect 17916 4922 17972 4924
rect 17996 4922 18052 4924
rect 18076 4922 18132 4924
rect 18156 4922 18212 4924
rect 18236 4922 18292 4924
rect 18316 4922 18372 4924
rect 18396 4922 18452 4924
rect 18476 4922 18532 4924
rect 18556 4922 18612 4924
rect 18636 4922 18692 4924
rect 17516 4870 17554 4922
rect 17554 4870 17566 4922
rect 17566 4870 17572 4922
rect 17596 4870 17618 4922
rect 17618 4870 17630 4922
rect 17630 4870 17652 4922
rect 17676 4870 17682 4922
rect 17682 4870 17694 4922
rect 17694 4870 17732 4922
rect 17756 4870 17758 4922
rect 17758 4870 17810 4922
rect 17810 4870 17812 4922
rect 17836 4870 17874 4922
rect 17874 4870 17886 4922
rect 17886 4870 17892 4922
rect 17916 4870 17938 4922
rect 17938 4870 17950 4922
rect 17950 4870 17972 4922
rect 17996 4870 18002 4922
rect 18002 4870 18014 4922
rect 18014 4870 18052 4922
rect 18076 4870 18078 4922
rect 18078 4870 18130 4922
rect 18130 4870 18132 4922
rect 18156 4870 18194 4922
rect 18194 4870 18206 4922
rect 18206 4870 18212 4922
rect 18236 4870 18258 4922
rect 18258 4870 18270 4922
rect 18270 4870 18292 4922
rect 18316 4870 18322 4922
rect 18322 4870 18334 4922
rect 18334 4870 18372 4922
rect 18396 4870 18398 4922
rect 18398 4870 18450 4922
rect 18450 4870 18452 4922
rect 18476 4870 18514 4922
rect 18514 4870 18526 4922
rect 18526 4870 18532 4922
rect 18556 4870 18578 4922
rect 18578 4870 18590 4922
rect 18590 4870 18612 4922
rect 18636 4870 18642 4922
rect 18642 4870 18654 4922
rect 18654 4870 18692 4922
rect 17516 4868 17572 4870
rect 17596 4868 17652 4870
rect 17676 4868 17732 4870
rect 17756 4868 17812 4870
rect 17836 4868 17892 4870
rect 17916 4868 17972 4870
rect 17996 4868 18052 4870
rect 18076 4868 18132 4870
rect 18156 4868 18212 4870
rect 18236 4868 18292 4870
rect 18316 4868 18372 4870
rect 18396 4868 18452 4870
rect 18476 4868 18532 4870
rect 18556 4868 18612 4870
rect 18636 4868 18692 4870
rect 18694 3984 18750 4040
rect 17516 3834 17572 3836
rect 17596 3834 17652 3836
rect 17676 3834 17732 3836
rect 17756 3834 17812 3836
rect 17836 3834 17892 3836
rect 17916 3834 17972 3836
rect 17996 3834 18052 3836
rect 18076 3834 18132 3836
rect 18156 3834 18212 3836
rect 18236 3834 18292 3836
rect 18316 3834 18372 3836
rect 18396 3834 18452 3836
rect 18476 3834 18532 3836
rect 18556 3834 18612 3836
rect 18636 3834 18692 3836
rect 17516 3782 17554 3834
rect 17554 3782 17566 3834
rect 17566 3782 17572 3834
rect 17596 3782 17618 3834
rect 17618 3782 17630 3834
rect 17630 3782 17652 3834
rect 17676 3782 17682 3834
rect 17682 3782 17694 3834
rect 17694 3782 17732 3834
rect 17756 3782 17758 3834
rect 17758 3782 17810 3834
rect 17810 3782 17812 3834
rect 17836 3782 17874 3834
rect 17874 3782 17886 3834
rect 17886 3782 17892 3834
rect 17916 3782 17938 3834
rect 17938 3782 17950 3834
rect 17950 3782 17972 3834
rect 17996 3782 18002 3834
rect 18002 3782 18014 3834
rect 18014 3782 18052 3834
rect 18076 3782 18078 3834
rect 18078 3782 18130 3834
rect 18130 3782 18132 3834
rect 18156 3782 18194 3834
rect 18194 3782 18206 3834
rect 18206 3782 18212 3834
rect 18236 3782 18258 3834
rect 18258 3782 18270 3834
rect 18270 3782 18292 3834
rect 18316 3782 18322 3834
rect 18322 3782 18334 3834
rect 18334 3782 18372 3834
rect 18396 3782 18398 3834
rect 18398 3782 18450 3834
rect 18450 3782 18452 3834
rect 18476 3782 18514 3834
rect 18514 3782 18526 3834
rect 18526 3782 18532 3834
rect 18556 3782 18578 3834
rect 18578 3782 18590 3834
rect 18590 3782 18612 3834
rect 18636 3782 18642 3834
rect 18642 3782 18654 3834
rect 18654 3782 18692 3834
rect 17516 3780 17572 3782
rect 17596 3780 17652 3782
rect 17676 3780 17732 3782
rect 17756 3780 17812 3782
rect 17836 3780 17892 3782
rect 17916 3780 17972 3782
rect 17996 3780 18052 3782
rect 18076 3780 18132 3782
rect 18156 3780 18212 3782
rect 18236 3780 18292 3782
rect 18316 3780 18372 3782
rect 18396 3780 18452 3782
rect 18476 3780 18532 3782
rect 18556 3780 18612 3782
rect 18636 3780 18692 3782
rect 17038 3440 17094 3496
rect 16670 2760 16726 2816
rect 17516 2746 17572 2748
rect 17596 2746 17652 2748
rect 17676 2746 17732 2748
rect 17756 2746 17812 2748
rect 17836 2746 17892 2748
rect 17916 2746 17972 2748
rect 17996 2746 18052 2748
rect 18076 2746 18132 2748
rect 18156 2746 18212 2748
rect 18236 2746 18292 2748
rect 18316 2746 18372 2748
rect 18396 2746 18452 2748
rect 18476 2746 18532 2748
rect 18556 2746 18612 2748
rect 18636 2746 18692 2748
rect 17516 2694 17554 2746
rect 17554 2694 17566 2746
rect 17566 2694 17572 2746
rect 17596 2694 17618 2746
rect 17618 2694 17630 2746
rect 17630 2694 17652 2746
rect 17676 2694 17682 2746
rect 17682 2694 17694 2746
rect 17694 2694 17732 2746
rect 17756 2694 17758 2746
rect 17758 2694 17810 2746
rect 17810 2694 17812 2746
rect 17836 2694 17874 2746
rect 17874 2694 17886 2746
rect 17886 2694 17892 2746
rect 17916 2694 17938 2746
rect 17938 2694 17950 2746
rect 17950 2694 17972 2746
rect 17996 2694 18002 2746
rect 18002 2694 18014 2746
rect 18014 2694 18052 2746
rect 18076 2694 18078 2746
rect 18078 2694 18130 2746
rect 18130 2694 18132 2746
rect 18156 2694 18194 2746
rect 18194 2694 18206 2746
rect 18206 2694 18212 2746
rect 18236 2694 18258 2746
rect 18258 2694 18270 2746
rect 18270 2694 18292 2746
rect 18316 2694 18322 2746
rect 18322 2694 18334 2746
rect 18334 2694 18372 2746
rect 18396 2694 18398 2746
rect 18398 2694 18450 2746
rect 18450 2694 18452 2746
rect 18476 2694 18514 2746
rect 18514 2694 18526 2746
rect 18526 2694 18532 2746
rect 18556 2694 18578 2746
rect 18578 2694 18590 2746
rect 18590 2694 18612 2746
rect 18636 2694 18642 2746
rect 18642 2694 18654 2746
rect 18654 2694 18692 2746
rect 17516 2692 17572 2694
rect 17596 2692 17652 2694
rect 17676 2692 17732 2694
rect 17756 2692 17812 2694
rect 17836 2692 17892 2694
rect 17916 2692 17972 2694
rect 17996 2692 18052 2694
rect 18076 2692 18132 2694
rect 18156 2692 18212 2694
rect 18236 2692 18292 2694
rect 18316 2692 18372 2694
rect 18396 2692 18452 2694
rect 18476 2692 18532 2694
rect 18556 2692 18612 2694
rect 18636 2692 18692 2694
rect 19062 7520 19118 7576
rect 19062 5752 19118 5808
rect 18970 5208 19026 5264
rect 15842 1536 15898 1592
rect 15382 1284 15438 1320
rect 15382 1264 15384 1284
rect 15384 1264 15436 1284
rect 15436 1264 15438 1284
rect 18878 720 18934 776
rect 19154 5480 19210 5536
rect 19154 3984 19210 4040
rect 19062 992 19118 1048
rect 18970 448 19026 504
rect 19062 176 19118 232
rect 19430 13368 19486 13424
rect 19338 7520 19394 7576
rect 19706 5072 19762 5128
rect 19706 2896 19762 2952
rect 19798 2488 19854 2544
<< metal3 >>
rect 5506 17440 6702 17441
rect 5506 17376 5512 17440
rect 5576 17376 5592 17440
rect 5656 17376 5672 17440
rect 5736 17376 5752 17440
rect 5816 17376 5832 17440
rect 5896 17376 5912 17440
rect 5976 17376 5992 17440
rect 6056 17376 6072 17440
rect 6136 17376 6152 17440
rect 6216 17376 6232 17440
rect 6296 17376 6312 17440
rect 6376 17376 6392 17440
rect 6456 17376 6472 17440
rect 6536 17376 6552 17440
rect 6616 17376 6632 17440
rect 6696 17376 6702 17440
rect 5506 17375 6702 17376
rect 13506 17440 14702 17441
rect 13506 17376 13512 17440
rect 13576 17376 13592 17440
rect 13656 17376 13672 17440
rect 13736 17376 13752 17440
rect 13816 17376 13832 17440
rect 13896 17376 13912 17440
rect 13976 17376 13992 17440
rect 14056 17376 14072 17440
rect 14136 17376 14152 17440
rect 14216 17376 14232 17440
rect 14296 17376 14312 17440
rect 14376 17376 14392 17440
rect 14456 17376 14472 17440
rect 14536 17376 14552 17440
rect 14616 17376 14632 17440
rect 14696 17376 14702 17440
rect 13506 17375 14702 17376
rect 3325 17234 3391 17237
rect 10869 17234 10935 17237
rect 3325 17232 10935 17234
rect 3325 17176 3330 17232
rect 3386 17176 10874 17232
rect 10930 17176 10935 17232
rect 3325 17174 10935 17176
rect 3325 17171 3391 17174
rect 10869 17171 10935 17174
rect 1506 16896 2702 16897
rect 1506 16832 1512 16896
rect 1576 16832 1592 16896
rect 1656 16832 1672 16896
rect 1736 16832 1752 16896
rect 1816 16832 1832 16896
rect 1896 16832 1912 16896
rect 1976 16832 1992 16896
rect 2056 16832 2072 16896
rect 2136 16832 2152 16896
rect 2216 16832 2232 16896
rect 2296 16832 2312 16896
rect 2376 16832 2392 16896
rect 2456 16832 2472 16896
rect 2536 16832 2552 16896
rect 2616 16832 2632 16896
rect 2696 16832 2702 16896
rect 1506 16831 2702 16832
rect 9506 16896 10702 16897
rect 9506 16832 9512 16896
rect 9576 16832 9592 16896
rect 9656 16832 9672 16896
rect 9736 16832 9752 16896
rect 9816 16832 9832 16896
rect 9896 16832 9912 16896
rect 9976 16832 9992 16896
rect 10056 16832 10072 16896
rect 10136 16832 10152 16896
rect 10216 16832 10232 16896
rect 10296 16832 10312 16896
rect 10376 16832 10392 16896
rect 10456 16832 10472 16896
rect 10536 16832 10552 16896
rect 10616 16832 10632 16896
rect 10696 16832 10702 16896
rect 9506 16831 10702 16832
rect 17506 16896 18702 16897
rect 17506 16832 17512 16896
rect 17576 16832 17592 16896
rect 17656 16832 17672 16896
rect 17736 16832 17752 16896
rect 17816 16832 17832 16896
rect 17896 16832 17912 16896
rect 17976 16832 17992 16896
rect 18056 16832 18072 16896
rect 18136 16832 18152 16896
rect 18216 16832 18232 16896
rect 18296 16832 18312 16896
rect 18376 16832 18392 16896
rect 18456 16832 18472 16896
rect 18536 16832 18552 16896
rect 18616 16832 18632 16896
rect 18696 16832 18702 16896
rect 17506 16831 18702 16832
rect 5441 16690 5507 16693
rect 18781 16690 18847 16693
rect 5441 16688 18847 16690
rect 5441 16632 5446 16688
rect 5502 16632 18786 16688
rect 18842 16632 18847 16688
rect 5441 16630 18847 16632
rect 5441 16627 5507 16630
rect 18781 16627 18847 16630
rect 5506 16352 6702 16353
rect 5506 16288 5512 16352
rect 5576 16288 5592 16352
rect 5656 16288 5672 16352
rect 5736 16288 5752 16352
rect 5816 16288 5832 16352
rect 5896 16288 5912 16352
rect 5976 16288 5992 16352
rect 6056 16288 6072 16352
rect 6136 16288 6152 16352
rect 6216 16288 6232 16352
rect 6296 16288 6312 16352
rect 6376 16288 6392 16352
rect 6456 16288 6472 16352
rect 6536 16288 6552 16352
rect 6616 16288 6632 16352
rect 6696 16288 6702 16352
rect 5506 16287 6702 16288
rect 13506 16352 14702 16353
rect 13506 16288 13512 16352
rect 13576 16288 13592 16352
rect 13656 16288 13672 16352
rect 13736 16288 13752 16352
rect 13816 16288 13832 16352
rect 13896 16288 13912 16352
rect 13976 16288 13992 16352
rect 14056 16288 14072 16352
rect 14136 16288 14152 16352
rect 14216 16288 14232 16352
rect 14296 16288 14312 16352
rect 14376 16288 14392 16352
rect 14456 16288 14472 16352
rect 14536 16288 14552 16352
rect 14616 16288 14632 16352
rect 14696 16288 14702 16352
rect 13506 16287 14702 16288
rect 7649 16010 7715 16013
rect 16573 16010 16639 16013
rect 7649 16008 16639 16010
rect 7649 15952 7654 16008
rect 7710 15952 16578 16008
rect 16634 15952 16639 16008
rect 7649 15950 16639 15952
rect 7649 15947 7715 15950
rect 16573 15947 16639 15950
rect 1506 15808 2702 15809
rect 1506 15744 1512 15808
rect 1576 15744 1592 15808
rect 1656 15744 1672 15808
rect 1736 15744 1752 15808
rect 1816 15744 1832 15808
rect 1896 15744 1912 15808
rect 1976 15744 1992 15808
rect 2056 15744 2072 15808
rect 2136 15744 2152 15808
rect 2216 15744 2232 15808
rect 2296 15744 2312 15808
rect 2376 15744 2392 15808
rect 2456 15744 2472 15808
rect 2536 15744 2552 15808
rect 2616 15744 2632 15808
rect 2696 15744 2702 15808
rect 1506 15743 2702 15744
rect 9506 15808 10702 15809
rect 9506 15744 9512 15808
rect 9576 15744 9592 15808
rect 9656 15744 9672 15808
rect 9736 15744 9752 15808
rect 9816 15744 9832 15808
rect 9896 15744 9912 15808
rect 9976 15744 9992 15808
rect 10056 15744 10072 15808
rect 10136 15744 10152 15808
rect 10216 15744 10232 15808
rect 10296 15744 10312 15808
rect 10376 15744 10392 15808
rect 10456 15744 10472 15808
rect 10536 15744 10552 15808
rect 10616 15744 10632 15808
rect 10696 15744 10702 15808
rect 9506 15743 10702 15744
rect 17506 15808 18702 15809
rect 17506 15744 17512 15808
rect 17576 15744 17592 15808
rect 17656 15744 17672 15808
rect 17736 15744 17752 15808
rect 17816 15744 17832 15808
rect 17896 15744 17912 15808
rect 17976 15744 17992 15808
rect 18056 15744 18072 15808
rect 18136 15744 18152 15808
rect 18216 15744 18232 15808
rect 18296 15744 18312 15808
rect 18376 15744 18392 15808
rect 18456 15744 18472 15808
rect 18536 15744 18552 15808
rect 18616 15744 18632 15808
rect 18696 15744 18702 15808
rect 17506 15743 18702 15744
rect 6177 15738 6243 15741
rect 7189 15738 7255 15741
rect 6177 15736 7255 15738
rect 6177 15680 6182 15736
rect 6238 15680 7194 15736
rect 7250 15680 7255 15736
rect 6177 15678 7255 15680
rect 6177 15675 6243 15678
rect 7189 15675 7255 15678
rect 5441 15602 5507 15605
rect 11421 15602 11487 15605
rect 5441 15600 11487 15602
rect 5441 15544 5446 15600
rect 5502 15544 11426 15600
rect 11482 15544 11487 15600
rect 5441 15542 11487 15544
rect 5441 15539 5507 15542
rect 11421 15539 11487 15542
rect 5165 15466 5231 15469
rect 7741 15466 7807 15469
rect 5165 15464 7807 15466
rect 5165 15408 5170 15464
rect 5226 15408 7746 15464
rect 7802 15408 7807 15464
rect 5165 15406 7807 15408
rect 5165 15403 5231 15406
rect 7741 15403 7807 15406
rect 7465 15330 7531 15333
rect 11513 15330 11579 15333
rect 7465 15328 11579 15330
rect 7465 15272 7470 15328
rect 7526 15272 11518 15328
rect 11574 15272 11579 15328
rect 7465 15270 11579 15272
rect 7465 15267 7531 15270
rect 11513 15267 11579 15270
rect 5506 15264 6702 15265
rect 5506 15200 5512 15264
rect 5576 15200 5592 15264
rect 5656 15200 5672 15264
rect 5736 15200 5752 15264
rect 5816 15200 5832 15264
rect 5896 15200 5912 15264
rect 5976 15200 5992 15264
rect 6056 15200 6072 15264
rect 6136 15200 6152 15264
rect 6216 15200 6232 15264
rect 6296 15200 6312 15264
rect 6376 15200 6392 15264
rect 6456 15200 6472 15264
rect 6536 15200 6552 15264
rect 6616 15200 6632 15264
rect 6696 15200 6702 15264
rect 5506 15199 6702 15200
rect 13506 15264 14702 15265
rect 13506 15200 13512 15264
rect 13576 15200 13592 15264
rect 13656 15200 13672 15264
rect 13736 15200 13752 15264
rect 13816 15200 13832 15264
rect 13896 15200 13912 15264
rect 13976 15200 13992 15264
rect 14056 15200 14072 15264
rect 14136 15200 14152 15264
rect 14216 15200 14232 15264
rect 14296 15200 14312 15264
rect 14376 15200 14392 15264
rect 14456 15200 14472 15264
rect 14536 15200 14552 15264
rect 14616 15200 14632 15264
rect 14696 15200 14702 15264
rect 13506 15199 14702 15200
rect 7281 15194 7347 15197
rect 7238 15192 7347 15194
rect 7238 15136 7286 15192
rect 7342 15136 7347 15192
rect 7238 15131 7347 15136
rect 4981 15058 5047 15061
rect 5625 15058 5691 15061
rect 6545 15058 6611 15061
rect 4981 15056 6611 15058
rect 4981 15000 4986 15056
rect 5042 15000 5630 15056
rect 5686 15000 6550 15056
rect 6606 15000 6611 15056
rect 4981 14998 6611 15000
rect 4981 14995 5047 14998
rect 5625 14995 5691 14998
rect 6545 14995 6611 14998
rect 2773 14920 2839 14925
rect 2773 14864 2778 14920
rect 2834 14864 2839 14920
rect 2773 14859 2839 14864
rect 4889 14920 4955 14925
rect 7238 14922 7298 15131
rect 9397 14922 9463 14925
rect 11697 14922 11763 14925
rect 4889 14864 4894 14920
rect 4950 14864 4955 14920
rect 4889 14859 4955 14864
rect 5720 14862 7298 14922
rect 8250 14920 11763 14922
rect 8250 14864 9402 14920
rect 9458 14864 11702 14920
rect 11758 14864 11763 14920
rect 8250 14862 11763 14864
rect 1506 14720 2702 14721
rect 1506 14656 1512 14720
rect 1576 14656 1592 14720
rect 1656 14656 1672 14720
rect 1736 14656 1752 14720
rect 1816 14656 1832 14720
rect 1896 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2312 14720
rect 2376 14656 2392 14720
rect 2456 14656 2472 14720
rect 2536 14656 2552 14720
rect 2616 14656 2632 14720
rect 2696 14656 2702 14720
rect 1506 14655 2702 14656
rect 749 14514 815 14517
rect 246 14512 815 14514
rect 246 14456 754 14512
rect 810 14456 815 14512
rect 246 14454 815 14456
rect 105 12746 171 12749
rect 246 12746 306 14454
rect 749 14451 815 14454
rect 1577 14514 1643 14517
rect 2776 14514 2836 14859
rect 4892 14786 4952 14859
rect 5720 14789 5780 14862
rect 5717 14786 5783 14789
rect 4524 14784 5783 14786
rect 4524 14728 5722 14784
rect 5778 14728 5783 14784
rect 4524 14726 5783 14728
rect 4524 14517 4584 14726
rect 5717 14723 5783 14726
rect 6453 14786 6519 14789
rect 7373 14786 7439 14789
rect 8250 14786 8310 14862
rect 9397 14859 9463 14862
rect 11697 14859 11763 14862
rect 6453 14784 8310 14786
rect 6453 14728 6458 14784
rect 6514 14728 7378 14784
rect 7434 14728 8310 14784
rect 6453 14726 8310 14728
rect 6453 14723 6519 14726
rect 7373 14723 7439 14726
rect 9506 14720 10702 14721
rect 9506 14656 9512 14720
rect 9576 14656 9592 14720
rect 9656 14656 9672 14720
rect 9736 14656 9752 14720
rect 9816 14656 9832 14720
rect 9896 14656 9912 14720
rect 9976 14656 9992 14720
rect 10056 14656 10072 14720
rect 10136 14656 10152 14720
rect 10216 14656 10232 14720
rect 10296 14656 10312 14720
rect 10376 14656 10392 14720
rect 10456 14656 10472 14720
rect 10536 14656 10552 14720
rect 10616 14656 10632 14720
rect 10696 14656 10702 14720
rect 9506 14655 10702 14656
rect 17506 14720 18702 14721
rect 17506 14656 17512 14720
rect 17576 14656 17592 14720
rect 17656 14656 17672 14720
rect 17736 14656 17752 14720
rect 17816 14656 17832 14720
rect 17896 14656 17912 14720
rect 17976 14656 17992 14720
rect 18056 14656 18072 14720
rect 18136 14656 18152 14720
rect 18216 14656 18232 14720
rect 18296 14656 18312 14720
rect 18376 14656 18392 14720
rect 18456 14656 18472 14720
rect 18536 14656 18552 14720
rect 18616 14656 18632 14720
rect 18696 14656 18702 14720
rect 17506 14655 18702 14656
rect 5441 14650 5507 14653
rect 6637 14650 6703 14653
rect 4662 14648 6703 14650
rect 4662 14592 5446 14648
rect 5502 14592 6642 14648
rect 6698 14592 6703 14648
rect 4662 14590 6703 14592
rect 1577 14512 2836 14514
rect 1577 14456 1582 14512
rect 1638 14456 2836 14512
rect 1577 14454 2836 14456
rect 4521 14512 4587 14517
rect 4521 14456 4526 14512
rect 4582 14456 4587 14512
rect 1577 14451 1643 14454
rect 4521 14451 4587 14456
rect 565 14378 631 14381
rect 4662 14378 4722 14590
rect 5441 14587 5507 14590
rect 6637 14587 6703 14590
rect 5533 14514 5599 14517
rect 6269 14514 6335 14517
rect 6913 14514 6979 14517
rect 15745 14514 15811 14517
rect 5533 14512 5826 14514
rect 5533 14456 5538 14512
rect 5594 14456 5826 14512
rect 5533 14454 5826 14456
rect 5533 14451 5599 14454
rect 5625 14378 5691 14381
rect 565 14376 4722 14378
rect 565 14320 570 14376
rect 626 14320 4722 14376
rect 565 14318 4722 14320
rect 565 14315 631 14318
rect 4521 14242 4587 14245
rect 2960 14240 4587 14242
rect 2960 14184 4526 14240
rect 4582 14184 4587 14240
rect 2960 14182 4587 14184
rect 1853 13834 1919 13837
rect 1350 13832 1919 13834
rect 1350 13776 1858 13832
rect 1914 13776 1919 13832
rect 1350 13774 1919 13776
rect 1350 13426 1410 13774
rect 1853 13771 1919 13774
rect 2221 13834 2287 13837
rect 2221 13832 2836 13834
rect 2221 13776 2226 13832
rect 2282 13776 2836 13832
rect 2221 13774 2836 13776
rect 2221 13771 2287 13774
rect 1506 13632 2702 13633
rect 1506 13568 1512 13632
rect 1576 13568 1592 13632
rect 1656 13568 1672 13632
rect 1736 13568 1752 13632
rect 1816 13568 1832 13632
rect 1896 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2312 13632
rect 2376 13568 2392 13632
rect 2456 13568 2472 13632
rect 2536 13568 2552 13632
rect 2616 13568 2632 13632
rect 2696 13568 2702 13632
rect 1506 13567 2702 13568
rect 1761 13426 1827 13429
rect 1350 13424 1827 13426
rect 1350 13368 1766 13424
rect 1822 13368 1827 13424
rect 1350 13366 1827 13368
rect 1761 13363 1827 13366
rect 2313 13426 2379 13429
rect 2776 13426 2836 13774
rect 2960 13701 3020 14182
rect 4521 14179 4587 14182
rect 4521 14106 4587 14109
rect 4662 14106 4722 14318
rect 4521 14104 4722 14106
rect 4521 14048 4526 14104
rect 4582 14048 4722 14104
rect 4521 14046 4722 14048
rect 5214 14376 5691 14378
rect 5214 14320 5630 14376
rect 5686 14320 5691 14376
rect 5214 14318 5691 14320
rect 5766 14378 5826 14454
rect 6269 14512 15811 14514
rect 6269 14456 6274 14512
rect 6330 14456 6918 14512
rect 6974 14456 15750 14512
rect 15806 14456 15811 14512
rect 6269 14454 15811 14456
rect 6269 14451 6335 14454
rect 6913 14451 6979 14454
rect 15745 14451 15811 14454
rect 7649 14378 7715 14381
rect 5766 14376 7715 14378
rect 5766 14320 7654 14376
rect 7710 14320 7715 14376
rect 5766 14318 7715 14320
rect 4521 14043 4587 14046
rect 5073 13834 5139 13837
rect 5214 13834 5274 14318
rect 5625 14315 5691 14318
rect 7649 14315 7715 14318
rect 5506 14176 6702 14177
rect 5506 14112 5512 14176
rect 5576 14112 5592 14176
rect 5656 14112 5672 14176
rect 5736 14112 5752 14176
rect 5816 14112 5832 14176
rect 5896 14112 5912 14176
rect 5976 14112 5992 14176
rect 6056 14112 6072 14176
rect 6136 14112 6152 14176
rect 6216 14112 6232 14176
rect 6296 14112 6312 14176
rect 6376 14112 6392 14176
rect 6456 14112 6472 14176
rect 6536 14112 6552 14176
rect 6616 14112 6632 14176
rect 6696 14112 6702 14176
rect 5506 14111 6702 14112
rect 13506 14176 14702 14177
rect 13506 14112 13512 14176
rect 13576 14112 13592 14176
rect 13656 14112 13672 14176
rect 13736 14112 13752 14176
rect 13816 14112 13832 14176
rect 13896 14112 13912 14176
rect 13976 14112 13992 14176
rect 14056 14112 14072 14176
rect 14136 14112 14152 14176
rect 14216 14112 14232 14176
rect 14296 14112 14312 14176
rect 14376 14112 14392 14176
rect 14456 14112 14472 14176
rect 14536 14112 14552 14176
rect 14616 14112 14632 14176
rect 14696 14112 14702 14176
rect 13506 14111 14702 14112
rect 9029 14106 9095 14109
rect 10317 14106 10383 14109
rect 9029 14104 10383 14106
rect 9029 14048 9034 14104
rect 9090 14048 10322 14104
rect 10378 14048 10383 14104
rect 9029 14046 10383 14048
rect 9029 14043 9095 14046
rect 10317 14043 10383 14046
rect 8201 13834 8267 13837
rect 5073 13832 5274 13834
rect 5073 13776 5078 13832
rect 5134 13776 5274 13832
rect 5073 13774 5274 13776
rect 5720 13832 8267 13834
rect 5720 13776 8206 13832
rect 8262 13776 8267 13832
rect 5720 13774 8267 13776
rect 5073 13771 5139 13774
rect 2957 13696 3023 13701
rect 2957 13640 2962 13696
rect 3018 13640 3023 13696
rect 2957 13635 3023 13640
rect 4429 13562 4495 13565
rect 5533 13562 5599 13565
rect 2313 13424 2836 13426
rect 2313 13368 2318 13424
rect 2374 13368 2836 13424
rect 2313 13366 2836 13368
rect 3788 13560 5599 13562
rect 3788 13504 4434 13560
rect 4490 13504 5538 13560
rect 5594 13504 5599 13560
rect 3788 13502 5599 13504
rect 2313 13363 2379 13366
rect 1945 13290 2011 13293
rect 3788 13290 3848 13502
rect 4429 13499 4495 13502
rect 5533 13499 5599 13502
rect 4153 13426 4219 13429
rect 5720 13426 5780 13774
rect 8201 13771 8267 13774
rect 6821 13698 6887 13701
rect 6821 13696 8402 13698
rect 6821 13640 6826 13696
rect 6882 13640 8402 13696
rect 6821 13638 8402 13640
rect 6821 13635 6887 13638
rect 5901 13562 5967 13565
rect 5901 13560 7666 13562
rect 5901 13504 5906 13560
rect 5962 13504 7666 13560
rect 5901 13502 7666 13504
rect 5901 13499 5967 13502
rect 1945 13288 3848 13290
rect 1945 13232 1950 13288
rect 2006 13232 3848 13288
rect 1945 13230 3848 13232
rect 3926 13424 4219 13426
rect 3926 13368 4158 13424
rect 4214 13368 4219 13424
rect 3926 13366 4219 13368
rect 1945 13227 2011 13230
rect 657 13154 723 13157
rect 3509 13154 3575 13157
rect 657 13152 3575 13154
rect 657 13096 662 13152
rect 718 13096 3514 13152
rect 3570 13096 3575 13152
rect 657 13094 3575 13096
rect 657 13091 723 13094
rect 3509 13091 3575 13094
rect 3926 13018 3986 13366
rect 4153 13363 4219 13366
rect 4294 13366 5780 13426
rect 4294 13293 4354 13366
rect 4245 13288 4354 13293
rect 4245 13232 4250 13288
rect 4306 13232 4354 13288
rect 4245 13230 4354 13232
rect 5165 13288 5231 13293
rect 5717 13290 5783 13293
rect 5165 13232 5170 13288
rect 5226 13232 5231 13288
rect 4245 13227 4311 13230
rect 5165 13227 5231 13232
rect 5352 13288 5783 13290
rect 5352 13232 5722 13288
rect 5778 13232 5783 13288
rect 5352 13230 5783 13232
rect 5168 13021 5228 13227
rect 3006 12958 3986 13018
rect 4061 13016 4127 13021
rect 4981 13018 5047 13021
rect 4061 12960 4066 13016
rect 4122 12960 4127 13016
rect 2313 12882 2379 12885
rect 105 12744 306 12746
rect 105 12688 110 12744
rect 166 12688 306 12744
rect 105 12686 306 12688
rect 1166 12880 2379 12882
rect 1166 12824 2318 12880
rect 2374 12824 2379 12880
rect 1166 12822 2379 12824
rect 105 12683 171 12686
rect 1166 12202 1226 12822
rect 2313 12819 2379 12822
rect 2865 12880 2931 12885
rect 2865 12824 2870 12880
rect 2926 12824 2931 12880
rect 2865 12819 2931 12824
rect 2681 12746 2747 12749
rect 1350 12744 2747 12746
rect 1350 12688 2686 12744
rect 2742 12688 2747 12744
rect 1350 12686 2747 12688
rect 1350 12338 1410 12686
rect 2681 12683 2747 12686
rect 1506 12544 2702 12545
rect 1506 12480 1512 12544
rect 1576 12480 1592 12544
rect 1656 12480 1672 12544
rect 1736 12480 1752 12544
rect 1816 12480 1832 12544
rect 1896 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2312 12544
rect 2376 12480 2392 12544
rect 2456 12480 2472 12544
rect 2536 12480 2552 12544
rect 2616 12480 2632 12544
rect 2696 12480 2702 12544
rect 1506 12479 2702 12480
rect 2868 12341 2928 12819
rect 2313 12338 2379 12341
rect 1350 12336 2379 12338
rect 1350 12280 2318 12336
rect 2374 12280 2379 12336
rect 1350 12278 2379 12280
rect 2313 12275 2379 12278
rect 2865 12336 2931 12341
rect 2865 12280 2870 12336
rect 2926 12280 2931 12336
rect 2865 12275 2931 12280
rect 2221 12202 2287 12205
rect 1166 12200 2287 12202
rect 1166 12144 2226 12200
rect 2282 12144 2287 12200
rect 1166 12142 2287 12144
rect 2221 12139 2287 12142
rect 3006 11930 3066 12958
rect 4061 12955 4127 12960
rect 4248 13016 5047 13018
rect 4248 12960 4986 13016
rect 5042 12960 5047 13016
rect 4248 12958 5047 12960
rect 4064 12610 4124 12955
rect 3144 12550 4124 12610
rect 3144 12477 3204 12550
rect 3141 12472 3207 12477
rect 3877 12474 3943 12477
rect 3141 12416 3146 12472
rect 3202 12416 3207 12472
rect 3141 12411 3207 12416
rect 3558 12472 3943 12474
rect 3558 12416 3882 12472
rect 3938 12416 3943 12472
rect 3558 12414 3943 12416
rect 3558 12338 3618 12414
rect 3877 12411 3943 12414
rect 4248 12338 4308 12958
rect 4981 12955 5047 12958
rect 5165 13016 5231 13021
rect 5165 12960 5170 13016
rect 5226 12960 5231 13016
rect 5165 12955 5231 12960
rect 5352 12916 5412 13230
rect 5717 13227 5783 13230
rect 6637 13290 6703 13293
rect 6637 13288 6884 13290
rect 6637 13232 6642 13288
rect 6698 13232 6884 13288
rect 6637 13230 6884 13232
rect 6637 13227 6703 13230
rect 5506 13088 6702 13089
rect 5506 13024 5512 13088
rect 5576 13024 5592 13088
rect 5656 13024 5672 13088
rect 5736 13024 5752 13088
rect 5816 13024 5832 13088
rect 5896 13024 5912 13088
rect 5976 13024 5992 13088
rect 6056 13024 6072 13088
rect 6136 13024 6152 13088
rect 6216 13024 6232 13088
rect 6296 13024 6312 13088
rect 6376 13024 6392 13088
rect 6456 13024 6472 13088
rect 6536 13024 6552 13088
rect 6616 13024 6632 13088
rect 6696 13024 6702 13088
rect 5506 13023 6702 13024
rect 4889 12880 4955 12885
rect 4889 12824 4894 12880
rect 4950 12824 4955 12880
rect 5352 12882 5504 12916
rect 5809 12882 5875 12885
rect 5352 12880 5875 12882
rect 5352 12856 5814 12880
rect 4889 12819 4955 12824
rect 5444 12824 5814 12856
rect 5870 12824 5875 12880
rect 5444 12822 5875 12824
rect 5809 12819 5875 12822
rect 6545 12882 6611 12885
rect 6824 12882 6884 13230
rect 7373 13288 7439 13293
rect 7373 13232 7378 13288
rect 7434 13232 7439 13288
rect 7373 13227 7439 13232
rect 7189 13016 7255 13021
rect 7189 12960 7194 13016
rect 7250 12960 7255 13016
rect 7189 12955 7255 12960
rect 6545 12880 6884 12882
rect 6545 12824 6550 12880
rect 6606 12824 6884 12880
rect 6545 12822 6884 12824
rect 6545 12819 6611 12822
rect 4892 12746 4952 12819
rect 5717 12746 5783 12749
rect 4892 12744 5783 12746
rect 4892 12688 5722 12744
rect 5778 12688 5783 12744
rect 4892 12686 5783 12688
rect 5717 12683 5783 12686
rect 6821 12746 6887 12749
rect 7192 12746 7252 12955
rect 6821 12744 7252 12746
rect 6821 12688 6826 12744
rect 6882 12688 7252 12744
rect 6821 12686 7252 12688
rect 6821 12683 6887 12686
rect 4889 12474 4955 12477
rect 5993 12474 6059 12477
rect 4889 12472 6059 12474
rect 4889 12416 4894 12472
rect 4950 12416 5998 12472
rect 6054 12416 6059 12472
rect 4889 12414 6059 12416
rect 7376 12474 7436 13227
rect 7606 13157 7666 13502
rect 8017 13560 8083 13565
rect 8017 13504 8022 13560
rect 8078 13504 8083 13560
rect 8017 13499 8083 13504
rect 8342 13562 8402 13638
rect 9506 13632 10702 13633
rect 9506 13568 9512 13632
rect 9576 13568 9592 13632
rect 9656 13568 9672 13632
rect 9736 13568 9752 13632
rect 9816 13568 9832 13632
rect 9896 13568 9912 13632
rect 9976 13568 9992 13632
rect 10056 13568 10072 13632
rect 10136 13568 10152 13632
rect 10216 13568 10232 13632
rect 10296 13568 10312 13632
rect 10376 13568 10392 13632
rect 10456 13568 10472 13632
rect 10536 13568 10552 13632
rect 10616 13568 10632 13632
rect 10696 13568 10702 13632
rect 9506 13567 10702 13568
rect 17506 13632 18702 13633
rect 17506 13568 17512 13632
rect 17576 13568 17592 13632
rect 17656 13568 17672 13632
rect 17736 13568 17752 13632
rect 17816 13568 17832 13632
rect 17896 13568 17912 13632
rect 17976 13568 17992 13632
rect 18056 13568 18072 13632
rect 18136 13568 18152 13632
rect 18216 13568 18232 13632
rect 18296 13568 18312 13632
rect 18376 13568 18392 13632
rect 18456 13568 18472 13632
rect 18536 13568 18552 13632
rect 18616 13568 18632 13632
rect 18696 13568 18702 13632
rect 17506 13567 18702 13568
rect 8753 13562 8819 13565
rect 8342 13560 8819 13562
rect 8342 13504 8758 13560
rect 8814 13504 8819 13560
rect 8342 13502 8819 13504
rect 8753 13499 8819 13502
rect 7557 13152 7666 13157
rect 7557 13096 7562 13152
rect 7618 13096 7666 13152
rect 7557 13094 7666 13096
rect 7557 13091 7623 13094
rect 8020 13018 8080 13499
rect 19425 13426 19491 13429
rect 9630 13424 19491 13426
rect 9630 13368 19430 13424
rect 19486 13368 19491 13424
rect 9630 13366 19491 13368
rect 8201 13288 8267 13293
rect 8201 13232 8206 13288
rect 8262 13232 8267 13288
rect 8201 13227 8267 13232
rect 8204 13154 8264 13227
rect 9630 13154 9690 13366
rect 19425 13363 19491 13366
rect 10777 13288 10843 13293
rect 10777 13232 10782 13288
rect 10838 13232 10843 13288
rect 10777 13227 10843 13232
rect 8204 13094 9690 13154
rect 10780 13154 10840 13227
rect 10780 13094 11484 13154
rect 8020 12958 8310 13018
rect 8109 12744 8175 12749
rect 8109 12688 8114 12744
rect 8170 12688 8175 12744
rect 8109 12683 8175 12688
rect 7376 12414 7988 12474
rect 4889 12411 4955 12414
rect 5993 12411 6059 12414
rect 3144 12278 3618 12338
rect 3742 12278 4308 12338
rect 4429 12338 4495 12341
rect 5257 12338 5323 12341
rect 4429 12336 5323 12338
rect 4429 12280 4434 12336
rect 4490 12280 5262 12336
rect 5318 12280 5323 12336
rect 4429 12278 5323 12280
rect 3144 12069 3204 12278
rect 3742 12202 3802 12278
rect 4429 12275 4495 12278
rect 5257 12275 5323 12278
rect 5441 12338 5507 12341
rect 5625 12338 5691 12341
rect 5441 12336 5691 12338
rect 5441 12280 5446 12336
rect 5502 12280 5630 12336
rect 5686 12280 5691 12336
rect 5441 12278 5691 12280
rect 5441 12275 5507 12278
rect 5625 12275 5691 12278
rect 6177 12338 6243 12341
rect 6913 12338 6979 12341
rect 7741 12338 7807 12341
rect 6177 12336 6979 12338
rect 6177 12280 6182 12336
rect 6238 12280 6918 12336
rect 6974 12280 6979 12336
rect 6177 12278 6979 12280
rect 6177 12275 6243 12278
rect 6913 12275 6979 12278
rect 7054 12336 7807 12338
rect 7054 12280 7746 12336
rect 7802 12280 7807 12336
rect 7054 12278 7807 12280
rect 6453 12202 6519 12205
rect 3558 12142 3802 12202
rect 4110 12200 6519 12202
rect 4110 12144 6458 12200
rect 6514 12144 6519 12200
rect 4110 12142 6519 12144
rect 3141 12064 3207 12069
rect 3141 12008 3146 12064
rect 3202 12008 3207 12064
rect 3141 12003 3207 12008
rect 3417 11930 3483 11933
rect 3006 11928 3483 11930
rect 3006 11872 3422 11928
rect 3478 11872 3483 11928
rect 3006 11870 3483 11872
rect 3417 11867 3483 11870
rect 2589 11794 2655 11797
rect 3558 11794 3618 12142
rect 4110 11930 4170 12142
rect 6453 12139 6519 12142
rect 6637 12202 6703 12205
rect 6637 12200 6884 12202
rect 6637 12144 6642 12200
rect 6698 12144 6884 12200
rect 6637 12142 6884 12144
rect 6637 12139 6703 12142
rect 5506 12000 6702 12001
rect 5506 11936 5512 12000
rect 5576 11936 5592 12000
rect 5656 11936 5672 12000
rect 5736 11936 5752 12000
rect 5816 11936 5832 12000
rect 5896 11936 5912 12000
rect 5976 11936 5992 12000
rect 6056 11936 6072 12000
rect 6136 11936 6152 12000
rect 6216 11936 6232 12000
rect 6296 11936 6312 12000
rect 6376 11936 6392 12000
rect 6456 11936 6472 12000
rect 6536 11936 6552 12000
rect 6616 11936 6632 12000
rect 6696 11936 6702 12000
rect 5506 11935 6702 11936
rect 3972 11870 4170 11930
rect 6824 11930 6884 12142
rect 7054 12069 7114 12278
rect 7741 12275 7807 12278
rect 7928 12205 7988 12414
rect 8112 12338 8172 12683
rect 8250 12610 8310 12958
rect 10869 12882 10935 12885
rect 10869 12880 10978 12882
rect 10869 12824 10874 12880
rect 10930 12824 10978 12880
rect 10869 12819 10978 12824
rect 8661 12746 8727 12749
rect 9397 12746 9463 12749
rect 8661 12744 9463 12746
rect 8661 12688 8666 12744
rect 8722 12688 9402 12744
rect 9458 12688 9463 12744
rect 8661 12686 9463 12688
rect 8661 12683 8727 12686
rect 9397 12683 9463 12686
rect 10133 12746 10199 12749
rect 10133 12744 10840 12746
rect 10133 12688 10138 12744
rect 10194 12688 10840 12744
rect 10133 12686 10840 12688
rect 10133 12683 10199 12686
rect 8250 12550 9092 12610
rect 8661 12338 8727 12341
rect 8112 12336 8727 12338
rect 8112 12280 8666 12336
rect 8722 12280 8727 12336
rect 8112 12278 8727 12280
rect 8661 12275 8727 12278
rect 9032 12205 9092 12550
rect 9506 12544 10702 12545
rect 9506 12480 9512 12544
rect 9576 12480 9592 12544
rect 9656 12480 9672 12544
rect 9736 12480 9752 12544
rect 9816 12480 9832 12544
rect 9896 12480 9912 12544
rect 9976 12480 9992 12544
rect 10056 12480 10072 12544
rect 10136 12480 10152 12544
rect 10216 12480 10232 12544
rect 10296 12480 10312 12544
rect 10376 12480 10392 12544
rect 10456 12480 10472 12544
rect 10536 12480 10552 12544
rect 10616 12480 10632 12544
rect 10696 12480 10702 12544
rect 9506 12479 10702 12480
rect 10780 12372 10840 12686
rect 10734 12341 10840 12372
rect 9397 12338 9463 12341
rect 10317 12338 10383 12341
rect 9397 12336 10383 12338
rect 9397 12280 9402 12336
rect 9458 12280 10322 12336
rect 10378 12280 10383 12336
rect 9397 12278 10383 12280
rect 9397 12275 9463 12278
rect 10317 12275 10383 12278
rect 10685 12336 10840 12341
rect 10685 12280 10690 12336
rect 10746 12312 10840 12336
rect 10746 12280 10794 12312
rect 10685 12278 10794 12280
rect 10685 12275 10751 12278
rect 7281 12200 7347 12205
rect 7281 12144 7286 12200
rect 7342 12144 7347 12200
rect 7281 12139 7347 12144
rect 7925 12200 7991 12205
rect 7925 12144 7930 12200
rect 7986 12144 7991 12200
rect 7925 12139 7991 12144
rect 9029 12200 9095 12205
rect 9029 12144 9034 12200
rect 9090 12144 9095 12200
rect 9029 12139 9095 12144
rect 9765 12202 9831 12205
rect 10777 12202 10843 12205
rect 9765 12200 10843 12202
rect 9765 12144 9770 12200
rect 9826 12144 10782 12200
rect 10838 12144 10843 12200
rect 9765 12142 10843 12144
rect 9765 12139 9831 12142
rect 10777 12139 10843 12142
rect 7005 12064 7114 12069
rect 7005 12008 7010 12064
rect 7066 12008 7114 12064
rect 7005 12006 7114 12008
rect 7005 12003 7071 12006
rect 6824 11870 7068 11930
rect 3785 11794 3851 11797
rect 2589 11792 3020 11794
rect 2589 11736 2594 11792
rect 2650 11736 3020 11792
rect 2589 11734 3020 11736
rect 3558 11792 3851 11794
rect 3558 11736 3790 11792
rect 3846 11736 3851 11792
rect 3558 11734 3851 11736
rect 2589 11731 2655 11734
rect 2405 11658 2471 11661
rect 2405 11656 2836 11658
rect 2405 11600 2410 11656
rect 2466 11600 2836 11656
rect 2405 11598 2836 11600
rect 2405 11595 2471 11598
rect 1506 11456 2702 11457
rect 1506 11392 1512 11456
rect 1576 11392 1592 11456
rect 1656 11392 1672 11456
rect 1736 11392 1752 11456
rect 1816 11392 1832 11456
rect 1896 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2312 11456
rect 2376 11392 2392 11456
rect 2456 11392 2472 11456
rect 2536 11392 2552 11456
rect 2616 11392 2632 11456
rect 2696 11392 2702 11456
rect 1506 11391 2702 11392
rect 2776 11386 2836 11598
rect 2960 11522 3020 11734
rect 3785 11731 3851 11734
rect 3141 11658 3207 11661
rect 3972 11658 4032 11870
rect 5625 11794 5691 11797
rect 6821 11794 6887 11797
rect 3141 11656 4032 11658
rect 3141 11600 3146 11656
rect 3202 11600 4032 11656
rect 3141 11598 4032 11600
rect 4110 11734 4538 11794
rect 3141 11595 3207 11598
rect 4110 11522 4170 11734
rect 2960 11462 4170 11522
rect 4478 11522 4538 11734
rect 5625 11792 6887 11794
rect 5625 11736 5630 11792
rect 5686 11736 6826 11792
rect 6882 11736 6887 11792
rect 5625 11734 6887 11736
rect 5625 11731 5691 11734
rect 6821 11731 6887 11734
rect 5257 11658 5323 11661
rect 7008 11658 7068 11870
rect 5257 11656 7068 11658
rect 5257 11600 5262 11656
rect 5318 11600 7068 11656
rect 5257 11598 7068 11600
rect 5257 11595 5323 11598
rect 4889 11522 4955 11525
rect 5809 11522 5875 11525
rect 4478 11520 5875 11522
rect 4478 11464 4894 11520
rect 4950 11464 5814 11520
rect 5870 11464 5875 11520
rect 4478 11462 5875 11464
rect 4889 11459 4955 11462
rect 5809 11459 5875 11462
rect 6545 11522 6611 11525
rect 7284 11522 7344 12139
rect 10918 12066 10978 12819
rect 11145 12610 11211 12613
rect 11102 12608 11211 12610
rect 11102 12552 11150 12608
rect 11206 12552 11211 12608
rect 11102 12547 11211 12552
rect 11102 12069 11162 12547
rect 6545 11520 7344 11522
rect 6545 11464 6550 11520
rect 6606 11464 7344 11520
rect 6545 11462 7344 11464
rect 7468 12006 10978 12066
rect 11053 12064 11162 12069
rect 11053 12008 11058 12064
rect 11114 12008 11162 12064
rect 11053 12006 11162 12008
rect 6545 11459 6611 11462
rect 5993 11386 6059 11389
rect 2776 11384 6059 11386
rect 2776 11328 5998 11384
rect 6054 11328 6059 11384
rect 2776 11326 6059 11328
rect 5993 11323 6059 11326
rect 7468 11250 7528 12006
rect 11053 12003 11119 12006
rect 7649 11930 7715 11933
rect 7649 11928 7896 11930
rect 7649 11872 7654 11928
rect 7710 11872 7896 11928
rect 7649 11870 7896 11872
rect 7649 11867 7715 11870
rect 7649 11656 7715 11661
rect 7649 11600 7654 11656
rect 7710 11600 7715 11656
rect 7649 11595 7715 11600
rect 752 11190 7528 11250
rect 752 11117 812 11190
rect 749 11112 815 11117
rect 749 11056 754 11112
rect 810 11056 815 11112
rect 749 11051 815 11056
rect 3969 11114 4035 11117
rect 7652 11114 7712 11595
rect 3969 11112 7712 11114
rect 3969 11056 3974 11112
rect 4030 11056 7712 11112
rect 3969 11054 7712 11056
rect 3969 11051 4035 11054
rect 1853 10978 1919 10981
rect 4613 10978 4679 10981
rect 1853 10976 4679 10978
rect 1853 10920 1858 10976
rect 1914 10920 4618 10976
rect 4674 10920 4679 10976
rect 1853 10918 4679 10920
rect 1853 10915 1919 10918
rect 4613 10915 4679 10918
rect 7281 10976 7347 10981
rect 7281 10920 7286 10976
rect 7342 10920 7347 10976
rect 7281 10915 7347 10920
rect 5506 10912 6702 10913
rect 5506 10848 5512 10912
rect 5576 10848 5592 10912
rect 5656 10848 5672 10912
rect 5736 10848 5752 10912
rect 5816 10848 5832 10912
rect 5896 10848 5912 10912
rect 5976 10848 5992 10912
rect 6056 10848 6072 10912
rect 6136 10848 6152 10912
rect 6216 10848 6232 10912
rect 6296 10848 6312 10912
rect 6376 10848 6392 10912
rect 6456 10848 6472 10912
rect 6536 10848 6552 10912
rect 6616 10848 6632 10912
rect 6696 10848 6702 10912
rect 5506 10847 6702 10848
rect 4153 10842 4219 10845
rect 4337 10842 4403 10845
rect 4153 10840 4403 10842
rect 4153 10784 4158 10840
rect 4214 10784 4342 10840
rect 4398 10784 4403 10840
rect 4153 10782 4403 10784
rect 4153 10779 4219 10782
rect 4337 10779 4403 10782
rect 5257 10706 5323 10709
rect 5257 10704 5780 10706
rect 5257 10648 5262 10704
rect 5318 10648 5780 10704
rect 5257 10646 5780 10648
rect 5257 10643 5323 10646
rect 4061 10570 4127 10573
rect 5533 10570 5599 10573
rect 4061 10568 5599 10570
rect 4061 10512 4066 10568
rect 4122 10512 5538 10568
rect 5594 10512 5599 10568
rect 4061 10510 5599 10512
rect 4061 10507 4127 10510
rect 5533 10507 5599 10510
rect 5720 10434 5780 10646
rect 7284 10570 7344 10915
rect 7652 10706 7712 11054
rect 7836 10981 7896 11870
rect 8109 11928 8175 11933
rect 9121 11930 9187 11933
rect 8109 11872 8114 11928
rect 8170 11872 8175 11928
rect 8109 11867 8175 11872
rect 8756 11928 9187 11930
rect 8756 11872 9126 11928
rect 9182 11872 9187 11928
rect 8756 11870 9187 11872
rect 8112 11386 8172 11867
rect 8477 11658 8543 11661
rect 7974 11326 8172 11386
rect 8250 11656 8543 11658
rect 8250 11600 8482 11656
rect 8538 11600 8543 11656
rect 8250 11598 8543 11600
rect 7974 10981 8034 11326
rect 8250 11253 8310 11598
rect 8477 11595 8543 11598
rect 8385 11386 8451 11389
rect 8756 11386 8816 11870
rect 9121 11867 9187 11870
rect 9305 11930 9371 11933
rect 9305 11928 10978 11930
rect 9305 11872 9310 11928
rect 9366 11872 10978 11928
rect 9305 11870 10978 11872
rect 9305 11867 9371 11870
rect 9213 11794 9279 11797
rect 9078 11792 9279 11794
rect 9078 11736 9218 11792
rect 9274 11736 9279 11792
rect 9078 11734 9279 11736
rect 8937 11522 9003 11525
rect 8385 11384 8816 11386
rect 8385 11328 8390 11384
rect 8446 11328 8816 11384
rect 8385 11326 8816 11328
rect 8894 11520 9003 11522
rect 8894 11464 8942 11520
rect 8998 11464 9003 11520
rect 8894 11459 9003 11464
rect 8385 11323 8451 11326
rect 8201 11248 8310 11253
rect 8201 11192 8206 11248
rect 8262 11192 8310 11248
rect 8201 11190 8310 11192
rect 8569 11250 8635 11253
rect 8894 11250 8954 11459
rect 9078 11389 9138 11734
rect 9213 11731 9279 11734
rect 9397 11794 9463 11797
rect 9857 11794 9923 11797
rect 10777 11794 10843 11797
rect 9397 11792 10843 11794
rect 9397 11736 9402 11792
rect 9458 11736 9862 11792
rect 9918 11736 10782 11792
rect 10838 11736 10843 11792
rect 9397 11734 10843 11736
rect 9397 11731 9463 11734
rect 9857 11731 9923 11734
rect 10777 11731 10843 11734
rect 10041 11658 10107 11661
rect 9029 11384 9138 11389
rect 9029 11328 9034 11384
rect 9090 11328 9138 11384
rect 9029 11326 9138 11328
rect 9262 11656 10107 11658
rect 9262 11600 10046 11656
rect 10102 11600 10107 11656
rect 9262 11598 10107 11600
rect 9029 11323 9095 11326
rect 8569 11248 8954 11250
rect 8569 11192 8574 11248
rect 8630 11192 8954 11248
rect 8569 11190 8954 11192
rect 9262 11250 9322 11598
rect 10041 11595 10107 11598
rect 10225 11658 10291 11661
rect 10225 11656 10840 11658
rect 10225 11600 10230 11656
rect 10286 11600 10840 11656
rect 10225 11598 10840 11600
rect 10225 11595 10291 11598
rect 9506 11456 10702 11457
rect 9506 11392 9512 11456
rect 9576 11392 9592 11456
rect 9656 11392 9672 11456
rect 9736 11392 9752 11456
rect 9816 11392 9832 11456
rect 9896 11392 9912 11456
rect 9976 11392 9992 11456
rect 10056 11392 10072 11456
rect 10136 11392 10152 11456
rect 10216 11392 10232 11456
rect 10296 11392 10312 11456
rect 10376 11392 10392 11456
rect 10456 11392 10472 11456
rect 10536 11392 10552 11456
rect 10616 11392 10632 11456
rect 10696 11392 10702 11456
rect 9506 11391 10702 11392
rect 9949 11250 10015 11253
rect 9262 11248 10015 11250
rect 9262 11192 9954 11248
rect 10010 11192 10015 11248
rect 9262 11190 10015 11192
rect 8201 11187 8267 11190
rect 8569 11187 8635 11190
rect 9949 11187 10015 11190
rect 10593 11250 10659 11253
rect 10780 11250 10840 11598
rect 10593 11248 10840 11250
rect 10593 11192 10598 11248
rect 10654 11192 10840 11248
rect 10593 11190 10840 11192
rect 10593 11187 10659 11190
rect 8109 11114 8175 11117
rect 8477 11114 8543 11117
rect 8109 11112 8543 11114
rect 8109 11056 8114 11112
rect 8170 11056 8482 11112
rect 8538 11056 8543 11112
rect 8109 11054 8543 11056
rect 8109 11051 8175 11054
rect 8477 11051 8543 11054
rect 9673 11114 9739 11117
rect 10918 11114 10978 11870
rect 11424 11250 11484 13094
rect 13506 13088 14702 13089
rect 13506 13024 13512 13088
rect 13576 13024 13592 13088
rect 13656 13024 13672 13088
rect 13736 13024 13752 13088
rect 13816 13024 13832 13088
rect 13896 13024 13912 13088
rect 13976 13024 13992 13088
rect 14056 13024 14072 13088
rect 14136 13024 14152 13088
rect 14216 13024 14232 13088
rect 14296 13024 14312 13088
rect 14376 13024 14392 13088
rect 14456 13024 14472 13088
rect 14536 13024 14552 13088
rect 14616 13024 14632 13088
rect 14696 13024 14702 13088
rect 13506 13023 14702 13024
rect 11789 13016 11855 13021
rect 11789 12960 11794 13016
rect 11850 12960 11855 13016
rect 11789 12955 11855 12960
rect 11792 12613 11852 12955
rect 11789 12608 11855 12613
rect 11789 12552 11794 12608
rect 11850 12552 11855 12608
rect 11789 12547 11855 12552
rect 12249 12610 12315 12613
rect 12249 12608 12634 12610
rect 12249 12552 12254 12608
rect 12310 12552 12634 12608
rect 12249 12550 12634 12552
rect 12249 12547 12315 12550
rect 12341 12474 12407 12477
rect 12206 12472 12407 12474
rect 12206 12416 12346 12472
rect 12402 12416 12407 12472
rect 12206 12414 12407 12416
rect 12206 12069 12266 12414
rect 12341 12411 12407 12414
rect 12341 12202 12407 12205
rect 12574 12202 12634 12550
rect 17506 12544 18702 12545
rect 17506 12480 17512 12544
rect 17576 12480 17592 12544
rect 17656 12480 17672 12544
rect 17736 12480 17752 12544
rect 17816 12480 17832 12544
rect 17896 12480 17912 12544
rect 17976 12480 17992 12544
rect 18056 12480 18072 12544
rect 18136 12480 18152 12544
rect 18216 12480 18232 12544
rect 18296 12480 18312 12544
rect 18376 12480 18392 12544
rect 18456 12480 18472 12544
rect 18536 12480 18552 12544
rect 18616 12480 18632 12544
rect 18696 12480 18702 12544
rect 17506 12479 18702 12480
rect 12341 12200 12634 12202
rect 12341 12144 12346 12200
rect 12402 12144 12634 12200
rect 12341 12142 12634 12144
rect 12341 12139 12407 12142
rect 12206 12064 12315 12069
rect 12206 12008 12254 12064
rect 12310 12008 12315 12064
rect 12206 12006 12315 12008
rect 12249 12003 12315 12006
rect 13506 12000 14702 12001
rect 13506 11936 13512 12000
rect 13576 11936 13592 12000
rect 13656 11936 13672 12000
rect 13736 11936 13752 12000
rect 13816 11936 13832 12000
rect 13896 11936 13912 12000
rect 13976 11936 13992 12000
rect 14056 11936 14072 12000
rect 14136 11936 14152 12000
rect 14216 11936 14232 12000
rect 14296 11936 14312 12000
rect 14376 11936 14392 12000
rect 14456 11936 14472 12000
rect 14536 11936 14552 12000
rect 14616 11936 14632 12000
rect 14696 11936 14702 12000
rect 13506 11935 14702 11936
rect 11697 11792 11763 11797
rect 11697 11736 11702 11792
rect 11758 11736 11763 11792
rect 11697 11731 11763 11736
rect 12801 11794 12867 11797
rect 14641 11794 14707 11797
rect 12801 11792 14707 11794
rect 12801 11736 12806 11792
rect 12862 11736 14646 11792
rect 14702 11736 14707 11792
rect 12801 11734 14707 11736
rect 12801 11731 12867 11734
rect 14641 11731 14707 11734
rect 11700 11386 11760 11731
rect 18689 11658 18755 11661
rect 18822 11658 18828 11660
rect 18689 11656 18828 11658
rect 18689 11600 18694 11656
rect 18750 11600 18828 11656
rect 18689 11598 18828 11600
rect 18689 11595 18755 11598
rect 18822 11596 18828 11598
rect 18892 11596 18898 11660
rect 17506 11456 18702 11457
rect 17506 11392 17512 11456
rect 17576 11392 17592 11456
rect 17656 11392 17672 11456
rect 17736 11392 17752 11456
rect 17816 11392 17832 11456
rect 17896 11392 17912 11456
rect 17976 11392 17992 11456
rect 18056 11392 18072 11456
rect 18136 11392 18152 11456
rect 18216 11392 18232 11456
rect 18296 11392 18312 11456
rect 18376 11392 18392 11456
rect 18456 11392 18472 11456
rect 18536 11392 18552 11456
rect 18616 11392 18632 11456
rect 18696 11392 18702 11456
rect 17506 11391 18702 11392
rect 12341 11386 12407 11389
rect 11700 11350 11898 11386
rect 11700 11326 11794 11350
rect 11789 11294 11794 11326
rect 11850 11294 11898 11350
rect 11789 11292 11898 11294
rect 12206 11384 12407 11386
rect 12206 11328 12346 11384
rect 12402 11328 12407 11384
rect 12206 11326 12407 11328
rect 11789 11289 11855 11292
rect 12065 11250 12131 11253
rect 12206 11250 12266 11326
rect 12341 11323 12407 11326
rect 14457 11250 14523 11253
rect 11424 11190 11714 11250
rect 9673 11112 10978 11114
rect 9673 11056 9678 11112
rect 9734 11056 10978 11112
rect 9673 11054 10978 11056
rect 11654 11117 11714 11190
rect 12065 11248 12266 11250
rect 12065 11192 12070 11248
rect 12126 11192 12266 11248
rect 12065 11190 12266 11192
rect 12804 11248 14523 11250
rect 12804 11192 14462 11248
rect 14518 11192 14523 11248
rect 12804 11190 14523 11192
rect 12065 11187 12131 11190
rect 11654 11112 11763 11117
rect 11654 11056 11702 11112
rect 11758 11056 11763 11112
rect 11654 11054 11763 11056
rect 9673 11051 9739 11054
rect 11697 11051 11763 11054
rect 11973 11114 12039 11117
rect 12804 11114 12864 11190
rect 14457 11187 14523 11190
rect 15101 11250 15167 11253
rect 15285 11250 15351 11253
rect 16849 11250 16915 11253
rect 15101 11248 15351 11250
rect 15101 11192 15106 11248
rect 15162 11192 15290 11248
rect 15346 11192 15351 11248
rect 15101 11190 15351 11192
rect 15101 11187 15167 11190
rect 15285 11187 15351 11190
rect 16806 11248 16915 11250
rect 16806 11192 16854 11248
rect 16910 11192 16915 11248
rect 16806 11187 16915 11192
rect 11973 11112 12864 11114
rect 11973 11056 11978 11112
rect 12034 11056 12864 11112
rect 11973 11054 12864 11056
rect 11973 11051 12039 11054
rect 7833 10976 7899 10981
rect 7833 10920 7838 10976
rect 7894 10920 7899 10976
rect 7833 10915 7899 10920
rect 7974 10976 8083 10981
rect 7974 10920 8022 10976
rect 8078 10920 8083 10976
rect 7974 10918 8083 10920
rect 8017 10915 8083 10918
rect 8845 10978 8911 10981
rect 9857 10978 9923 10981
rect 8845 10976 9923 10978
rect 8845 10920 8850 10976
rect 8906 10920 9862 10976
rect 9918 10920 9923 10976
rect 8845 10918 9923 10920
rect 8845 10915 8911 10918
rect 9857 10915 9923 10918
rect 10961 10978 11027 10981
rect 11421 10978 11487 10981
rect 10961 10976 11487 10978
rect 10961 10920 10966 10976
rect 11022 10920 11426 10976
rect 11482 10920 11487 10976
rect 10961 10918 11487 10920
rect 10961 10915 11027 10918
rect 11421 10915 11487 10918
rect 16665 10978 16731 10981
rect 16806 10978 16866 11187
rect 16665 10976 16866 10978
rect 16665 10920 16670 10976
rect 16726 10920 16866 10976
rect 16665 10918 16866 10920
rect 16665 10915 16731 10918
rect 13506 10912 14702 10913
rect 13506 10848 13512 10912
rect 13576 10848 13592 10912
rect 13656 10848 13672 10912
rect 13736 10848 13752 10912
rect 13816 10848 13832 10912
rect 13896 10848 13912 10912
rect 13976 10848 13992 10912
rect 14056 10848 14072 10912
rect 14136 10848 14152 10912
rect 14216 10848 14232 10912
rect 14296 10848 14312 10912
rect 14376 10848 14392 10912
rect 14456 10848 14472 10912
rect 14536 10848 14552 10912
rect 14616 10848 14632 10912
rect 14696 10848 14702 10912
rect 13506 10847 14702 10848
rect 7925 10842 7991 10845
rect 7925 10840 12634 10842
rect 7925 10784 7930 10840
rect 7986 10784 12634 10840
rect 7925 10782 12634 10784
rect 7925 10779 7991 10782
rect 11789 10706 11855 10709
rect 7652 10646 8448 10706
rect 8388 10570 8448 10646
rect 9032 10704 11855 10706
rect 9032 10648 11794 10704
rect 11850 10648 11855 10704
rect 9032 10646 11855 10648
rect 8569 10570 8635 10573
rect 7284 10510 8080 10570
rect 8388 10568 8635 10570
rect 8388 10512 8574 10568
rect 8630 10512 8635 10568
rect 8388 10510 8635 10512
rect 7833 10434 7899 10437
rect 5720 10432 7899 10434
rect 5720 10376 7838 10432
rect 7894 10376 7899 10432
rect 5720 10374 7899 10376
rect 7833 10371 7899 10374
rect 1506 10368 2702 10369
rect 1506 10304 1512 10368
rect 1576 10304 1592 10368
rect 1656 10304 1672 10368
rect 1736 10304 1752 10368
rect 1816 10304 1832 10368
rect 1896 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2312 10368
rect 2376 10304 2392 10368
rect 2456 10304 2472 10368
rect 2536 10304 2552 10368
rect 2616 10304 2632 10368
rect 2696 10304 2702 10368
rect 1506 10303 2702 10304
rect 6545 10298 6611 10301
rect 7097 10298 7163 10301
rect 6545 10296 7163 10298
rect 6545 10240 6550 10296
rect 6606 10240 7102 10296
rect 7158 10240 7163 10296
rect 6545 10238 7163 10240
rect 6545 10235 6611 10238
rect 7097 10235 7163 10238
rect 7557 10298 7623 10301
rect 7741 10298 7807 10301
rect 7557 10296 7807 10298
rect 7557 10240 7562 10296
rect 7618 10240 7746 10296
rect 7802 10240 7807 10296
rect 7557 10238 7807 10240
rect 8020 10298 8080 10510
rect 8569 10507 8635 10510
rect 8201 10434 8267 10437
rect 9032 10434 9092 10646
rect 11789 10643 11855 10646
rect 9397 10570 9463 10573
rect 8201 10432 9092 10434
rect 8201 10376 8206 10432
rect 8262 10376 9092 10432
rect 8201 10374 9092 10376
rect 9262 10568 9463 10570
rect 9262 10512 9402 10568
rect 9458 10512 9463 10568
rect 9262 10510 9463 10512
rect 8201 10371 8267 10374
rect 9029 10298 9095 10301
rect 8020 10296 9095 10298
rect 8020 10240 9034 10296
rect 9090 10240 9095 10296
rect 8020 10238 9095 10240
rect 7557 10235 7623 10238
rect 7741 10235 7807 10238
rect 9029 10235 9095 10238
rect 13 10162 79 10165
rect 7741 10162 7807 10165
rect 13 10160 7807 10162
rect 13 10104 18 10160
rect 74 10104 7746 10160
rect 7802 10104 7807 10160
rect 13 10102 7807 10104
rect 13 10099 79 10102
rect 7741 10099 7807 10102
rect 8109 10160 8175 10165
rect 8109 10104 8114 10160
rect 8170 10104 8175 10160
rect 8109 10099 8175 10104
rect 9262 10162 9322 10510
rect 9397 10507 9463 10510
rect 9581 10570 9647 10573
rect 10133 10570 10199 10573
rect 9581 10568 10199 10570
rect 9581 10512 9586 10568
rect 9642 10512 10138 10568
rect 10194 10512 10199 10568
rect 9581 10510 10199 10512
rect 9581 10507 9647 10510
rect 10133 10507 10199 10510
rect 10685 10570 10751 10573
rect 11789 10570 11855 10573
rect 12433 10570 12499 10573
rect 10685 10568 11300 10570
rect 10685 10512 10690 10568
rect 10746 10512 11300 10568
rect 10685 10510 11300 10512
rect 10685 10507 10751 10510
rect 10777 10432 10843 10437
rect 10777 10376 10782 10432
rect 10838 10376 10843 10432
rect 10777 10371 10843 10376
rect 9506 10368 10702 10369
rect 9506 10304 9512 10368
rect 9576 10304 9592 10368
rect 9656 10304 9672 10368
rect 9736 10304 9752 10368
rect 9816 10304 9832 10368
rect 9896 10304 9912 10368
rect 9976 10304 9992 10368
rect 10056 10304 10072 10368
rect 10136 10304 10152 10368
rect 10216 10304 10232 10368
rect 10296 10304 10312 10368
rect 10376 10304 10392 10368
rect 10456 10304 10472 10368
rect 10536 10304 10552 10368
rect 10616 10304 10632 10368
rect 10696 10304 10702 10368
rect 9506 10303 10702 10304
rect 9397 10162 9463 10165
rect 9262 10160 9463 10162
rect 9262 10104 9402 10160
rect 9458 10104 9463 10160
rect 9262 10102 9463 10104
rect 9397 10099 9463 10102
rect 9765 10162 9831 10165
rect 10780 10162 10840 10371
rect 9765 10160 10840 10162
rect 9765 10104 9770 10160
rect 9826 10104 10840 10160
rect 9765 10102 10840 10104
rect 9765 10099 9831 10102
rect 3417 10026 3483 10029
rect 4981 10026 5047 10029
rect 3417 10024 5047 10026
rect 3417 9968 3422 10024
rect 3478 9968 4986 10024
rect 5042 9968 5047 10024
rect 3417 9966 5047 9968
rect 3417 9963 3483 9966
rect 4981 9963 5047 9966
rect 6637 10026 6703 10029
rect 8112 10026 8172 10099
rect 6637 10024 8172 10026
rect 6637 9968 6642 10024
rect 6698 9968 8172 10024
rect 6637 9966 8172 9968
rect 6637 9963 6703 9966
rect 11240 9893 11300 10510
rect 11789 10568 12499 10570
rect 11789 10512 11794 10568
rect 11850 10512 12438 10568
rect 12494 10512 12499 10568
rect 11789 10510 12499 10512
rect 11789 10507 11855 10510
rect 12433 10507 12499 10510
rect 12433 10434 12499 10437
rect 12574 10434 12634 10782
rect 18873 10706 18939 10709
rect 19006 10706 19012 10708
rect 18873 10704 19012 10706
rect 18873 10648 18878 10704
rect 18934 10648 19012 10704
rect 18873 10646 19012 10648
rect 18873 10643 18939 10646
rect 19006 10644 19012 10646
rect 19076 10644 19082 10708
rect 14733 10570 14799 10573
rect 16021 10570 16087 10573
rect 14733 10568 16087 10570
rect 14733 10512 14738 10568
rect 14794 10512 16026 10568
rect 16082 10512 16087 10568
rect 14733 10510 16087 10512
rect 14733 10507 14799 10510
rect 16021 10507 16087 10510
rect 12433 10432 12634 10434
rect 12433 10376 12438 10432
rect 12494 10376 12634 10432
rect 12433 10374 12634 10376
rect 12433 10371 12499 10374
rect 17506 10368 18702 10369
rect 17506 10304 17512 10368
rect 17576 10304 17592 10368
rect 17656 10304 17672 10368
rect 17736 10304 17752 10368
rect 17816 10304 17832 10368
rect 17896 10304 17912 10368
rect 17976 10304 17992 10368
rect 18056 10304 18072 10368
rect 18136 10304 18152 10368
rect 18216 10304 18232 10368
rect 18296 10304 18312 10368
rect 18376 10304 18392 10368
rect 18456 10304 18472 10368
rect 18536 10304 18552 10368
rect 18616 10304 18632 10368
rect 18696 10304 18702 10368
rect 17506 10303 18702 10304
rect 11697 10160 11763 10165
rect 11697 10104 11702 10160
rect 11758 10104 11763 10160
rect 11697 10099 11763 10104
rect 12157 10162 12223 10165
rect 14457 10162 14523 10165
rect 12157 10160 15578 10162
rect 12157 10104 12162 10160
rect 12218 10104 14462 10160
rect 14518 10104 15578 10160
rect 12157 10102 15578 10104
rect 12157 10099 12223 10102
rect 14457 10099 14523 10102
rect 11237 9888 11303 9893
rect 11237 9832 11242 9888
rect 11298 9832 11303 9888
rect 11237 9827 11303 9832
rect 5506 9824 6702 9825
rect 5506 9760 5512 9824
rect 5576 9760 5592 9824
rect 5656 9760 5672 9824
rect 5736 9760 5752 9824
rect 5816 9760 5832 9824
rect 5896 9760 5912 9824
rect 5976 9760 5992 9824
rect 6056 9760 6072 9824
rect 6136 9760 6152 9824
rect 6216 9760 6232 9824
rect 6296 9760 6312 9824
rect 6376 9760 6392 9824
rect 6456 9760 6472 9824
rect 6536 9760 6552 9824
rect 6616 9760 6632 9824
rect 6696 9760 6702 9824
rect 5506 9759 6702 9760
rect 5073 9618 5139 9621
rect 8017 9618 8083 9621
rect 5073 9616 8083 9618
rect 5073 9560 5078 9616
rect 5134 9560 8022 9616
rect 8078 9560 8083 9616
rect 5073 9558 8083 9560
rect 5073 9555 5139 9558
rect 8017 9555 8083 9558
rect 11329 9618 11395 9621
rect 11700 9618 11760 10099
rect 14273 10026 14339 10029
rect 14273 10024 14842 10026
rect 14273 9968 14278 10024
rect 14334 9968 14842 10024
rect 14273 9966 14842 9968
rect 14273 9963 14339 9966
rect 13261 9890 13327 9893
rect 13261 9888 13370 9890
rect 13261 9832 13266 9888
rect 13322 9832 13370 9888
rect 13261 9827 13370 9832
rect 11329 9616 11760 9618
rect 11329 9560 11334 9616
rect 11390 9560 11760 9616
rect 11329 9558 11760 9560
rect 13310 9621 13370 9827
rect 13506 9824 14702 9825
rect 13506 9760 13512 9824
rect 13576 9760 13592 9824
rect 13656 9760 13672 9824
rect 13736 9760 13752 9824
rect 13816 9760 13832 9824
rect 13896 9760 13912 9824
rect 13976 9760 13992 9824
rect 14056 9760 14072 9824
rect 14136 9760 14152 9824
rect 14216 9760 14232 9824
rect 14296 9760 14312 9824
rect 14376 9760 14392 9824
rect 14456 9760 14472 9824
rect 14536 9760 14552 9824
rect 14616 9760 14632 9824
rect 14696 9760 14702 9824
rect 13506 9759 14702 9760
rect 13310 9616 13419 9621
rect 13310 9560 13358 9616
rect 13414 9560 13419 9616
rect 13310 9558 13419 9560
rect 11329 9555 11395 9558
rect 7833 9482 7899 9485
rect 10685 9482 10751 9485
rect 7833 9480 10751 9482
rect 7833 9424 7838 9480
rect 7894 9424 10690 9480
rect 10746 9424 10751 9480
rect 7833 9422 10751 9424
rect 7833 9419 7899 9422
rect 10685 9419 10751 9422
rect 11700 9346 11760 9558
rect 13353 9555 13419 9558
rect 14641 9618 14707 9621
rect 14782 9618 14842 9966
rect 14641 9616 14842 9618
rect 14641 9560 14646 9616
rect 14702 9560 14842 9616
rect 14641 9558 14842 9560
rect 14641 9555 14707 9558
rect 13813 9482 13879 9485
rect 15518 9482 15578 10102
rect 15745 9618 15811 9621
rect 15745 9616 16130 9618
rect 15745 9560 15750 9616
rect 15806 9560 16130 9616
rect 15745 9558 16130 9560
rect 15745 9555 15811 9558
rect 15745 9482 15811 9485
rect 13813 9480 15811 9482
rect 13813 9424 13818 9480
rect 13874 9424 15750 9480
rect 15806 9424 15811 9480
rect 13813 9422 15811 9424
rect 13813 9419 13879 9422
rect 15745 9419 15811 9422
rect 16070 9346 16130 9558
rect 17953 9482 18019 9485
rect 16392 9480 18019 9482
rect 16392 9424 17958 9480
rect 18014 9424 18019 9480
rect 16392 9422 18019 9424
rect 16205 9346 16271 9349
rect 11700 9286 15946 9346
rect 16070 9344 16271 9346
rect 16070 9288 16210 9344
rect 16266 9288 16271 9344
rect 16070 9286 16271 9288
rect 1506 9280 2702 9281
rect 1506 9216 1512 9280
rect 1576 9216 1592 9280
rect 1656 9216 1672 9280
rect 1736 9216 1752 9280
rect 1816 9216 1832 9280
rect 1896 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2312 9280
rect 2376 9216 2392 9280
rect 2456 9216 2472 9280
rect 2536 9216 2552 9280
rect 2616 9216 2632 9280
rect 2696 9216 2702 9280
rect 1506 9215 2702 9216
rect 9506 9280 10702 9281
rect 9506 9216 9512 9280
rect 9576 9216 9592 9280
rect 9656 9216 9672 9280
rect 9736 9216 9752 9280
rect 9816 9216 9832 9280
rect 9896 9216 9912 9280
rect 9976 9216 9992 9280
rect 10056 9216 10072 9280
rect 10136 9216 10152 9280
rect 10216 9216 10232 9280
rect 10296 9216 10312 9280
rect 10376 9216 10392 9280
rect 10456 9216 10472 9280
rect 10536 9216 10552 9280
rect 10616 9216 10632 9280
rect 10696 9216 10702 9280
rect 9506 9215 10702 9216
rect 11053 9210 11119 9213
rect 13537 9210 13603 9213
rect 11053 9208 13603 9210
rect 11053 9152 11058 9208
rect 11114 9152 13542 9208
rect 13598 9152 13603 9208
rect 11053 9150 13603 9152
rect 15886 9210 15946 9286
rect 16205 9283 16271 9286
rect 16392 9210 16452 9422
rect 17953 9419 18019 9422
rect 18689 9482 18755 9485
rect 19190 9482 19196 9484
rect 18689 9480 19196 9482
rect 18689 9424 18694 9480
rect 18750 9424 19196 9480
rect 18689 9422 19196 9424
rect 18689 9419 18755 9422
rect 19190 9420 19196 9422
rect 19260 9420 19266 9484
rect 17506 9280 18702 9281
rect 17506 9216 17512 9280
rect 17576 9216 17592 9280
rect 17656 9216 17672 9280
rect 17736 9216 17752 9280
rect 17816 9216 17832 9280
rect 17896 9216 17912 9280
rect 17976 9216 17992 9280
rect 18056 9216 18072 9280
rect 18136 9216 18152 9280
rect 18216 9216 18232 9280
rect 18296 9216 18312 9280
rect 18376 9216 18392 9280
rect 18456 9216 18472 9280
rect 18536 9216 18552 9280
rect 18616 9216 18632 9280
rect 18696 9216 18702 9280
rect 17506 9215 18702 9216
rect 15886 9150 16452 9210
rect 11053 9147 11119 9150
rect 13537 9147 13603 9150
rect 4153 9074 4219 9077
rect 11053 9074 11119 9077
rect 18137 9074 18203 9077
rect 4153 9072 8310 9074
rect 4153 9016 4158 9072
rect 4214 9016 8310 9072
rect 4153 9014 8310 9016
rect 4153 9011 4219 9014
rect 8250 8938 8310 9014
rect 11053 9072 18203 9074
rect 11053 9016 11058 9072
rect 11114 9016 18142 9072
rect 18198 9016 18203 9072
rect 11053 9014 18203 9016
rect 11053 9011 11119 9014
rect 18137 9011 18203 9014
rect 13169 8938 13235 8941
rect 13813 8938 13879 8941
rect 8250 8936 13235 8938
rect 8250 8880 13174 8936
rect 13230 8880 13235 8936
rect 8250 8878 13235 8880
rect 13169 8875 13235 8878
rect 13310 8936 13879 8938
rect 13310 8880 13818 8936
rect 13874 8880 13879 8936
rect 13310 8878 13879 8880
rect 13169 8802 13235 8805
rect 13310 8802 13370 8878
rect 13813 8875 13879 8878
rect 14549 8938 14615 8941
rect 14549 8936 14842 8938
rect 14549 8880 14554 8936
rect 14610 8880 14842 8936
rect 14549 8878 14842 8880
rect 14549 8875 14615 8878
rect 13169 8800 13370 8802
rect 13169 8744 13174 8800
rect 13230 8744 13370 8800
rect 13169 8742 13370 8744
rect 13169 8739 13235 8742
rect 5506 8736 6702 8737
rect 5506 8672 5512 8736
rect 5576 8672 5592 8736
rect 5656 8672 5672 8736
rect 5736 8672 5752 8736
rect 5816 8672 5832 8736
rect 5896 8672 5912 8736
rect 5976 8672 5992 8736
rect 6056 8672 6072 8736
rect 6136 8672 6152 8736
rect 6216 8672 6232 8736
rect 6296 8672 6312 8736
rect 6376 8672 6392 8736
rect 6456 8672 6472 8736
rect 6536 8672 6552 8736
rect 6616 8672 6632 8736
rect 6696 8672 6702 8736
rect 5506 8671 6702 8672
rect 13506 8736 14702 8737
rect 13506 8672 13512 8736
rect 13576 8672 13592 8736
rect 13656 8672 13672 8736
rect 13736 8672 13752 8736
rect 13816 8672 13832 8736
rect 13896 8672 13912 8736
rect 13976 8672 13992 8736
rect 14056 8672 14072 8736
rect 14136 8672 14152 8736
rect 14216 8672 14232 8736
rect 14296 8672 14312 8736
rect 14376 8672 14392 8736
rect 14456 8672 14472 8736
rect 14536 8672 14552 8736
rect 14616 8672 14632 8736
rect 14696 8672 14702 8736
rect 13506 8671 14702 8672
rect 7097 8666 7163 8669
rect 12709 8666 12775 8669
rect 7097 8664 12775 8666
rect 7097 8608 7102 8664
rect 7158 8608 12714 8664
rect 12770 8608 12775 8664
rect 7097 8606 12775 8608
rect 7097 8603 7163 8606
rect 12709 8603 12775 8606
rect 7373 8530 7439 8533
rect 7741 8530 7807 8533
rect 7373 8528 7807 8530
rect 7373 8472 7378 8528
rect 7434 8472 7746 8528
rect 7802 8472 7807 8528
rect 7373 8470 7807 8472
rect 7373 8467 7439 8470
rect 7741 8467 7807 8470
rect 14089 8530 14155 8533
rect 14782 8530 14842 8878
rect 14089 8528 14842 8530
rect 14089 8472 14094 8528
rect 14150 8472 14842 8528
rect 14089 8470 14842 8472
rect 14089 8467 14155 8470
rect 5441 8394 5507 8397
rect 14825 8394 14891 8397
rect 5441 8392 14891 8394
rect 5441 8336 5446 8392
rect 5502 8336 14830 8392
rect 14886 8336 14891 8392
rect 5441 8334 14891 8336
rect 5441 8331 5507 8334
rect 14825 8331 14891 8334
rect 1506 8192 2702 8193
rect 1506 8128 1512 8192
rect 1576 8128 1592 8192
rect 1656 8128 1672 8192
rect 1736 8128 1752 8192
rect 1816 8128 1832 8192
rect 1896 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2312 8192
rect 2376 8128 2392 8192
rect 2456 8128 2472 8192
rect 2536 8128 2552 8192
rect 2616 8128 2632 8192
rect 2696 8128 2702 8192
rect 1506 8127 2702 8128
rect 9506 8192 10702 8193
rect 9506 8128 9512 8192
rect 9576 8128 9592 8192
rect 9656 8128 9672 8192
rect 9736 8128 9752 8192
rect 9816 8128 9832 8192
rect 9896 8128 9912 8192
rect 9976 8128 9992 8192
rect 10056 8128 10072 8192
rect 10136 8128 10152 8192
rect 10216 8128 10232 8192
rect 10296 8128 10312 8192
rect 10376 8128 10392 8192
rect 10456 8128 10472 8192
rect 10536 8128 10552 8192
rect 10616 8128 10632 8192
rect 10696 8128 10702 8192
rect 9506 8127 10702 8128
rect 17506 8192 18702 8193
rect 17506 8128 17512 8192
rect 17576 8128 17592 8192
rect 17656 8128 17672 8192
rect 17736 8128 17752 8192
rect 17816 8128 17832 8192
rect 17896 8128 17912 8192
rect 17976 8128 17992 8192
rect 18056 8128 18072 8192
rect 18136 8128 18152 8192
rect 18216 8128 18232 8192
rect 18296 8128 18312 8192
rect 18376 8128 18392 8192
rect 18456 8128 18472 8192
rect 18536 8128 18552 8192
rect 18616 8128 18632 8192
rect 18696 8128 18702 8192
rect 17506 8127 18702 8128
rect 12433 8122 12499 8125
rect 15377 8122 15443 8125
rect 12433 8120 15443 8122
rect 12433 8064 12438 8120
rect 12494 8064 15382 8120
rect 15438 8064 15443 8120
rect 12433 8062 15443 8064
rect 12433 8059 12499 8062
rect 15377 8059 15443 8062
rect 8845 7850 8911 7853
rect 14549 7850 14615 7853
rect 7606 7848 14615 7850
rect 7606 7792 8850 7848
rect 8906 7792 14554 7848
rect 14610 7792 14615 7848
rect 7606 7790 14615 7792
rect 5506 7648 6702 7649
rect 5506 7584 5512 7648
rect 5576 7584 5592 7648
rect 5656 7584 5672 7648
rect 5736 7584 5752 7648
rect 5816 7584 5832 7648
rect 5896 7584 5912 7648
rect 5976 7584 5992 7648
rect 6056 7584 6072 7648
rect 6136 7584 6152 7648
rect 6216 7584 6232 7648
rect 6296 7584 6312 7648
rect 6376 7584 6392 7648
rect 6456 7584 6472 7648
rect 6536 7584 6552 7648
rect 6616 7584 6632 7648
rect 6696 7584 6702 7648
rect 5506 7583 6702 7584
rect 5717 7442 5783 7445
rect 7465 7442 7531 7445
rect 5717 7440 7531 7442
rect 5717 7384 5722 7440
rect 5778 7384 7470 7440
rect 7526 7384 7531 7440
rect 5717 7382 7531 7384
rect 5717 7379 5783 7382
rect 7465 7379 7531 7382
rect 5533 7306 5599 7309
rect 7606 7306 7666 7790
rect 8845 7787 8911 7790
rect 14549 7787 14615 7790
rect 11237 7714 11303 7717
rect 11421 7714 11487 7717
rect 11237 7712 11487 7714
rect 11237 7656 11242 7712
rect 11298 7656 11426 7712
rect 11482 7656 11487 7712
rect 11237 7654 11487 7656
rect 11237 7651 11303 7654
rect 11421 7651 11487 7654
rect 13506 7648 14702 7649
rect 13506 7584 13512 7648
rect 13576 7584 13592 7648
rect 13656 7584 13672 7648
rect 13736 7584 13752 7648
rect 13816 7584 13832 7648
rect 13896 7584 13912 7648
rect 13976 7584 13992 7648
rect 14056 7584 14072 7648
rect 14136 7584 14152 7648
rect 14216 7584 14232 7648
rect 14296 7584 14312 7648
rect 14376 7584 14392 7648
rect 14456 7584 14472 7648
rect 14536 7584 14552 7648
rect 14616 7584 14632 7648
rect 14696 7584 14702 7648
rect 13506 7583 14702 7584
rect 19057 7578 19123 7581
rect 19333 7578 19399 7581
rect 19057 7576 19399 7578
rect 19057 7520 19062 7576
rect 19118 7520 19338 7576
rect 19394 7520 19399 7576
rect 19057 7518 19399 7520
rect 19057 7515 19123 7518
rect 19333 7515 19399 7518
rect 5533 7304 7666 7306
rect 5533 7248 5538 7304
rect 5594 7248 7666 7304
rect 5533 7246 7666 7248
rect 5533 7243 5599 7246
rect 12617 7170 12683 7173
rect 16205 7170 16271 7173
rect 12617 7168 16271 7170
rect 12617 7112 12622 7168
rect 12678 7112 16210 7168
rect 16266 7112 16271 7168
rect 12617 7110 16271 7112
rect 12617 7107 12683 7110
rect 16205 7107 16271 7110
rect 1506 7104 2702 7105
rect 1506 7040 1512 7104
rect 1576 7040 1592 7104
rect 1656 7040 1672 7104
rect 1736 7040 1752 7104
rect 1816 7040 1832 7104
rect 1896 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2312 7104
rect 2376 7040 2392 7104
rect 2456 7040 2472 7104
rect 2536 7040 2552 7104
rect 2616 7040 2632 7104
rect 2696 7040 2702 7104
rect 1506 7039 2702 7040
rect 9506 7104 10702 7105
rect 9506 7040 9512 7104
rect 9576 7040 9592 7104
rect 9656 7040 9672 7104
rect 9736 7040 9752 7104
rect 9816 7040 9832 7104
rect 9896 7040 9912 7104
rect 9976 7040 9992 7104
rect 10056 7040 10072 7104
rect 10136 7040 10152 7104
rect 10216 7040 10232 7104
rect 10296 7040 10312 7104
rect 10376 7040 10392 7104
rect 10456 7040 10472 7104
rect 10536 7040 10552 7104
rect 10616 7040 10632 7104
rect 10696 7040 10702 7104
rect 9506 7039 10702 7040
rect 17506 7104 18702 7105
rect 17506 7040 17512 7104
rect 17576 7040 17592 7104
rect 17656 7040 17672 7104
rect 17736 7040 17752 7104
rect 17816 7040 17832 7104
rect 17896 7040 17912 7104
rect 17976 7040 17992 7104
rect 18056 7040 18072 7104
rect 18136 7040 18152 7104
rect 18216 7040 18232 7104
rect 18296 7040 18312 7104
rect 18376 7040 18392 7104
rect 18456 7040 18472 7104
rect 18536 7040 18552 7104
rect 18616 7040 18632 7104
rect 18696 7040 18702 7104
rect 17506 7039 18702 7040
rect 11697 7034 11763 7037
rect 15469 7034 15535 7037
rect 11697 7032 15535 7034
rect 11697 6976 11702 7032
rect 11758 6976 15474 7032
rect 15530 6976 15535 7032
rect 11697 6974 15535 6976
rect 11697 6971 11763 6974
rect 15469 6971 15535 6974
rect 6821 6898 6887 6901
rect 11053 6898 11119 6901
rect 6821 6896 11119 6898
rect 6821 6840 6826 6896
rect 6882 6840 11058 6896
rect 11114 6840 11119 6896
rect 6821 6838 11119 6840
rect 6821 6835 6887 6838
rect 11053 6835 11119 6838
rect 12433 6762 12499 6765
rect 15193 6762 15259 6765
rect 16021 6762 16087 6765
rect 16481 6762 16547 6765
rect 12433 6760 16547 6762
rect 12433 6704 12438 6760
rect 12494 6704 15198 6760
rect 15254 6704 16026 6760
rect 16082 6704 16486 6760
rect 16542 6704 16547 6760
rect 12433 6702 16547 6704
rect 12433 6699 12499 6702
rect 15193 6699 15259 6702
rect 16021 6699 16087 6702
rect 16481 6699 16547 6702
rect 5506 6560 6702 6561
rect 5506 6496 5512 6560
rect 5576 6496 5592 6560
rect 5656 6496 5672 6560
rect 5736 6496 5752 6560
rect 5816 6496 5832 6560
rect 5896 6496 5912 6560
rect 5976 6496 5992 6560
rect 6056 6496 6072 6560
rect 6136 6496 6152 6560
rect 6216 6496 6232 6560
rect 6296 6496 6312 6560
rect 6376 6496 6392 6560
rect 6456 6496 6472 6560
rect 6536 6496 6552 6560
rect 6616 6496 6632 6560
rect 6696 6496 6702 6560
rect 5506 6495 6702 6496
rect 13506 6560 14702 6561
rect 13506 6496 13512 6560
rect 13576 6496 13592 6560
rect 13656 6496 13672 6560
rect 13736 6496 13752 6560
rect 13816 6496 13832 6560
rect 13896 6496 13912 6560
rect 13976 6496 13992 6560
rect 14056 6496 14072 6560
rect 14136 6496 14152 6560
rect 14216 6496 14232 6560
rect 14296 6496 14312 6560
rect 14376 6496 14392 6560
rect 14456 6496 14472 6560
rect 14536 6496 14552 6560
rect 14616 6496 14632 6560
rect 14696 6496 14702 6560
rect 13506 6495 14702 6496
rect 12525 6354 12591 6357
rect 14549 6354 14615 6357
rect 15561 6354 15627 6357
rect 12525 6352 15627 6354
rect 12525 6296 12530 6352
rect 12586 6296 14554 6352
rect 14610 6296 15566 6352
rect 15622 6296 15627 6352
rect 12525 6294 15627 6296
rect 12525 6291 12591 6294
rect 14549 6291 14615 6294
rect 15561 6291 15627 6294
rect 5349 6218 5415 6221
rect 18781 6218 18847 6221
rect 5349 6216 18847 6218
rect 5349 6160 5354 6216
rect 5410 6160 18786 6216
rect 18842 6160 18847 6216
rect 5349 6158 18847 6160
rect 5349 6155 5415 6158
rect 18781 6155 18847 6158
rect 14549 6082 14615 6085
rect 15377 6082 15443 6085
rect 16849 6082 16915 6085
rect 14549 6080 16915 6082
rect 14549 6024 14554 6080
rect 14610 6024 15382 6080
rect 15438 6024 16854 6080
rect 16910 6024 16915 6080
rect 14549 6022 16915 6024
rect 14549 6019 14615 6022
rect 15377 6019 15443 6022
rect 16849 6019 16915 6022
rect 1506 6016 2702 6017
rect 1506 5952 1512 6016
rect 1576 5952 1592 6016
rect 1656 5952 1672 6016
rect 1736 5952 1752 6016
rect 1816 5952 1832 6016
rect 1896 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2312 6016
rect 2376 5952 2392 6016
rect 2456 5952 2472 6016
rect 2536 5952 2552 6016
rect 2616 5952 2632 6016
rect 2696 5952 2702 6016
rect 1506 5951 2702 5952
rect 9506 6016 10702 6017
rect 9506 5952 9512 6016
rect 9576 5952 9592 6016
rect 9656 5952 9672 6016
rect 9736 5952 9752 6016
rect 9816 5952 9832 6016
rect 9896 5952 9912 6016
rect 9976 5952 9992 6016
rect 10056 5952 10072 6016
rect 10136 5952 10152 6016
rect 10216 5952 10232 6016
rect 10296 5952 10312 6016
rect 10376 5952 10392 6016
rect 10456 5952 10472 6016
rect 10536 5952 10552 6016
rect 10616 5952 10632 6016
rect 10696 5952 10702 6016
rect 9506 5951 10702 5952
rect 17506 6016 18702 6017
rect 17506 5952 17512 6016
rect 17576 5952 17592 6016
rect 17656 5952 17672 6016
rect 17736 5952 17752 6016
rect 17816 5952 17832 6016
rect 17896 5952 17912 6016
rect 17976 5952 17992 6016
rect 18056 5952 18072 6016
rect 18136 5952 18152 6016
rect 18216 5952 18232 6016
rect 18296 5952 18312 6016
rect 18376 5952 18392 6016
rect 18456 5952 18472 6016
rect 18536 5952 18552 6016
rect 18616 5952 18632 6016
rect 18696 5952 18702 6016
rect 17506 5951 18702 5952
rect 18045 5810 18111 5813
rect 19057 5810 19123 5813
rect 18045 5808 19123 5810
rect 18045 5752 18050 5808
rect 18106 5752 19062 5808
rect 19118 5752 19123 5808
rect 18045 5750 19123 5752
rect 18045 5747 18111 5750
rect 19057 5747 19123 5750
rect 16389 5538 16455 5541
rect 19149 5538 19215 5541
rect 16389 5536 19215 5538
rect 16389 5480 16394 5536
rect 16450 5480 19154 5536
rect 19210 5480 19215 5536
rect 16389 5478 19215 5480
rect 16389 5475 16455 5478
rect 19149 5475 19215 5478
rect 5506 5472 6702 5473
rect 5506 5408 5512 5472
rect 5576 5408 5592 5472
rect 5656 5408 5672 5472
rect 5736 5408 5752 5472
rect 5816 5408 5832 5472
rect 5896 5408 5912 5472
rect 5976 5408 5992 5472
rect 6056 5408 6072 5472
rect 6136 5408 6152 5472
rect 6216 5408 6232 5472
rect 6296 5408 6312 5472
rect 6376 5408 6392 5472
rect 6456 5408 6472 5472
rect 6536 5408 6552 5472
rect 6616 5408 6632 5472
rect 6696 5408 6702 5472
rect 5506 5407 6702 5408
rect 13506 5472 14702 5473
rect 13506 5408 13512 5472
rect 13576 5408 13592 5472
rect 13656 5408 13672 5472
rect 13736 5408 13752 5472
rect 13816 5408 13832 5472
rect 13896 5408 13912 5472
rect 13976 5408 13992 5472
rect 14056 5408 14072 5472
rect 14136 5408 14152 5472
rect 14216 5408 14232 5472
rect 14296 5408 14312 5472
rect 14376 5408 14392 5472
rect 14456 5408 14472 5472
rect 14536 5408 14552 5472
rect 14616 5408 14632 5472
rect 14696 5408 14702 5472
rect 13506 5407 14702 5408
rect 6453 5266 6519 5269
rect 18965 5266 19031 5269
rect 6453 5264 19031 5266
rect 6453 5208 6458 5264
rect 6514 5208 18970 5264
rect 19026 5208 19031 5264
rect 6453 5206 19031 5208
rect 6453 5203 6519 5206
rect 18965 5203 19031 5206
rect 18822 5068 18828 5132
rect 18892 5130 18898 5132
rect 19701 5130 19767 5133
rect 18892 5128 19767 5130
rect 18892 5072 19706 5128
rect 19762 5072 19767 5128
rect 18892 5070 19767 5072
rect 18892 5068 18898 5070
rect 19701 5067 19767 5070
rect 1506 4928 2702 4929
rect 1506 4864 1512 4928
rect 1576 4864 1592 4928
rect 1656 4864 1672 4928
rect 1736 4864 1752 4928
rect 1816 4864 1832 4928
rect 1896 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2312 4928
rect 2376 4864 2392 4928
rect 2456 4864 2472 4928
rect 2536 4864 2552 4928
rect 2616 4864 2632 4928
rect 2696 4864 2702 4928
rect 1506 4863 2702 4864
rect 9506 4928 10702 4929
rect 9506 4864 9512 4928
rect 9576 4864 9592 4928
rect 9656 4864 9672 4928
rect 9736 4864 9752 4928
rect 9816 4864 9832 4928
rect 9896 4864 9912 4928
rect 9976 4864 9992 4928
rect 10056 4864 10072 4928
rect 10136 4864 10152 4928
rect 10216 4864 10232 4928
rect 10296 4864 10312 4928
rect 10376 4864 10392 4928
rect 10456 4864 10472 4928
rect 10536 4864 10552 4928
rect 10616 4864 10632 4928
rect 10696 4864 10702 4928
rect 9506 4863 10702 4864
rect 17506 4928 18702 4929
rect 17506 4864 17512 4928
rect 17576 4864 17592 4928
rect 17656 4864 17672 4928
rect 17736 4864 17752 4928
rect 17816 4864 17832 4928
rect 17896 4864 17912 4928
rect 17976 4864 17992 4928
rect 18056 4864 18072 4928
rect 18136 4864 18152 4928
rect 18216 4864 18232 4928
rect 18296 4864 18312 4928
rect 18376 4864 18392 4928
rect 18456 4864 18472 4928
rect 18536 4864 18552 4928
rect 18616 4864 18632 4928
rect 18696 4864 18702 4928
rect 17506 4863 18702 4864
rect 657 4586 723 4589
rect 10685 4586 10751 4589
rect 19190 4586 19196 4588
rect 657 4584 996 4586
rect 657 4528 662 4584
rect 718 4528 996 4584
rect 657 4526 996 4528
rect 657 4523 723 4526
rect 0 4314 800 4344
rect 936 4314 996 4526
rect 10685 4584 19196 4586
rect 10685 4528 10690 4584
rect 10746 4528 19196 4584
rect 10685 4526 19196 4528
rect 10685 4523 10751 4526
rect 19190 4524 19196 4526
rect 19260 4524 19266 4588
rect 5506 4384 6702 4385
rect 5506 4320 5512 4384
rect 5576 4320 5592 4384
rect 5656 4320 5672 4384
rect 5736 4320 5752 4384
rect 5816 4320 5832 4384
rect 5896 4320 5912 4384
rect 5976 4320 5992 4384
rect 6056 4320 6072 4384
rect 6136 4320 6152 4384
rect 6216 4320 6232 4384
rect 6296 4320 6312 4384
rect 6376 4320 6392 4384
rect 6456 4320 6472 4384
rect 6536 4320 6552 4384
rect 6616 4320 6632 4384
rect 6696 4320 6702 4384
rect 5506 4319 6702 4320
rect 13506 4384 14702 4385
rect 13506 4320 13512 4384
rect 13576 4320 13592 4384
rect 13656 4320 13672 4384
rect 13736 4320 13752 4384
rect 13816 4320 13832 4384
rect 13896 4320 13912 4384
rect 13976 4320 13992 4384
rect 14056 4320 14072 4384
rect 14136 4320 14152 4384
rect 14216 4320 14232 4384
rect 14296 4320 14312 4384
rect 14376 4320 14392 4384
rect 14456 4320 14472 4384
rect 14536 4320 14552 4384
rect 14616 4320 14632 4384
rect 14696 4320 14702 4384
rect 13506 4319 14702 4320
rect 0 4254 996 4314
rect 0 4224 800 4254
rect 19006 4178 19012 4180
rect 18462 4118 19012 4178
rect 0 4042 800 4072
rect 1393 4042 1459 4045
rect 0 4040 1459 4042
rect 0 3984 1398 4040
rect 1454 3984 1459 4040
rect 0 3982 1459 3984
rect 0 3952 800 3982
rect 1393 3979 1459 3982
rect 7741 4042 7807 4045
rect 11053 4042 11119 4045
rect 7741 4040 11119 4042
rect 7741 3984 7746 4040
rect 7802 3984 11058 4040
rect 11114 3984 11119 4040
rect 7741 3982 11119 3984
rect 7741 3979 7807 3982
rect 11053 3979 11119 3982
rect 14181 4042 14247 4045
rect 18462 4042 18522 4118
rect 19006 4116 19012 4118
rect 19076 4116 19082 4180
rect 14181 4040 18522 4042
rect 14181 3984 14186 4040
rect 14242 3984 18522 4040
rect 14181 3982 18522 3984
rect 18689 4042 18755 4045
rect 19149 4042 19215 4045
rect 18689 4040 19215 4042
rect 18689 3984 18694 4040
rect 18750 3984 19154 4040
rect 19210 3984 19215 4040
rect 18689 3982 19215 3984
rect 14181 3979 14247 3982
rect 18689 3979 18755 3982
rect 19149 3979 19215 3982
rect 11237 3906 11303 3909
rect 12341 3906 12407 3909
rect 11237 3904 12407 3906
rect 11237 3848 11242 3904
rect 11298 3848 12346 3904
rect 12402 3848 12407 3904
rect 11237 3846 12407 3848
rect 11237 3843 11303 3846
rect 12341 3843 12407 3846
rect 1506 3840 2702 3841
rect 0 3770 800 3800
rect 1506 3776 1512 3840
rect 1576 3776 1592 3840
rect 1656 3776 1672 3840
rect 1736 3776 1752 3840
rect 1816 3776 1832 3840
rect 1896 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2312 3840
rect 2376 3776 2392 3840
rect 2456 3776 2472 3840
rect 2536 3776 2552 3840
rect 2616 3776 2632 3840
rect 2696 3776 2702 3840
rect 1506 3775 2702 3776
rect 9506 3840 10702 3841
rect 9506 3776 9512 3840
rect 9576 3776 9592 3840
rect 9656 3776 9672 3840
rect 9736 3776 9752 3840
rect 9816 3776 9832 3840
rect 9896 3776 9912 3840
rect 9976 3776 9992 3840
rect 10056 3776 10072 3840
rect 10136 3776 10152 3840
rect 10216 3776 10232 3840
rect 10296 3776 10312 3840
rect 10376 3776 10392 3840
rect 10456 3776 10472 3840
rect 10536 3776 10552 3840
rect 10616 3776 10632 3840
rect 10696 3776 10702 3840
rect 9506 3775 10702 3776
rect 17506 3840 18702 3841
rect 17506 3776 17512 3840
rect 17576 3776 17592 3840
rect 17656 3776 17672 3840
rect 17736 3776 17752 3840
rect 17816 3776 17832 3840
rect 17896 3776 17912 3840
rect 17976 3776 17992 3840
rect 18056 3776 18072 3840
rect 18136 3776 18152 3840
rect 18216 3776 18232 3840
rect 18296 3776 18312 3840
rect 18376 3776 18392 3840
rect 18456 3776 18472 3840
rect 18536 3776 18552 3840
rect 18616 3776 18632 3840
rect 18696 3776 18702 3840
rect 17506 3775 18702 3776
rect 933 3770 999 3773
rect 12709 3770 12775 3773
rect 14641 3770 14707 3773
rect 0 3768 999 3770
rect 0 3712 938 3768
rect 994 3712 999 3768
rect 0 3710 999 3712
rect 0 3680 800 3710
rect 933 3707 999 3710
rect 10918 3768 14707 3770
rect 10918 3712 12714 3768
rect 12770 3712 14646 3768
rect 14702 3712 14707 3768
rect 10918 3710 14707 3712
rect 5717 3634 5783 3637
rect 9121 3634 9187 3637
rect 5717 3632 9187 3634
rect 5717 3576 5722 3632
rect 5778 3576 9126 3632
rect 9182 3576 9187 3632
rect 5717 3574 9187 3576
rect 5717 3571 5783 3574
rect 9121 3571 9187 3574
rect 9581 3634 9647 3637
rect 10918 3634 10978 3710
rect 12709 3707 12775 3710
rect 14641 3707 14707 3710
rect 9581 3632 10978 3634
rect 9581 3576 9586 3632
rect 9642 3576 10978 3632
rect 9581 3574 10978 3576
rect 11053 3634 11119 3637
rect 16665 3634 16731 3637
rect 11053 3632 16731 3634
rect 11053 3576 11058 3632
rect 11114 3576 16670 3632
rect 16726 3576 16731 3632
rect 11053 3574 16731 3576
rect 9581 3571 9647 3574
rect 11053 3571 11119 3574
rect 16665 3571 16731 3574
rect 0 3498 800 3528
rect 1117 3498 1183 3501
rect 0 3496 1183 3498
rect 0 3440 1122 3496
rect 1178 3440 1183 3496
rect 0 3438 1183 3440
rect 0 3408 800 3438
rect 1117 3435 1183 3438
rect 8937 3498 9003 3501
rect 14273 3498 14339 3501
rect 8937 3496 14339 3498
rect 8937 3440 8942 3496
rect 8998 3440 14278 3496
rect 14334 3440 14339 3496
rect 8937 3438 14339 3440
rect 8937 3435 9003 3438
rect 14273 3435 14339 3438
rect 14457 3498 14523 3501
rect 17033 3498 17099 3501
rect 14457 3496 17099 3498
rect 14457 3440 14462 3496
rect 14518 3440 17038 3496
rect 17094 3440 17099 3496
rect 14457 3438 17099 3440
rect 14457 3435 14523 3438
rect 17033 3435 17099 3438
rect 10409 3362 10475 3365
rect 11053 3362 11119 3365
rect 10409 3360 11119 3362
rect 10409 3304 10414 3360
rect 10470 3304 11058 3360
rect 11114 3304 11119 3360
rect 10409 3302 11119 3304
rect 10409 3299 10475 3302
rect 11053 3299 11119 3302
rect 5506 3296 6702 3297
rect 0 3226 800 3256
rect 5506 3232 5512 3296
rect 5576 3232 5592 3296
rect 5656 3232 5672 3296
rect 5736 3232 5752 3296
rect 5816 3232 5832 3296
rect 5896 3232 5912 3296
rect 5976 3232 5992 3296
rect 6056 3232 6072 3296
rect 6136 3232 6152 3296
rect 6216 3232 6232 3296
rect 6296 3232 6312 3296
rect 6376 3232 6392 3296
rect 6456 3232 6472 3296
rect 6536 3232 6552 3296
rect 6616 3232 6632 3296
rect 6696 3232 6702 3296
rect 5506 3231 6702 3232
rect 13506 3296 14702 3297
rect 13506 3232 13512 3296
rect 13576 3232 13592 3296
rect 13656 3232 13672 3296
rect 13736 3232 13752 3296
rect 13816 3232 13832 3296
rect 13896 3232 13912 3296
rect 13976 3232 13992 3296
rect 14056 3232 14072 3296
rect 14136 3232 14152 3296
rect 14216 3232 14232 3296
rect 14296 3232 14312 3296
rect 14376 3232 14392 3296
rect 14456 3232 14472 3296
rect 14536 3232 14552 3296
rect 14616 3232 14632 3296
rect 14696 3232 14702 3296
rect 13506 3231 14702 3232
rect 1025 3226 1091 3229
rect 0 3224 1091 3226
rect 0 3168 1030 3224
rect 1086 3168 1091 3224
rect 0 3166 1091 3168
rect 0 3136 800 3166
rect 1025 3163 1091 3166
rect 10593 3226 10659 3229
rect 12985 3226 13051 3229
rect 10593 3224 13051 3226
rect 10593 3168 10598 3224
rect 10654 3168 12990 3224
rect 13046 3168 13051 3224
rect 10593 3166 13051 3168
rect 10593 3163 10659 3166
rect 12985 3163 13051 3166
rect 0 2954 800 2984
rect 933 2954 999 2957
rect 0 2952 999 2954
rect 0 2896 938 2952
rect 994 2896 999 2952
rect 0 2894 999 2896
rect 0 2864 800 2894
rect 933 2891 999 2894
rect 12709 2954 12775 2957
rect 19701 2954 19767 2957
rect 12709 2952 19767 2954
rect 12709 2896 12714 2952
rect 12770 2896 19706 2952
rect 19762 2896 19767 2952
rect 12709 2894 19767 2896
rect 12709 2891 12775 2894
rect 19701 2891 19767 2894
rect 10869 2818 10935 2821
rect 11697 2818 11763 2821
rect 10869 2816 11763 2818
rect 10869 2760 10874 2816
rect 10930 2760 11702 2816
rect 11758 2760 11763 2816
rect 10869 2758 11763 2760
rect 10869 2755 10935 2758
rect 11697 2755 11763 2758
rect 15101 2818 15167 2821
rect 16665 2818 16731 2821
rect 15101 2816 16731 2818
rect 15101 2760 15106 2816
rect 15162 2760 16670 2816
rect 16726 2760 16731 2816
rect 15101 2758 16731 2760
rect 15101 2755 15167 2758
rect 16665 2755 16731 2758
rect 1506 2752 2702 2753
rect 0 2682 800 2712
rect 1506 2688 1512 2752
rect 1576 2688 1592 2752
rect 1656 2688 1672 2752
rect 1736 2688 1752 2752
rect 1816 2688 1832 2752
rect 1896 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2312 2752
rect 2376 2688 2392 2752
rect 2456 2688 2472 2752
rect 2536 2688 2552 2752
rect 2616 2688 2632 2752
rect 2696 2688 2702 2752
rect 1506 2687 2702 2688
rect 9506 2752 10702 2753
rect 9506 2688 9512 2752
rect 9576 2688 9592 2752
rect 9656 2688 9672 2752
rect 9736 2688 9752 2752
rect 9816 2688 9832 2752
rect 9896 2688 9912 2752
rect 9976 2688 9992 2752
rect 10056 2688 10072 2752
rect 10136 2688 10152 2752
rect 10216 2688 10232 2752
rect 10296 2688 10312 2752
rect 10376 2688 10392 2752
rect 10456 2688 10472 2752
rect 10536 2688 10552 2752
rect 10616 2688 10632 2752
rect 10696 2688 10702 2752
rect 9506 2687 10702 2688
rect 17506 2752 18702 2753
rect 17506 2688 17512 2752
rect 17576 2688 17592 2752
rect 17656 2688 17672 2752
rect 17736 2688 17752 2752
rect 17816 2688 17832 2752
rect 17896 2688 17912 2752
rect 17976 2688 17992 2752
rect 18056 2688 18072 2752
rect 18136 2688 18152 2752
rect 18216 2688 18232 2752
rect 18296 2688 18312 2752
rect 18376 2688 18392 2752
rect 18456 2688 18472 2752
rect 18536 2688 18552 2752
rect 18616 2688 18632 2752
rect 18696 2688 18702 2752
rect 17506 2687 18702 2688
rect 0 2622 1410 2682
rect 0 2592 800 2622
rect 1350 2546 1410 2622
rect 3693 2546 3759 2549
rect 1350 2544 3759 2546
rect 1350 2488 3698 2544
rect 3754 2488 3759 2544
rect 1350 2486 3759 2488
rect 3693 2483 3759 2486
rect 13077 2546 13143 2549
rect 19793 2546 19859 2549
rect 13077 2544 19859 2546
rect 13077 2488 13082 2544
rect 13138 2488 19798 2544
rect 19854 2488 19859 2544
rect 13077 2486 19859 2488
rect 13077 2483 13143 2486
rect 19793 2483 19859 2486
rect 0 2410 800 2440
rect 933 2410 999 2413
rect 0 2408 999 2410
rect 0 2352 938 2408
rect 994 2352 999 2408
rect 0 2350 999 2352
rect 0 2320 800 2350
rect 933 2347 999 2350
rect 5506 2208 6702 2209
rect 0 2138 800 2168
rect 5506 2144 5512 2208
rect 5576 2144 5592 2208
rect 5656 2144 5672 2208
rect 5736 2144 5752 2208
rect 5816 2144 5832 2208
rect 5896 2144 5912 2208
rect 5976 2144 5992 2208
rect 6056 2144 6072 2208
rect 6136 2144 6152 2208
rect 6216 2144 6232 2208
rect 6296 2144 6312 2208
rect 6376 2144 6392 2208
rect 6456 2144 6472 2208
rect 6536 2144 6552 2208
rect 6616 2144 6632 2208
rect 6696 2144 6702 2208
rect 5506 2143 6702 2144
rect 13506 2208 14702 2209
rect 13506 2144 13512 2208
rect 13576 2144 13592 2208
rect 13656 2144 13672 2208
rect 13736 2144 13752 2208
rect 13816 2144 13832 2208
rect 13896 2144 13912 2208
rect 13976 2144 13992 2208
rect 14056 2144 14072 2208
rect 14136 2144 14152 2208
rect 14216 2144 14232 2208
rect 14296 2144 14312 2208
rect 14376 2144 14392 2208
rect 14456 2144 14472 2208
rect 14536 2144 14552 2208
rect 14616 2144 14632 2208
rect 14696 2144 14702 2208
rect 13506 2143 14702 2144
rect 1025 2138 1091 2141
rect 0 2136 1091 2138
rect 0 2080 1030 2136
rect 1086 2080 1091 2136
rect 0 2078 1091 2080
rect 0 2048 800 2078
rect 1025 2075 1091 2078
rect 0 1866 800 1896
rect 3417 1866 3483 1869
rect 0 1864 3483 1866
rect 0 1808 3422 1864
rect 3478 1808 3483 1864
rect 0 1806 3483 1808
rect 0 1776 800 1806
rect 3417 1803 3483 1806
rect 0 1594 800 1624
rect 3509 1594 3575 1597
rect 0 1592 3575 1594
rect 0 1536 3514 1592
rect 3570 1536 3575 1592
rect 0 1534 3575 1536
rect 0 1504 800 1534
rect 3509 1531 3575 1534
rect 15837 1594 15903 1597
rect 19200 1594 20000 1624
rect 15837 1592 20000 1594
rect 15837 1536 15842 1592
rect 15898 1536 20000 1592
rect 15837 1534 20000 1536
rect 15837 1531 15903 1534
rect 19200 1504 20000 1534
rect 0 1322 800 1352
rect 1117 1322 1183 1325
rect 0 1320 1183 1322
rect 0 1264 1122 1320
rect 1178 1264 1183 1320
rect 0 1262 1183 1264
rect 0 1232 800 1262
rect 1117 1259 1183 1262
rect 15377 1322 15443 1325
rect 19200 1322 20000 1352
rect 15377 1320 20000 1322
rect 15377 1264 15382 1320
rect 15438 1264 20000 1320
rect 15377 1262 20000 1264
rect 15377 1259 15443 1262
rect 19200 1232 20000 1262
rect 0 1050 800 1080
rect 3509 1050 3575 1053
rect 0 1048 3575 1050
rect 0 992 3514 1048
rect 3570 992 3575 1048
rect 0 990 3575 992
rect 0 960 800 990
rect 3509 987 3575 990
rect 19057 1050 19123 1053
rect 19200 1050 20000 1080
rect 19057 1048 20000 1050
rect 19057 992 19062 1048
rect 19118 992 20000 1048
rect 19057 990 20000 992
rect 19057 987 19123 990
rect 19200 960 20000 990
rect 0 778 800 808
rect 3325 778 3391 781
rect 0 776 3391 778
rect 0 720 3330 776
rect 3386 720 3391 776
rect 0 718 3391 720
rect 0 688 800 718
rect 3325 715 3391 718
rect 18873 778 18939 781
rect 19200 778 20000 808
rect 18873 776 20000 778
rect 18873 720 18878 776
rect 18934 720 20000 776
rect 18873 718 20000 720
rect 18873 715 18939 718
rect 19200 688 20000 718
rect 0 506 800 536
rect 3417 506 3483 509
rect 0 504 3483 506
rect 0 448 3422 504
rect 3478 448 3483 504
rect 0 446 3483 448
rect 0 416 800 446
rect 3417 443 3483 446
rect 18965 506 19031 509
rect 19200 506 20000 536
rect 18965 504 20000 506
rect 18965 448 18970 504
rect 19026 448 20000 504
rect 18965 446 20000 448
rect 18965 443 19031 446
rect 19200 416 20000 446
rect 0 234 800 264
rect 4061 234 4127 237
rect 0 232 4127 234
rect 0 176 4066 232
rect 4122 176 4127 232
rect 0 174 4127 176
rect 0 144 800 174
rect 4061 171 4127 174
rect 19057 234 19123 237
rect 19200 234 20000 264
rect 19057 232 20000 234
rect 19057 176 19062 232
rect 19118 176 20000 232
rect 19057 174 20000 176
rect 19057 171 19123 174
rect 19200 144 20000 174
<< via3 >>
rect 5512 17436 5576 17440
rect 5512 17380 5516 17436
rect 5516 17380 5572 17436
rect 5572 17380 5576 17436
rect 5512 17376 5576 17380
rect 5592 17436 5656 17440
rect 5592 17380 5596 17436
rect 5596 17380 5652 17436
rect 5652 17380 5656 17436
rect 5592 17376 5656 17380
rect 5672 17436 5736 17440
rect 5672 17380 5676 17436
rect 5676 17380 5732 17436
rect 5732 17380 5736 17436
rect 5672 17376 5736 17380
rect 5752 17436 5816 17440
rect 5752 17380 5756 17436
rect 5756 17380 5812 17436
rect 5812 17380 5816 17436
rect 5752 17376 5816 17380
rect 5832 17436 5896 17440
rect 5832 17380 5836 17436
rect 5836 17380 5892 17436
rect 5892 17380 5896 17436
rect 5832 17376 5896 17380
rect 5912 17436 5976 17440
rect 5912 17380 5916 17436
rect 5916 17380 5972 17436
rect 5972 17380 5976 17436
rect 5912 17376 5976 17380
rect 5992 17436 6056 17440
rect 5992 17380 5996 17436
rect 5996 17380 6052 17436
rect 6052 17380 6056 17436
rect 5992 17376 6056 17380
rect 6072 17436 6136 17440
rect 6072 17380 6076 17436
rect 6076 17380 6132 17436
rect 6132 17380 6136 17436
rect 6072 17376 6136 17380
rect 6152 17436 6216 17440
rect 6152 17380 6156 17436
rect 6156 17380 6212 17436
rect 6212 17380 6216 17436
rect 6152 17376 6216 17380
rect 6232 17436 6296 17440
rect 6232 17380 6236 17436
rect 6236 17380 6292 17436
rect 6292 17380 6296 17436
rect 6232 17376 6296 17380
rect 6312 17436 6376 17440
rect 6312 17380 6316 17436
rect 6316 17380 6372 17436
rect 6372 17380 6376 17436
rect 6312 17376 6376 17380
rect 6392 17436 6456 17440
rect 6392 17380 6396 17436
rect 6396 17380 6452 17436
rect 6452 17380 6456 17436
rect 6392 17376 6456 17380
rect 6472 17436 6536 17440
rect 6472 17380 6476 17436
rect 6476 17380 6532 17436
rect 6532 17380 6536 17436
rect 6472 17376 6536 17380
rect 6552 17436 6616 17440
rect 6552 17380 6556 17436
rect 6556 17380 6612 17436
rect 6612 17380 6616 17436
rect 6552 17376 6616 17380
rect 6632 17436 6696 17440
rect 6632 17380 6636 17436
rect 6636 17380 6692 17436
rect 6692 17380 6696 17436
rect 6632 17376 6696 17380
rect 13512 17436 13576 17440
rect 13512 17380 13516 17436
rect 13516 17380 13572 17436
rect 13572 17380 13576 17436
rect 13512 17376 13576 17380
rect 13592 17436 13656 17440
rect 13592 17380 13596 17436
rect 13596 17380 13652 17436
rect 13652 17380 13656 17436
rect 13592 17376 13656 17380
rect 13672 17436 13736 17440
rect 13672 17380 13676 17436
rect 13676 17380 13732 17436
rect 13732 17380 13736 17436
rect 13672 17376 13736 17380
rect 13752 17436 13816 17440
rect 13752 17380 13756 17436
rect 13756 17380 13812 17436
rect 13812 17380 13816 17436
rect 13752 17376 13816 17380
rect 13832 17436 13896 17440
rect 13832 17380 13836 17436
rect 13836 17380 13892 17436
rect 13892 17380 13896 17436
rect 13832 17376 13896 17380
rect 13912 17436 13976 17440
rect 13912 17380 13916 17436
rect 13916 17380 13972 17436
rect 13972 17380 13976 17436
rect 13912 17376 13976 17380
rect 13992 17436 14056 17440
rect 13992 17380 13996 17436
rect 13996 17380 14052 17436
rect 14052 17380 14056 17436
rect 13992 17376 14056 17380
rect 14072 17436 14136 17440
rect 14072 17380 14076 17436
rect 14076 17380 14132 17436
rect 14132 17380 14136 17436
rect 14072 17376 14136 17380
rect 14152 17436 14216 17440
rect 14152 17380 14156 17436
rect 14156 17380 14212 17436
rect 14212 17380 14216 17436
rect 14152 17376 14216 17380
rect 14232 17436 14296 17440
rect 14232 17380 14236 17436
rect 14236 17380 14292 17436
rect 14292 17380 14296 17436
rect 14232 17376 14296 17380
rect 14312 17436 14376 17440
rect 14312 17380 14316 17436
rect 14316 17380 14372 17436
rect 14372 17380 14376 17436
rect 14312 17376 14376 17380
rect 14392 17436 14456 17440
rect 14392 17380 14396 17436
rect 14396 17380 14452 17436
rect 14452 17380 14456 17436
rect 14392 17376 14456 17380
rect 14472 17436 14536 17440
rect 14472 17380 14476 17436
rect 14476 17380 14532 17436
rect 14532 17380 14536 17436
rect 14472 17376 14536 17380
rect 14552 17436 14616 17440
rect 14552 17380 14556 17436
rect 14556 17380 14612 17436
rect 14612 17380 14616 17436
rect 14552 17376 14616 17380
rect 14632 17436 14696 17440
rect 14632 17380 14636 17436
rect 14636 17380 14692 17436
rect 14692 17380 14696 17436
rect 14632 17376 14696 17380
rect 1512 16892 1576 16896
rect 1512 16836 1516 16892
rect 1516 16836 1572 16892
rect 1572 16836 1576 16892
rect 1512 16832 1576 16836
rect 1592 16892 1656 16896
rect 1592 16836 1596 16892
rect 1596 16836 1652 16892
rect 1652 16836 1656 16892
rect 1592 16832 1656 16836
rect 1672 16892 1736 16896
rect 1672 16836 1676 16892
rect 1676 16836 1732 16892
rect 1732 16836 1736 16892
rect 1672 16832 1736 16836
rect 1752 16892 1816 16896
rect 1752 16836 1756 16892
rect 1756 16836 1812 16892
rect 1812 16836 1816 16892
rect 1752 16832 1816 16836
rect 1832 16892 1896 16896
rect 1832 16836 1836 16892
rect 1836 16836 1892 16892
rect 1892 16836 1896 16892
rect 1832 16832 1896 16836
rect 1912 16892 1976 16896
rect 1912 16836 1916 16892
rect 1916 16836 1972 16892
rect 1972 16836 1976 16892
rect 1912 16832 1976 16836
rect 1992 16892 2056 16896
rect 1992 16836 1996 16892
rect 1996 16836 2052 16892
rect 2052 16836 2056 16892
rect 1992 16832 2056 16836
rect 2072 16892 2136 16896
rect 2072 16836 2076 16892
rect 2076 16836 2132 16892
rect 2132 16836 2136 16892
rect 2072 16832 2136 16836
rect 2152 16892 2216 16896
rect 2152 16836 2156 16892
rect 2156 16836 2212 16892
rect 2212 16836 2216 16892
rect 2152 16832 2216 16836
rect 2232 16892 2296 16896
rect 2232 16836 2236 16892
rect 2236 16836 2292 16892
rect 2292 16836 2296 16892
rect 2232 16832 2296 16836
rect 2312 16892 2376 16896
rect 2312 16836 2316 16892
rect 2316 16836 2372 16892
rect 2372 16836 2376 16892
rect 2312 16832 2376 16836
rect 2392 16892 2456 16896
rect 2392 16836 2396 16892
rect 2396 16836 2452 16892
rect 2452 16836 2456 16892
rect 2392 16832 2456 16836
rect 2472 16892 2536 16896
rect 2472 16836 2476 16892
rect 2476 16836 2532 16892
rect 2532 16836 2536 16892
rect 2472 16832 2536 16836
rect 2552 16892 2616 16896
rect 2552 16836 2556 16892
rect 2556 16836 2612 16892
rect 2612 16836 2616 16892
rect 2552 16832 2616 16836
rect 2632 16892 2696 16896
rect 2632 16836 2636 16892
rect 2636 16836 2692 16892
rect 2692 16836 2696 16892
rect 2632 16832 2696 16836
rect 9512 16892 9576 16896
rect 9512 16836 9516 16892
rect 9516 16836 9572 16892
rect 9572 16836 9576 16892
rect 9512 16832 9576 16836
rect 9592 16892 9656 16896
rect 9592 16836 9596 16892
rect 9596 16836 9652 16892
rect 9652 16836 9656 16892
rect 9592 16832 9656 16836
rect 9672 16892 9736 16896
rect 9672 16836 9676 16892
rect 9676 16836 9732 16892
rect 9732 16836 9736 16892
rect 9672 16832 9736 16836
rect 9752 16892 9816 16896
rect 9752 16836 9756 16892
rect 9756 16836 9812 16892
rect 9812 16836 9816 16892
rect 9752 16832 9816 16836
rect 9832 16892 9896 16896
rect 9832 16836 9836 16892
rect 9836 16836 9892 16892
rect 9892 16836 9896 16892
rect 9832 16832 9896 16836
rect 9912 16892 9976 16896
rect 9912 16836 9916 16892
rect 9916 16836 9972 16892
rect 9972 16836 9976 16892
rect 9912 16832 9976 16836
rect 9992 16892 10056 16896
rect 9992 16836 9996 16892
rect 9996 16836 10052 16892
rect 10052 16836 10056 16892
rect 9992 16832 10056 16836
rect 10072 16892 10136 16896
rect 10072 16836 10076 16892
rect 10076 16836 10132 16892
rect 10132 16836 10136 16892
rect 10072 16832 10136 16836
rect 10152 16892 10216 16896
rect 10152 16836 10156 16892
rect 10156 16836 10212 16892
rect 10212 16836 10216 16892
rect 10152 16832 10216 16836
rect 10232 16892 10296 16896
rect 10232 16836 10236 16892
rect 10236 16836 10292 16892
rect 10292 16836 10296 16892
rect 10232 16832 10296 16836
rect 10312 16892 10376 16896
rect 10312 16836 10316 16892
rect 10316 16836 10372 16892
rect 10372 16836 10376 16892
rect 10312 16832 10376 16836
rect 10392 16892 10456 16896
rect 10392 16836 10396 16892
rect 10396 16836 10452 16892
rect 10452 16836 10456 16892
rect 10392 16832 10456 16836
rect 10472 16892 10536 16896
rect 10472 16836 10476 16892
rect 10476 16836 10532 16892
rect 10532 16836 10536 16892
rect 10472 16832 10536 16836
rect 10552 16892 10616 16896
rect 10552 16836 10556 16892
rect 10556 16836 10612 16892
rect 10612 16836 10616 16892
rect 10552 16832 10616 16836
rect 10632 16892 10696 16896
rect 10632 16836 10636 16892
rect 10636 16836 10692 16892
rect 10692 16836 10696 16892
rect 10632 16832 10696 16836
rect 17512 16892 17576 16896
rect 17512 16836 17516 16892
rect 17516 16836 17572 16892
rect 17572 16836 17576 16892
rect 17512 16832 17576 16836
rect 17592 16892 17656 16896
rect 17592 16836 17596 16892
rect 17596 16836 17652 16892
rect 17652 16836 17656 16892
rect 17592 16832 17656 16836
rect 17672 16892 17736 16896
rect 17672 16836 17676 16892
rect 17676 16836 17732 16892
rect 17732 16836 17736 16892
rect 17672 16832 17736 16836
rect 17752 16892 17816 16896
rect 17752 16836 17756 16892
rect 17756 16836 17812 16892
rect 17812 16836 17816 16892
rect 17752 16832 17816 16836
rect 17832 16892 17896 16896
rect 17832 16836 17836 16892
rect 17836 16836 17892 16892
rect 17892 16836 17896 16892
rect 17832 16832 17896 16836
rect 17912 16892 17976 16896
rect 17912 16836 17916 16892
rect 17916 16836 17972 16892
rect 17972 16836 17976 16892
rect 17912 16832 17976 16836
rect 17992 16892 18056 16896
rect 17992 16836 17996 16892
rect 17996 16836 18052 16892
rect 18052 16836 18056 16892
rect 17992 16832 18056 16836
rect 18072 16892 18136 16896
rect 18072 16836 18076 16892
rect 18076 16836 18132 16892
rect 18132 16836 18136 16892
rect 18072 16832 18136 16836
rect 18152 16892 18216 16896
rect 18152 16836 18156 16892
rect 18156 16836 18212 16892
rect 18212 16836 18216 16892
rect 18152 16832 18216 16836
rect 18232 16892 18296 16896
rect 18232 16836 18236 16892
rect 18236 16836 18292 16892
rect 18292 16836 18296 16892
rect 18232 16832 18296 16836
rect 18312 16892 18376 16896
rect 18312 16836 18316 16892
rect 18316 16836 18372 16892
rect 18372 16836 18376 16892
rect 18312 16832 18376 16836
rect 18392 16892 18456 16896
rect 18392 16836 18396 16892
rect 18396 16836 18452 16892
rect 18452 16836 18456 16892
rect 18392 16832 18456 16836
rect 18472 16892 18536 16896
rect 18472 16836 18476 16892
rect 18476 16836 18532 16892
rect 18532 16836 18536 16892
rect 18472 16832 18536 16836
rect 18552 16892 18616 16896
rect 18552 16836 18556 16892
rect 18556 16836 18612 16892
rect 18612 16836 18616 16892
rect 18552 16832 18616 16836
rect 18632 16892 18696 16896
rect 18632 16836 18636 16892
rect 18636 16836 18692 16892
rect 18692 16836 18696 16892
rect 18632 16832 18696 16836
rect 5512 16348 5576 16352
rect 5512 16292 5516 16348
rect 5516 16292 5572 16348
rect 5572 16292 5576 16348
rect 5512 16288 5576 16292
rect 5592 16348 5656 16352
rect 5592 16292 5596 16348
rect 5596 16292 5652 16348
rect 5652 16292 5656 16348
rect 5592 16288 5656 16292
rect 5672 16348 5736 16352
rect 5672 16292 5676 16348
rect 5676 16292 5732 16348
rect 5732 16292 5736 16348
rect 5672 16288 5736 16292
rect 5752 16348 5816 16352
rect 5752 16292 5756 16348
rect 5756 16292 5812 16348
rect 5812 16292 5816 16348
rect 5752 16288 5816 16292
rect 5832 16348 5896 16352
rect 5832 16292 5836 16348
rect 5836 16292 5892 16348
rect 5892 16292 5896 16348
rect 5832 16288 5896 16292
rect 5912 16348 5976 16352
rect 5912 16292 5916 16348
rect 5916 16292 5972 16348
rect 5972 16292 5976 16348
rect 5912 16288 5976 16292
rect 5992 16348 6056 16352
rect 5992 16292 5996 16348
rect 5996 16292 6052 16348
rect 6052 16292 6056 16348
rect 5992 16288 6056 16292
rect 6072 16348 6136 16352
rect 6072 16292 6076 16348
rect 6076 16292 6132 16348
rect 6132 16292 6136 16348
rect 6072 16288 6136 16292
rect 6152 16348 6216 16352
rect 6152 16292 6156 16348
rect 6156 16292 6212 16348
rect 6212 16292 6216 16348
rect 6152 16288 6216 16292
rect 6232 16348 6296 16352
rect 6232 16292 6236 16348
rect 6236 16292 6292 16348
rect 6292 16292 6296 16348
rect 6232 16288 6296 16292
rect 6312 16348 6376 16352
rect 6312 16292 6316 16348
rect 6316 16292 6372 16348
rect 6372 16292 6376 16348
rect 6312 16288 6376 16292
rect 6392 16348 6456 16352
rect 6392 16292 6396 16348
rect 6396 16292 6452 16348
rect 6452 16292 6456 16348
rect 6392 16288 6456 16292
rect 6472 16348 6536 16352
rect 6472 16292 6476 16348
rect 6476 16292 6532 16348
rect 6532 16292 6536 16348
rect 6472 16288 6536 16292
rect 6552 16348 6616 16352
rect 6552 16292 6556 16348
rect 6556 16292 6612 16348
rect 6612 16292 6616 16348
rect 6552 16288 6616 16292
rect 6632 16348 6696 16352
rect 6632 16292 6636 16348
rect 6636 16292 6692 16348
rect 6692 16292 6696 16348
rect 6632 16288 6696 16292
rect 13512 16348 13576 16352
rect 13512 16292 13516 16348
rect 13516 16292 13572 16348
rect 13572 16292 13576 16348
rect 13512 16288 13576 16292
rect 13592 16348 13656 16352
rect 13592 16292 13596 16348
rect 13596 16292 13652 16348
rect 13652 16292 13656 16348
rect 13592 16288 13656 16292
rect 13672 16348 13736 16352
rect 13672 16292 13676 16348
rect 13676 16292 13732 16348
rect 13732 16292 13736 16348
rect 13672 16288 13736 16292
rect 13752 16348 13816 16352
rect 13752 16292 13756 16348
rect 13756 16292 13812 16348
rect 13812 16292 13816 16348
rect 13752 16288 13816 16292
rect 13832 16348 13896 16352
rect 13832 16292 13836 16348
rect 13836 16292 13892 16348
rect 13892 16292 13896 16348
rect 13832 16288 13896 16292
rect 13912 16348 13976 16352
rect 13912 16292 13916 16348
rect 13916 16292 13972 16348
rect 13972 16292 13976 16348
rect 13912 16288 13976 16292
rect 13992 16348 14056 16352
rect 13992 16292 13996 16348
rect 13996 16292 14052 16348
rect 14052 16292 14056 16348
rect 13992 16288 14056 16292
rect 14072 16348 14136 16352
rect 14072 16292 14076 16348
rect 14076 16292 14132 16348
rect 14132 16292 14136 16348
rect 14072 16288 14136 16292
rect 14152 16348 14216 16352
rect 14152 16292 14156 16348
rect 14156 16292 14212 16348
rect 14212 16292 14216 16348
rect 14152 16288 14216 16292
rect 14232 16348 14296 16352
rect 14232 16292 14236 16348
rect 14236 16292 14292 16348
rect 14292 16292 14296 16348
rect 14232 16288 14296 16292
rect 14312 16348 14376 16352
rect 14312 16292 14316 16348
rect 14316 16292 14372 16348
rect 14372 16292 14376 16348
rect 14312 16288 14376 16292
rect 14392 16348 14456 16352
rect 14392 16292 14396 16348
rect 14396 16292 14452 16348
rect 14452 16292 14456 16348
rect 14392 16288 14456 16292
rect 14472 16348 14536 16352
rect 14472 16292 14476 16348
rect 14476 16292 14532 16348
rect 14532 16292 14536 16348
rect 14472 16288 14536 16292
rect 14552 16348 14616 16352
rect 14552 16292 14556 16348
rect 14556 16292 14612 16348
rect 14612 16292 14616 16348
rect 14552 16288 14616 16292
rect 14632 16348 14696 16352
rect 14632 16292 14636 16348
rect 14636 16292 14692 16348
rect 14692 16292 14696 16348
rect 14632 16288 14696 16292
rect 1512 15804 1576 15808
rect 1512 15748 1516 15804
rect 1516 15748 1572 15804
rect 1572 15748 1576 15804
rect 1512 15744 1576 15748
rect 1592 15804 1656 15808
rect 1592 15748 1596 15804
rect 1596 15748 1652 15804
rect 1652 15748 1656 15804
rect 1592 15744 1656 15748
rect 1672 15804 1736 15808
rect 1672 15748 1676 15804
rect 1676 15748 1732 15804
rect 1732 15748 1736 15804
rect 1672 15744 1736 15748
rect 1752 15804 1816 15808
rect 1752 15748 1756 15804
rect 1756 15748 1812 15804
rect 1812 15748 1816 15804
rect 1752 15744 1816 15748
rect 1832 15804 1896 15808
rect 1832 15748 1836 15804
rect 1836 15748 1892 15804
rect 1892 15748 1896 15804
rect 1832 15744 1896 15748
rect 1912 15804 1976 15808
rect 1912 15748 1916 15804
rect 1916 15748 1972 15804
rect 1972 15748 1976 15804
rect 1912 15744 1976 15748
rect 1992 15804 2056 15808
rect 1992 15748 1996 15804
rect 1996 15748 2052 15804
rect 2052 15748 2056 15804
rect 1992 15744 2056 15748
rect 2072 15804 2136 15808
rect 2072 15748 2076 15804
rect 2076 15748 2132 15804
rect 2132 15748 2136 15804
rect 2072 15744 2136 15748
rect 2152 15804 2216 15808
rect 2152 15748 2156 15804
rect 2156 15748 2212 15804
rect 2212 15748 2216 15804
rect 2152 15744 2216 15748
rect 2232 15804 2296 15808
rect 2232 15748 2236 15804
rect 2236 15748 2292 15804
rect 2292 15748 2296 15804
rect 2232 15744 2296 15748
rect 2312 15804 2376 15808
rect 2312 15748 2316 15804
rect 2316 15748 2372 15804
rect 2372 15748 2376 15804
rect 2312 15744 2376 15748
rect 2392 15804 2456 15808
rect 2392 15748 2396 15804
rect 2396 15748 2452 15804
rect 2452 15748 2456 15804
rect 2392 15744 2456 15748
rect 2472 15804 2536 15808
rect 2472 15748 2476 15804
rect 2476 15748 2532 15804
rect 2532 15748 2536 15804
rect 2472 15744 2536 15748
rect 2552 15804 2616 15808
rect 2552 15748 2556 15804
rect 2556 15748 2612 15804
rect 2612 15748 2616 15804
rect 2552 15744 2616 15748
rect 2632 15804 2696 15808
rect 2632 15748 2636 15804
rect 2636 15748 2692 15804
rect 2692 15748 2696 15804
rect 2632 15744 2696 15748
rect 9512 15804 9576 15808
rect 9512 15748 9516 15804
rect 9516 15748 9572 15804
rect 9572 15748 9576 15804
rect 9512 15744 9576 15748
rect 9592 15804 9656 15808
rect 9592 15748 9596 15804
rect 9596 15748 9652 15804
rect 9652 15748 9656 15804
rect 9592 15744 9656 15748
rect 9672 15804 9736 15808
rect 9672 15748 9676 15804
rect 9676 15748 9732 15804
rect 9732 15748 9736 15804
rect 9672 15744 9736 15748
rect 9752 15804 9816 15808
rect 9752 15748 9756 15804
rect 9756 15748 9812 15804
rect 9812 15748 9816 15804
rect 9752 15744 9816 15748
rect 9832 15804 9896 15808
rect 9832 15748 9836 15804
rect 9836 15748 9892 15804
rect 9892 15748 9896 15804
rect 9832 15744 9896 15748
rect 9912 15804 9976 15808
rect 9912 15748 9916 15804
rect 9916 15748 9972 15804
rect 9972 15748 9976 15804
rect 9912 15744 9976 15748
rect 9992 15804 10056 15808
rect 9992 15748 9996 15804
rect 9996 15748 10052 15804
rect 10052 15748 10056 15804
rect 9992 15744 10056 15748
rect 10072 15804 10136 15808
rect 10072 15748 10076 15804
rect 10076 15748 10132 15804
rect 10132 15748 10136 15804
rect 10072 15744 10136 15748
rect 10152 15804 10216 15808
rect 10152 15748 10156 15804
rect 10156 15748 10212 15804
rect 10212 15748 10216 15804
rect 10152 15744 10216 15748
rect 10232 15804 10296 15808
rect 10232 15748 10236 15804
rect 10236 15748 10292 15804
rect 10292 15748 10296 15804
rect 10232 15744 10296 15748
rect 10312 15804 10376 15808
rect 10312 15748 10316 15804
rect 10316 15748 10372 15804
rect 10372 15748 10376 15804
rect 10312 15744 10376 15748
rect 10392 15804 10456 15808
rect 10392 15748 10396 15804
rect 10396 15748 10452 15804
rect 10452 15748 10456 15804
rect 10392 15744 10456 15748
rect 10472 15804 10536 15808
rect 10472 15748 10476 15804
rect 10476 15748 10532 15804
rect 10532 15748 10536 15804
rect 10472 15744 10536 15748
rect 10552 15804 10616 15808
rect 10552 15748 10556 15804
rect 10556 15748 10612 15804
rect 10612 15748 10616 15804
rect 10552 15744 10616 15748
rect 10632 15804 10696 15808
rect 10632 15748 10636 15804
rect 10636 15748 10692 15804
rect 10692 15748 10696 15804
rect 10632 15744 10696 15748
rect 17512 15804 17576 15808
rect 17512 15748 17516 15804
rect 17516 15748 17572 15804
rect 17572 15748 17576 15804
rect 17512 15744 17576 15748
rect 17592 15804 17656 15808
rect 17592 15748 17596 15804
rect 17596 15748 17652 15804
rect 17652 15748 17656 15804
rect 17592 15744 17656 15748
rect 17672 15804 17736 15808
rect 17672 15748 17676 15804
rect 17676 15748 17732 15804
rect 17732 15748 17736 15804
rect 17672 15744 17736 15748
rect 17752 15804 17816 15808
rect 17752 15748 17756 15804
rect 17756 15748 17812 15804
rect 17812 15748 17816 15804
rect 17752 15744 17816 15748
rect 17832 15804 17896 15808
rect 17832 15748 17836 15804
rect 17836 15748 17892 15804
rect 17892 15748 17896 15804
rect 17832 15744 17896 15748
rect 17912 15804 17976 15808
rect 17912 15748 17916 15804
rect 17916 15748 17972 15804
rect 17972 15748 17976 15804
rect 17912 15744 17976 15748
rect 17992 15804 18056 15808
rect 17992 15748 17996 15804
rect 17996 15748 18052 15804
rect 18052 15748 18056 15804
rect 17992 15744 18056 15748
rect 18072 15804 18136 15808
rect 18072 15748 18076 15804
rect 18076 15748 18132 15804
rect 18132 15748 18136 15804
rect 18072 15744 18136 15748
rect 18152 15804 18216 15808
rect 18152 15748 18156 15804
rect 18156 15748 18212 15804
rect 18212 15748 18216 15804
rect 18152 15744 18216 15748
rect 18232 15804 18296 15808
rect 18232 15748 18236 15804
rect 18236 15748 18292 15804
rect 18292 15748 18296 15804
rect 18232 15744 18296 15748
rect 18312 15804 18376 15808
rect 18312 15748 18316 15804
rect 18316 15748 18372 15804
rect 18372 15748 18376 15804
rect 18312 15744 18376 15748
rect 18392 15804 18456 15808
rect 18392 15748 18396 15804
rect 18396 15748 18452 15804
rect 18452 15748 18456 15804
rect 18392 15744 18456 15748
rect 18472 15804 18536 15808
rect 18472 15748 18476 15804
rect 18476 15748 18532 15804
rect 18532 15748 18536 15804
rect 18472 15744 18536 15748
rect 18552 15804 18616 15808
rect 18552 15748 18556 15804
rect 18556 15748 18612 15804
rect 18612 15748 18616 15804
rect 18552 15744 18616 15748
rect 18632 15804 18696 15808
rect 18632 15748 18636 15804
rect 18636 15748 18692 15804
rect 18692 15748 18696 15804
rect 18632 15744 18696 15748
rect 5512 15260 5576 15264
rect 5512 15204 5516 15260
rect 5516 15204 5572 15260
rect 5572 15204 5576 15260
rect 5512 15200 5576 15204
rect 5592 15260 5656 15264
rect 5592 15204 5596 15260
rect 5596 15204 5652 15260
rect 5652 15204 5656 15260
rect 5592 15200 5656 15204
rect 5672 15260 5736 15264
rect 5672 15204 5676 15260
rect 5676 15204 5732 15260
rect 5732 15204 5736 15260
rect 5672 15200 5736 15204
rect 5752 15260 5816 15264
rect 5752 15204 5756 15260
rect 5756 15204 5812 15260
rect 5812 15204 5816 15260
rect 5752 15200 5816 15204
rect 5832 15260 5896 15264
rect 5832 15204 5836 15260
rect 5836 15204 5892 15260
rect 5892 15204 5896 15260
rect 5832 15200 5896 15204
rect 5912 15260 5976 15264
rect 5912 15204 5916 15260
rect 5916 15204 5972 15260
rect 5972 15204 5976 15260
rect 5912 15200 5976 15204
rect 5992 15260 6056 15264
rect 5992 15204 5996 15260
rect 5996 15204 6052 15260
rect 6052 15204 6056 15260
rect 5992 15200 6056 15204
rect 6072 15260 6136 15264
rect 6072 15204 6076 15260
rect 6076 15204 6132 15260
rect 6132 15204 6136 15260
rect 6072 15200 6136 15204
rect 6152 15260 6216 15264
rect 6152 15204 6156 15260
rect 6156 15204 6212 15260
rect 6212 15204 6216 15260
rect 6152 15200 6216 15204
rect 6232 15260 6296 15264
rect 6232 15204 6236 15260
rect 6236 15204 6292 15260
rect 6292 15204 6296 15260
rect 6232 15200 6296 15204
rect 6312 15260 6376 15264
rect 6312 15204 6316 15260
rect 6316 15204 6372 15260
rect 6372 15204 6376 15260
rect 6312 15200 6376 15204
rect 6392 15260 6456 15264
rect 6392 15204 6396 15260
rect 6396 15204 6452 15260
rect 6452 15204 6456 15260
rect 6392 15200 6456 15204
rect 6472 15260 6536 15264
rect 6472 15204 6476 15260
rect 6476 15204 6532 15260
rect 6532 15204 6536 15260
rect 6472 15200 6536 15204
rect 6552 15260 6616 15264
rect 6552 15204 6556 15260
rect 6556 15204 6612 15260
rect 6612 15204 6616 15260
rect 6552 15200 6616 15204
rect 6632 15260 6696 15264
rect 6632 15204 6636 15260
rect 6636 15204 6692 15260
rect 6692 15204 6696 15260
rect 6632 15200 6696 15204
rect 13512 15260 13576 15264
rect 13512 15204 13516 15260
rect 13516 15204 13572 15260
rect 13572 15204 13576 15260
rect 13512 15200 13576 15204
rect 13592 15260 13656 15264
rect 13592 15204 13596 15260
rect 13596 15204 13652 15260
rect 13652 15204 13656 15260
rect 13592 15200 13656 15204
rect 13672 15260 13736 15264
rect 13672 15204 13676 15260
rect 13676 15204 13732 15260
rect 13732 15204 13736 15260
rect 13672 15200 13736 15204
rect 13752 15260 13816 15264
rect 13752 15204 13756 15260
rect 13756 15204 13812 15260
rect 13812 15204 13816 15260
rect 13752 15200 13816 15204
rect 13832 15260 13896 15264
rect 13832 15204 13836 15260
rect 13836 15204 13892 15260
rect 13892 15204 13896 15260
rect 13832 15200 13896 15204
rect 13912 15260 13976 15264
rect 13912 15204 13916 15260
rect 13916 15204 13972 15260
rect 13972 15204 13976 15260
rect 13912 15200 13976 15204
rect 13992 15260 14056 15264
rect 13992 15204 13996 15260
rect 13996 15204 14052 15260
rect 14052 15204 14056 15260
rect 13992 15200 14056 15204
rect 14072 15260 14136 15264
rect 14072 15204 14076 15260
rect 14076 15204 14132 15260
rect 14132 15204 14136 15260
rect 14072 15200 14136 15204
rect 14152 15260 14216 15264
rect 14152 15204 14156 15260
rect 14156 15204 14212 15260
rect 14212 15204 14216 15260
rect 14152 15200 14216 15204
rect 14232 15260 14296 15264
rect 14232 15204 14236 15260
rect 14236 15204 14292 15260
rect 14292 15204 14296 15260
rect 14232 15200 14296 15204
rect 14312 15260 14376 15264
rect 14312 15204 14316 15260
rect 14316 15204 14372 15260
rect 14372 15204 14376 15260
rect 14312 15200 14376 15204
rect 14392 15260 14456 15264
rect 14392 15204 14396 15260
rect 14396 15204 14452 15260
rect 14452 15204 14456 15260
rect 14392 15200 14456 15204
rect 14472 15260 14536 15264
rect 14472 15204 14476 15260
rect 14476 15204 14532 15260
rect 14532 15204 14536 15260
rect 14472 15200 14536 15204
rect 14552 15260 14616 15264
rect 14552 15204 14556 15260
rect 14556 15204 14612 15260
rect 14612 15204 14616 15260
rect 14552 15200 14616 15204
rect 14632 15260 14696 15264
rect 14632 15204 14636 15260
rect 14636 15204 14692 15260
rect 14692 15204 14696 15260
rect 14632 15200 14696 15204
rect 1512 14716 1576 14720
rect 1512 14660 1516 14716
rect 1516 14660 1572 14716
rect 1572 14660 1576 14716
rect 1512 14656 1576 14660
rect 1592 14716 1656 14720
rect 1592 14660 1596 14716
rect 1596 14660 1652 14716
rect 1652 14660 1656 14716
rect 1592 14656 1656 14660
rect 1672 14716 1736 14720
rect 1672 14660 1676 14716
rect 1676 14660 1732 14716
rect 1732 14660 1736 14716
rect 1672 14656 1736 14660
rect 1752 14716 1816 14720
rect 1752 14660 1756 14716
rect 1756 14660 1812 14716
rect 1812 14660 1816 14716
rect 1752 14656 1816 14660
rect 1832 14716 1896 14720
rect 1832 14660 1836 14716
rect 1836 14660 1892 14716
rect 1892 14660 1896 14716
rect 1832 14656 1896 14660
rect 1912 14716 1976 14720
rect 1912 14660 1916 14716
rect 1916 14660 1972 14716
rect 1972 14660 1976 14716
rect 1912 14656 1976 14660
rect 1992 14716 2056 14720
rect 1992 14660 1996 14716
rect 1996 14660 2052 14716
rect 2052 14660 2056 14716
rect 1992 14656 2056 14660
rect 2072 14716 2136 14720
rect 2072 14660 2076 14716
rect 2076 14660 2132 14716
rect 2132 14660 2136 14716
rect 2072 14656 2136 14660
rect 2152 14716 2216 14720
rect 2152 14660 2156 14716
rect 2156 14660 2212 14716
rect 2212 14660 2216 14716
rect 2152 14656 2216 14660
rect 2232 14716 2296 14720
rect 2232 14660 2236 14716
rect 2236 14660 2292 14716
rect 2292 14660 2296 14716
rect 2232 14656 2296 14660
rect 2312 14716 2376 14720
rect 2312 14660 2316 14716
rect 2316 14660 2372 14716
rect 2372 14660 2376 14716
rect 2312 14656 2376 14660
rect 2392 14716 2456 14720
rect 2392 14660 2396 14716
rect 2396 14660 2452 14716
rect 2452 14660 2456 14716
rect 2392 14656 2456 14660
rect 2472 14716 2536 14720
rect 2472 14660 2476 14716
rect 2476 14660 2532 14716
rect 2532 14660 2536 14716
rect 2472 14656 2536 14660
rect 2552 14716 2616 14720
rect 2552 14660 2556 14716
rect 2556 14660 2612 14716
rect 2612 14660 2616 14716
rect 2552 14656 2616 14660
rect 2632 14716 2696 14720
rect 2632 14660 2636 14716
rect 2636 14660 2692 14716
rect 2692 14660 2696 14716
rect 2632 14656 2696 14660
rect 9512 14716 9576 14720
rect 9512 14660 9516 14716
rect 9516 14660 9572 14716
rect 9572 14660 9576 14716
rect 9512 14656 9576 14660
rect 9592 14716 9656 14720
rect 9592 14660 9596 14716
rect 9596 14660 9652 14716
rect 9652 14660 9656 14716
rect 9592 14656 9656 14660
rect 9672 14716 9736 14720
rect 9672 14660 9676 14716
rect 9676 14660 9732 14716
rect 9732 14660 9736 14716
rect 9672 14656 9736 14660
rect 9752 14716 9816 14720
rect 9752 14660 9756 14716
rect 9756 14660 9812 14716
rect 9812 14660 9816 14716
rect 9752 14656 9816 14660
rect 9832 14716 9896 14720
rect 9832 14660 9836 14716
rect 9836 14660 9892 14716
rect 9892 14660 9896 14716
rect 9832 14656 9896 14660
rect 9912 14716 9976 14720
rect 9912 14660 9916 14716
rect 9916 14660 9972 14716
rect 9972 14660 9976 14716
rect 9912 14656 9976 14660
rect 9992 14716 10056 14720
rect 9992 14660 9996 14716
rect 9996 14660 10052 14716
rect 10052 14660 10056 14716
rect 9992 14656 10056 14660
rect 10072 14716 10136 14720
rect 10072 14660 10076 14716
rect 10076 14660 10132 14716
rect 10132 14660 10136 14716
rect 10072 14656 10136 14660
rect 10152 14716 10216 14720
rect 10152 14660 10156 14716
rect 10156 14660 10212 14716
rect 10212 14660 10216 14716
rect 10152 14656 10216 14660
rect 10232 14716 10296 14720
rect 10232 14660 10236 14716
rect 10236 14660 10292 14716
rect 10292 14660 10296 14716
rect 10232 14656 10296 14660
rect 10312 14716 10376 14720
rect 10312 14660 10316 14716
rect 10316 14660 10372 14716
rect 10372 14660 10376 14716
rect 10312 14656 10376 14660
rect 10392 14716 10456 14720
rect 10392 14660 10396 14716
rect 10396 14660 10452 14716
rect 10452 14660 10456 14716
rect 10392 14656 10456 14660
rect 10472 14716 10536 14720
rect 10472 14660 10476 14716
rect 10476 14660 10532 14716
rect 10532 14660 10536 14716
rect 10472 14656 10536 14660
rect 10552 14716 10616 14720
rect 10552 14660 10556 14716
rect 10556 14660 10612 14716
rect 10612 14660 10616 14716
rect 10552 14656 10616 14660
rect 10632 14716 10696 14720
rect 10632 14660 10636 14716
rect 10636 14660 10692 14716
rect 10692 14660 10696 14716
rect 10632 14656 10696 14660
rect 17512 14716 17576 14720
rect 17512 14660 17516 14716
rect 17516 14660 17572 14716
rect 17572 14660 17576 14716
rect 17512 14656 17576 14660
rect 17592 14716 17656 14720
rect 17592 14660 17596 14716
rect 17596 14660 17652 14716
rect 17652 14660 17656 14716
rect 17592 14656 17656 14660
rect 17672 14716 17736 14720
rect 17672 14660 17676 14716
rect 17676 14660 17732 14716
rect 17732 14660 17736 14716
rect 17672 14656 17736 14660
rect 17752 14716 17816 14720
rect 17752 14660 17756 14716
rect 17756 14660 17812 14716
rect 17812 14660 17816 14716
rect 17752 14656 17816 14660
rect 17832 14716 17896 14720
rect 17832 14660 17836 14716
rect 17836 14660 17892 14716
rect 17892 14660 17896 14716
rect 17832 14656 17896 14660
rect 17912 14716 17976 14720
rect 17912 14660 17916 14716
rect 17916 14660 17972 14716
rect 17972 14660 17976 14716
rect 17912 14656 17976 14660
rect 17992 14716 18056 14720
rect 17992 14660 17996 14716
rect 17996 14660 18052 14716
rect 18052 14660 18056 14716
rect 17992 14656 18056 14660
rect 18072 14716 18136 14720
rect 18072 14660 18076 14716
rect 18076 14660 18132 14716
rect 18132 14660 18136 14716
rect 18072 14656 18136 14660
rect 18152 14716 18216 14720
rect 18152 14660 18156 14716
rect 18156 14660 18212 14716
rect 18212 14660 18216 14716
rect 18152 14656 18216 14660
rect 18232 14716 18296 14720
rect 18232 14660 18236 14716
rect 18236 14660 18292 14716
rect 18292 14660 18296 14716
rect 18232 14656 18296 14660
rect 18312 14716 18376 14720
rect 18312 14660 18316 14716
rect 18316 14660 18372 14716
rect 18372 14660 18376 14716
rect 18312 14656 18376 14660
rect 18392 14716 18456 14720
rect 18392 14660 18396 14716
rect 18396 14660 18452 14716
rect 18452 14660 18456 14716
rect 18392 14656 18456 14660
rect 18472 14716 18536 14720
rect 18472 14660 18476 14716
rect 18476 14660 18532 14716
rect 18532 14660 18536 14716
rect 18472 14656 18536 14660
rect 18552 14716 18616 14720
rect 18552 14660 18556 14716
rect 18556 14660 18612 14716
rect 18612 14660 18616 14716
rect 18552 14656 18616 14660
rect 18632 14716 18696 14720
rect 18632 14660 18636 14716
rect 18636 14660 18692 14716
rect 18692 14660 18696 14716
rect 18632 14656 18696 14660
rect 1512 13628 1576 13632
rect 1512 13572 1516 13628
rect 1516 13572 1572 13628
rect 1572 13572 1576 13628
rect 1512 13568 1576 13572
rect 1592 13628 1656 13632
rect 1592 13572 1596 13628
rect 1596 13572 1652 13628
rect 1652 13572 1656 13628
rect 1592 13568 1656 13572
rect 1672 13628 1736 13632
rect 1672 13572 1676 13628
rect 1676 13572 1732 13628
rect 1732 13572 1736 13628
rect 1672 13568 1736 13572
rect 1752 13628 1816 13632
rect 1752 13572 1756 13628
rect 1756 13572 1812 13628
rect 1812 13572 1816 13628
rect 1752 13568 1816 13572
rect 1832 13628 1896 13632
rect 1832 13572 1836 13628
rect 1836 13572 1892 13628
rect 1892 13572 1896 13628
rect 1832 13568 1896 13572
rect 1912 13628 1976 13632
rect 1912 13572 1916 13628
rect 1916 13572 1972 13628
rect 1972 13572 1976 13628
rect 1912 13568 1976 13572
rect 1992 13628 2056 13632
rect 1992 13572 1996 13628
rect 1996 13572 2052 13628
rect 2052 13572 2056 13628
rect 1992 13568 2056 13572
rect 2072 13628 2136 13632
rect 2072 13572 2076 13628
rect 2076 13572 2132 13628
rect 2132 13572 2136 13628
rect 2072 13568 2136 13572
rect 2152 13628 2216 13632
rect 2152 13572 2156 13628
rect 2156 13572 2212 13628
rect 2212 13572 2216 13628
rect 2152 13568 2216 13572
rect 2232 13628 2296 13632
rect 2232 13572 2236 13628
rect 2236 13572 2292 13628
rect 2292 13572 2296 13628
rect 2232 13568 2296 13572
rect 2312 13628 2376 13632
rect 2312 13572 2316 13628
rect 2316 13572 2372 13628
rect 2372 13572 2376 13628
rect 2312 13568 2376 13572
rect 2392 13628 2456 13632
rect 2392 13572 2396 13628
rect 2396 13572 2452 13628
rect 2452 13572 2456 13628
rect 2392 13568 2456 13572
rect 2472 13628 2536 13632
rect 2472 13572 2476 13628
rect 2476 13572 2532 13628
rect 2532 13572 2536 13628
rect 2472 13568 2536 13572
rect 2552 13628 2616 13632
rect 2552 13572 2556 13628
rect 2556 13572 2612 13628
rect 2612 13572 2616 13628
rect 2552 13568 2616 13572
rect 2632 13628 2696 13632
rect 2632 13572 2636 13628
rect 2636 13572 2692 13628
rect 2692 13572 2696 13628
rect 2632 13568 2696 13572
rect 5512 14172 5576 14176
rect 5512 14116 5516 14172
rect 5516 14116 5572 14172
rect 5572 14116 5576 14172
rect 5512 14112 5576 14116
rect 5592 14172 5656 14176
rect 5592 14116 5596 14172
rect 5596 14116 5652 14172
rect 5652 14116 5656 14172
rect 5592 14112 5656 14116
rect 5672 14172 5736 14176
rect 5672 14116 5676 14172
rect 5676 14116 5732 14172
rect 5732 14116 5736 14172
rect 5672 14112 5736 14116
rect 5752 14172 5816 14176
rect 5752 14116 5756 14172
rect 5756 14116 5812 14172
rect 5812 14116 5816 14172
rect 5752 14112 5816 14116
rect 5832 14172 5896 14176
rect 5832 14116 5836 14172
rect 5836 14116 5892 14172
rect 5892 14116 5896 14172
rect 5832 14112 5896 14116
rect 5912 14172 5976 14176
rect 5912 14116 5916 14172
rect 5916 14116 5972 14172
rect 5972 14116 5976 14172
rect 5912 14112 5976 14116
rect 5992 14172 6056 14176
rect 5992 14116 5996 14172
rect 5996 14116 6052 14172
rect 6052 14116 6056 14172
rect 5992 14112 6056 14116
rect 6072 14172 6136 14176
rect 6072 14116 6076 14172
rect 6076 14116 6132 14172
rect 6132 14116 6136 14172
rect 6072 14112 6136 14116
rect 6152 14172 6216 14176
rect 6152 14116 6156 14172
rect 6156 14116 6212 14172
rect 6212 14116 6216 14172
rect 6152 14112 6216 14116
rect 6232 14172 6296 14176
rect 6232 14116 6236 14172
rect 6236 14116 6292 14172
rect 6292 14116 6296 14172
rect 6232 14112 6296 14116
rect 6312 14172 6376 14176
rect 6312 14116 6316 14172
rect 6316 14116 6372 14172
rect 6372 14116 6376 14172
rect 6312 14112 6376 14116
rect 6392 14172 6456 14176
rect 6392 14116 6396 14172
rect 6396 14116 6452 14172
rect 6452 14116 6456 14172
rect 6392 14112 6456 14116
rect 6472 14172 6536 14176
rect 6472 14116 6476 14172
rect 6476 14116 6532 14172
rect 6532 14116 6536 14172
rect 6472 14112 6536 14116
rect 6552 14172 6616 14176
rect 6552 14116 6556 14172
rect 6556 14116 6612 14172
rect 6612 14116 6616 14172
rect 6552 14112 6616 14116
rect 6632 14172 6696 14176
rect 6632 14116 6636 14172
rect 6636 14116 6692 14172
rect 6692 14116 6696 14172
rect 6632 14112 6696 14116
rect 13512 14172 13576 14176
rect 13512 14116 13516 14172
rect 13516 14116 13572 14172
rect 13572 14116 13576 14172
rect 13512 14112 13576 14116
rect 13592 14172 13656 14176
rect 13592 14116 13596 14172
rect 13596 14116 13652 14172
rect 13652 14116 13656 14172
rect 13592 14112 13656 14116
rect 13672 14172 13736 14176
rect 13672 14116 13676 14172
rect 13676 14116 13732 14172
rect 13732 14116 13736 14172
rect 13672 14112 13736 14116
rect 13752 14172 13816 14176
rect 13752 14116 13756 14172
rect 13756 14116 13812 14172
rect 13812 14116 13816 14172
rect 13752 14112 13816 14116
rect 13832 14172 13896 14176
rect 13832 14116 13836 14172
rect 13836 14116 13892 14172
rect 13892 14116 13896 14172
rect 13832 14112 13896 14116
rect 13912 14172 13976 14176
rect 13912 14116 13916 14172
rect 13916 14116 13972 14172
rect 13972 14116 13976 14172
rect 13912 14112 13976 14116
rect 13992 14172 14056 14176
rect 13992 14116 13996 14172
rect 13996 14116 14052 14172
rect 14052 14116 14056 14172
rect 13992 14112 14056 14116
rect 14072 14172 14136 14176
rect 14072 14116 14076 14172
rect 14076 14116 14132 14172
rect 14132 14116 14136 14172
rect 14072 14112 14136 14116
rect 14152 14172 14216 14176
rect 14152 14116 14156 14172
rect 14156 14116 14212 14172
rect 14212 14116 14216 14172
rect 14152 14112 14216 14116
rect 14232 14172 14296 14176
rect 14232 14116 14236 14172
rect 14236 14116 14292 14172
rect 14292 14116 14296 14172
rect 14232 14112 14296 14116
rect 14312 14172 14376 14176
rect 14312 14116 14316 14172
rect 14316 14116 14372 14172
rect 14372 14116 14376 14172
rect 14312 14112 14376 14116
rect 14392 14172 14456 14176
rect 14392 14116 14396 14172
rect 14396 14116 14452 14172
rect 14452 14116 14456 14172
rect 14392 14112 14456 14116
rect 14472 14172 14536 14176
rect 14472 14116 14476 14172
rect 14476 14116 14532 14172
rect 14532 14116 14536 14172
rect 14472 14112 14536 14116
rect 14552 14172 14616 14176
rect 14552 14116 14556 14172
rect 14556 14116 14612 14172
rect 14612 14116 14616 14172
rect 14552 14112 14616 14116
rect 14632 14172 14696 14176
rect 14632 14116 14636 14172
rect 14636 14116 14692 14172
rect 14692 14116 14696 14172
rect 14632 14112 14696 14116
rect 1512 12540 1576 12544
rect 1512 12484 1516 12540
rect 1516 12484 1572 12540
rect 1572 12484 1576 12540
rect 1512 12480 1576 12484
rect 1592 12540 1656 12544
rect 1592 12484 1596 12540
rect 1596 12484 1652 12540
rect 1652 12484 1656 12540
rect 1592 12480 1656 12484
rect 1672 12540 1736 12544
rect 1672 12484 1676 12540
rect 1676 12484 1732 12540
rect 1732 12484 1736 12540
rect 1672 12480 1736 12484
rect 1752 12540 1816 12544
rect 1752 12484 1756 12540
rect 1756 12484 1812 12540
rect 1812 12484 1816 12540
rect 1752 12480 1816 12484
rect 1832 12540 1896 12544
rect 1832 12484 1836 12540
rect 1836 12484 1892 12540
rect 1892 12484 1896 12540
rect 1832 12480 1896 12484
rect 1912 12540 1976 12544
rect 1912 12484 1916 12540
rect 1916 12484 1972 12540
rect 1972 12484 1976 12540
rect 1912 12480 1976 12484
rect 1992 12540 2056 12544
rect 1992 12484 1996 12540
rect 1996 12484 2052 12540
rect 2052 12484 2056 12540
rect 1992 12480 2056 12484
rect 2072 12540 2136 12544
rect 2072 12484 2076 12540
rect 2076 12484 2132 12540
rect 2132 12484 2136 12540
rect 2072 12480 2136 12484
rect 2152 12540 2216 12544
rect 2152 12484 2156 12540
rect 2156 12484 2212 12540
rect 2212 12484 2216 12540
rect 2152 12480 2216 12484
rect 2232 12540 2296 12544
rect 2232 12484 2236 12540
rect 2236 12484 2292 12540
rect 2292 12484 2296 12540
rect 2232 12480 2296 12484
rect 2312 12540 2376 12544
rect 2312 12484 2316 12540
rect 2316 12484 2372 12540
rect 2372 12484 2376 12540
rect 2312 12480 2376 12484
rect 2392 12540 2456 12544
rect 2392 12484 2396 12540
rect 2396 12484 2452 12540
rect 2452 12484 2456 12540
rect 2392 12480 2456 12484
rect 2472 12540 2536 12544
rect 2472 12484 2476 12540
rect 2476 12484 2532 12540
rect 2532 12484 2536 12540
rect 2472 12480 2536 12484
rect 2552 12540 2616 12544
rect 2552 12484 2556 12540
rect 2556 12484 2612 12540
rect 2612 12484 2616 12540
rect 2552 12480 2616 12484
rect 2632 12540 2696 12544
rect 2632 12484 2636 12540
rect 2636 12484 2692 12540
rect 2692 12484 2696 12540
rect 2632 12480 2696 12484
rect 5512 13084 5576 13088
rect 5512 13028 5516 13084
rect 5516 13028 5572 13084
rect 5572 13028 5576 13084
rect 5512 13024 5576 13028
rect 5592 13084 5656 13088
rect 5592 13028 5596 13084
rect 5596 13028 5652 13084
rect 5652 13028 5656 13084
rect 5592 13024 5656 13028
rect 5672 13084 5736 13088
rect 5672 13028 5676 13084
rect 5676 13028 5732 13084
rect 5732 13028 5736 13084
rect 5672 13024 5736 13028
rect 5752 13084 5816 13088
rect 5752 13028 5756 13084
rect 5756 13028 5812 13084
rect 5812 13028 5816 13084
rect 5752 13024 5816 13028
rect 5832 13084 5896 13088
rect 5832 13028 5836 13084
rect 5836 13028 5892 13084
rect 5892 13028 5896 13084
rect 5832 13024 5896 13028
rect 5912 13084 5976 13088
rect 5912 13028 5916 13084
rect 5916 13028 5972 13084
rect 5972 13028 5976 13084
rect 5912 13024 5976 13028
rect 5992 13084 6056 13088
rect 5992 13028 5996 13084
rect 5996 13028 6052 13084
rect 6052 13028 6056 13084
rect 5992 13024 6056 13028
rect 6072 13084 6136 13088
rect 6072 13028 6076 13084
rect 6076 13028 6132 13084
rect 6132 13028 6136 13084
rect 6072 13024 6136 13028
rect 6152 13084 6216 13088
rect 6152 13028 6156 13084
rect 6156 13028 6212 13084
rect 6212 13028 6216 13084
rect 6152 13024 6216 13028
rect 6232 13084 6296 13088
rect 6232 13028 6236 13084
rect 6236 13028 6292 13084
rect 6292 13028 6296 13084
rect 6232 13024 6296 13028
rect 6312 13084 6376 13088
rect 6312 13028 6316 13084
rect 6316 13028 6372 13084
rect 6372 13028 6376 13084
rect 6312 13024 6376 13028
rect 6392 13084 6456 13088
rect 6392 13028 6396 13084
rect 6396 13028 6452 13084
rect 6452 13028 6456 13084
rect 6392 13024 6456 13028
rect 6472 13084 6536 13088
rect 6472 13028 6476 13084
rect 6476 13028 6532 13084
rect 6532 13028 6536 13084
rect 6472 13024 6536 13028
rect 6552 13084 6616 13088
rect 6552 13028 6556 13084
rect 6556 13028 6612 13084
rect 6612 13028 6616 13084
rect 6552 13024 6616 13028
rect 6632 13084 6696 13088
rect 6632 13028 6636 13084
rect 6636 13028 6692 13084
rect 6692 13028 6696 13084
rect 6632 13024 6696 13028
rect 9512 13628 9576 13632
rect 9512 13572 9516 13628
rect 9516 13572 9572 13628
rect 9572 13572 9576 13628
rect 9512 13568 9576 13572
rect 9592 13628 9656 13632
rect 9592 13572 9596 13628
rect 9596 13572 9652 13628
rect 9652 13572 9656 13628
rect 9592 13568 9656 13572
rect 9672 13628 9736 13632
rect 9672 13572 9676 13628
rect 9676 13572 9732 13628
rect 9732 13572 9736 13628
rect 9672 13568 9736 13572
rect 9752 13628 9816 13632
rect 9752 13572 9756 13628
rect 9756 13572 9812 13628
rect 9812 13572 9816 13628
rect 9752 13568 9816 13572
rect 9832 13628 9896 13632
rect 9832 13572 9836 13628
rect 9836 13572 9892 13628
rect 9892 13572 9896 13628
rect 9832 13568 9896 13572
rect 9912 13628 9976 13632
rect 9912 13572 9916 13628
rect 9916 13572 9972 13628
rect 9972 13572 9976 13628
rect 9912 13568 9976 13572
rect 9992 13628 10056 13632
rect 9992 13572 9996 13628
rect 9996 13572 10052 13628
rect 10052 13572 10056 13628
rect 9992 13568 10056 13572
rect 10072 13628 10136 13632
rect 10072 13572 10076 13628
rect 10076 13572 10132 13628
rect 10132 13572 10136 13628
rect 10072 13568 10136 13572
rect 10152 13628 10216 13632
rect 10152 13572 10156 13628
rect 10156 13572 10212 13628
rect 10212 13572 10216 13628
rect 10152 13568 10216 13572
rect 10232 13628 10296 13632
rect 10232 13572 10236 13628
rect 10236 13572 10292 13628
rect 10292 13572 10296 13628
rect 10232 13568 10296 13572
rect 10312 13628 10376 13632
rect 10312 13572 10316 13628
rect 10316 13572 10372 13628
rect 10372 13572 10376 13628
rect 10312 13568 10376 13572
rect 10392 13628 10456 13632
rect 10392 13572 10396 13628
rect 10396 13572 10452 13628
rect 10452 13572 10456 13628
rect 10392 13568 10456 13572
rect 10472 13628 10536 13632
rect 10472 13572 10476 13628
rect 10476 13572 10532 13628
rect 10532 13572 10536 13628
rect 10472 13568 10536 13572
rect 10552 13628 10616 13632
rect 10552 13572 10556 13628
rect 10556 13572 10612 13628
rect 10612 13572 10616 13628
rect 10552 13568 10616 13572
rect 10632 13628 10696 13632
rect 10632 13572 10636 13628
rect 10636 13572 10692 13628
rect 10692 13572 10696 13628
rect 10632 13568 10696 13572
rect 17512 13628 17576 13632
rect 17512 13572 17516 13628
rect 17516 13572 17572 13628
rect 17572 13572 17576 13628
rect 17512 13568 17576 13572
rect 17592 13628 17656 13632
rect 17592 13572 17596 13628
rect 17596 13572 17652 13628
rect 17652 13572 17656 13628
rect 17592 13568 17656 13572
rect 17672 13628 17736 13632
rect 17672 13572 17676 13628
rect 17676 13572 17732 13628
rect 17732 13572 17736 13628
rect 17672 13568 17736 13572
rect 17752 13628 17816 13632
rect 17752 13572 17756 13628
rect 17756 13572 17812 13628
rect 17812 13572 17816 13628
rect 17752 13568 17816 13572
rect 17832 13628 17896 13632
rect 17832 13572 17836 13628
rect 17836 13572 17892 13628
rect 17892 13572 17896 13628
rect 17832 13568 17896 13572
rect 17912 13628 17976 13632
rect 17912 13572 17916 13628
rect 17916 13572 17972 13628
rect 17972 13572 17976 13628
rect 17912 13568 17976 13572
rect 17992 13628 18056 13632
rect 17992 13572 17996 13628
rect 17996 13572 18052 13628
rect 18052 13572 18056 13628
rect 17992 13568 18056 13572
rect 18072 13628 18136 13632
rect 18072 13572 18076 13628
rect 18076 13572 18132 13628
rect 18132 13572 18136 13628
rect 18072 13568 18136 13572
rect 18152 13628 18216 13632
rect 18152 13572 18156 13628
rect 18156 13572 18212 13628
rect 18212 13572 18216 13628
rect 18152 13568 18216 13572
rect 18232 13628 18296 13632
rect 18232 13572 18236 13628
rect 18236 13572 18292 13628
rect 18292 13572 18296 13628
rect 18232 13568 18296 13572
rect 18312 13628 18376 13632
rect 18312 13572 18316 13628
rect 18316 13572 18372 13628
rect 18372 13572 18376 13628
rect 18312 13568 18376 13572
rect 18392 13628 18456 13632
rect 18392 13572 18396 13628
rect 18396 13572 18452 13628
rect 18452 13572 18456 13628
rect 18392 13568 18456 13572
rect 18472 13628 18536 13632
rect 18472 13572 18476 13628
rect 18476 13572 18532 13628
rect 18532 13572 18536 13628
rect 18472 13568 18536 13572
rect 18552 13628 18616 13632
rect 18552 13572 18556 13628
rect 18556 13572 18612 13628
rect 18612 13572 18616 13628
rect 18552 13568 18616 13572
rect 18632 13628 18696 13632
rect 18632 13572 18636 13628
rect 18636 13572 18692 13628
rect 18692 13572 18696 13628
rect 18632 13568 18696 13572
rect 5512 11996 5576 12000
rect 5512 11940 5516 11996
rect 5516 11940 5572 11996
rect 5572 11940 5576 11996
rect 5512 11936 5576 11940
rect 5592 11996 5656 12000
rect 5592 11940 5596 11996
rect 5596 11940 5652 11996
rect 5652 11940 5656 11996
rect 5592 11936 5656 11940
rect 5672 11996 5736 12000
rect 5672 11940 5676 11996
rect 5676 11940 5732 11996
rect 5732 11940 5736 11996
rect 5672 11936 5736 11940
rect 5752 11996 5816 12000
rect 5752 11940 5756 11996
rect 5756 11940 5812 11996
rect 5812 11940 5816 11996
rect 5752 11936 5816 11940
rect 5832 11996 5896 12000
rect 5832 11940 5836 11996
rect 5836 11940 5892 11996
rect 5892 11940 5896 11996
rect 5832 11936 5896 11940
rect 5912 11996 5976 12000
rect 5912 11940 5916 11996
rect 5916 11940 5972 11996
rect 5972 11940 5976 11996
rect 5912 11936 5976 11940
rect 5992 11996 6056 12000
rect 5992 11940 5996 11996
rect 5996 11940 6052 11996
rect 6052 11940 6056 11996
rect 5992 11936 6056 11940
rect 6072 11996 6136 12000
rect 6072 11940 6076 11996
rect 6076 11940 6132 11996
rect 6132 11940 6136 11996
rect 6072 11936 6136 11940
rect 6152 11996 6216 12000
rect 6152 11940 6156 11996
rect 6156 11940 6212 11996
rect 6212 11940 6216 11996
rect 6152 11936 6216 11940
rect 6232 11996 6296 12000
rect 6232 11940 6236 11996
rect 6236 11940 6292 11996
rect 6292 11940 6296 11996
rect 6232 11936 6296 11940
rect 6312 11996 6376 12000
rect 6312 11940 6316 11996
rect 6316 11940 6372 11996
rect 6372 11940 6376 11996
rect 6312 11936 6376 11940
rect 6392 11996 6456 12000
rect 6392 11940 6396 11996
rect 6396 11940 6452 11996
rect 6452 11940 6456 11996
rect 6392 11936 6456 11940
rect 6472 11996 6536 12000
rect 6472 11940 6476 11996
rect 6476 11940 6532 11996
rect 6532 11940 6536 11996
rect 6472 11936 6536 11940
rect 6552 11996 6616 12000
rect 6552 11940 6556 11996
rect 6556 11940 6612 11996
rect 6612 11940 6616 11996
rect 6552 11936 6616 11940
rect 6632 11996 6696 12000
rect 6632 11940 6636 11996
rect 6636 11940 6692 11996
rect 6692 11940 6696 11996
rect 6632 11936 6696 11940
rect 9512 12540 9576 12544
rect 9512 12484 9516 12540
rect 9516 12484 9572 12540
rect 9572 12484 9576 12540
rect 9512 12480 9576 12484
rect 9592 12540 9656 12544
rect 9592 12484 9596 12540
rect 9596 12484 9652 12540
rect 9652 12484 9656 12540
rect 9592 12480 9656 12484
rect 9672 12540 9736 12544
rect 9672 12484 9676 12540
rect 9676 12484 9732 12540
rect 9732 12484 9736 12540
rect 9672 12480 9736 12484
rect 9752 12540 9816 12544
rect 9752 12484 9756 12540
rect 9756 12484 9812 12540
rect 9812 12484 9816 12540
rect 9752 12480 9816 12484
rect 9832 12540 9896 12544
rect 9832 12484 9836 12540
rect 9836 12484 9892 12540
rect 9892 12484 9896 12540
rect 9832 12480 9896 12484
rect 9912 12540 9976 12544
rect 9912 12484 9916 12540
rect 9916 12484 9972 12540
rect 9972 12484 9976 12540
rect 9912 12480 9976 12484
rect 9992 12540 10056 12544
rect 9992 12484 9996 12540
rect 9996 12484 10052 12540
rect 10052 12484 10056 12540
rect 9992 12480 10056 12484
rect 10072 12540 10136 12544
rect 10072 12484 10076 12540
rect 10076 12484 10132 12540
rect 10132 12484 10136 12540
rect 10072 12480 10136 12484
rect 10152 12540 10216 12544
rect 10152 12484 10156 12540
rect 10156 12484 10212 12540
rect 10212 12484 10216 12540
rect 10152 12480 10216 12484
rect 10232 12540 10296 12544
rect 10232 12484 10236 12540
rect 10236 12484 10292 12540
rect 10292 12484 10296 12540
rect 10232 12480 10296 12484
rect 10312 12540 10376 12544
rect 10312 12484 10316 12540
rect 10316 12484 10372 12540
rect 10372 12484 10376 12540
rect 10312 12480 10376 12484
rect 10392 12540 10456 12544
rect 10392 12484 10396 12540
rect 10396 12484 10452 12540
rect 10452 12484 10456 12540
rect 10392 12480 10456 12484
rect 10472 12540 10536 12544
rect 10472 12484 10476 12540
rect 10476 12484 10532 12540
rect 10532 12484 10536 12540
rect 10472 12480 10536 12484
rect 10552 12540 10616 12544
rect 10552 12484 10556 12540
rect 10556 12484 10612 12540
rect 10612 12484 10616 12540
rect 10552 12480 10616 12484
rect 10632 12540 10696 12544
rect 10632 12484 10636 12540
rect 10636 12484 10692 12540
rect 10692 12484 10696 12540
rect 10632 12480 10696 12484
rect 1512 11452 1576 11456
rect 1512 11396 1516 11452
rect 1516 11396 1572 11452
rect 1572 11396 1576 11452
rect 1512 11392 1576 11396
rect 1592 11452 1656 11456
rect 1592 11396 1596 11452
rect 1596 11396 1652 11452
rect 1652 11396 1656 11452
rect 1592 11392 1656 11396
rect 1672 11452 1736 11456
rect 1672 11396 1676 11452
rect 1676 11396 1732 11452
rect 1732 11396 1736 11452
rect 1672 11392 1736 11396
rect 1752 11452 1816 11456
rect 1752 11396 1756 11452
rect 1756 11396 1812 11452
rect 1812 11396 1816 11452
rect 1752 11392 1816 11396
rect 1832 11452 1896 11456
rect 1832 11396 1836 11452
rect 1836 11396 1892 11452
rect 1892 11396 1896 11452
rect 1832 11392 1896 11396
rect 1912 11452 1976 11456
rect 1912 11396 1916 11452
rect 1916 11396 1972 11452
rect 1972 11396 1976 11452
rect 1912 11392 1976 11396
rect 1992 11452 2056 11456
rect 1992 11396 1996 11452
rect 1996 11396 2052 11452
rect 2052 11396 2056 11452
rect 1992 11392 2056 11396
rect 2072 11452 2136 11456
rect 2072 11396 2076 11452
rect 2076 11396 2132 11452
rect 2132 11396 2136 11452
rect 2072 11392 2136 11396
rect 2152 11452 2216 11456
rect 2152 11396 2156 11452
rect 2156 11396 2212 11452
rect 2212 11396 2216 11452
rect 2152 11392 2216 11396
rect 2232 11452 2296 11456
rect 2232 11396 2236 11452
rect 2236 11396 2292 11452
rect 2292 11396 2296 11452
rect 2232 11392 2296 11396
rect 2312 11452 2376 11456
rect 2312 11396 2316 11452
rect 2316 11396 2372 11452
rect 2372 11396 2376 11452
rect 2312 11392 2376 11396
rect 2392 11452 2456 11456
rect 2392 11396 2396 11452
rect 2396 11396 2452 11452
rect 2452 11396 2456 11452
rect 2392 11392 2456 11396
rect 2472 11452 2536 11456
rect 2472 11396 2476 11452
rect 2476 11396 2532 11452
rect 2532 11396 2536 11452
rect 2472 11392 2536 11396
rect 2552 11452 2616 11456
rect 2552 11396 2556 11452
rect 2556 11396 2612 11452
rect 2612 11396 2616 11452
rect 2552 11392 2616 11396
rect 2632 11452 2696 11456
rect 2632 11396 2636 11452
rect 2636 11396 2692 11452
rect 2692 11396 2696 11452
rect 2632 11392 2696 11396
rect 5512 10908 5576 10912
rect 5512 10852 5516 10908
rect 5516 10852 5572 10908
rect 5572 10852 5576 10908
rect 5512 10848 5576 10852
rect 5592 10908 5656 10912
rect 5592 10852 5596 10908
rect 5596 10852 5652 10908
rect 5652 10852 5656 10908
rect 5592 10848 5656 10852
rect 5672 10908 5736 10912
rect 5672 10852 5676 10908
rect 5676 10852 5732 10908
rect 5732 10852 5736 10908
rect 5672 10848 5736 10852
rect 5752 10908 5816 10912
rect 5752 10852 5756 10908
rect 5756 10852 5812 10908
rect 5812 10852 5816 10908
rect 5752 10848 5816 10852
rect 5832 10908 5896 10912
rect 5832 10852 5836 10908
rect 5836 10852 5892 10908
rect 5892 10852 5896 10908
rect 5832 10848 5896 10852
rect 5912 10908 5976 10912
rect 5912 10852 5916 10908
rect 5916 10852 5972 10908
rect 5972 10852 5976 10908
rect 5912 10848 5976 10852
rect 5992 10908 6056 10912
rect 5992 10852 5996 10908
rect 5996 10852 6052 10908
rect 6052 10852 6056 10908
rect 5992 10848 6056 10852
rect 6072 10908 6136 10912
rect 6072 10852 6076 10908
rect 6076 10852 6132 10908
rect 6132 10852 6136 10908
rect 6072 10848 6136 10852
rect 6152 10908 6216 10912
rect 6152 10852 6156 10908
rect 6156 10852 6212 10908
rect 6212 10852 6216 10908
rect 6152 10848 6216 10852
rect 6232 10908 6296 10912
rect 6232 10852 6236 10908
rect 6236 10852 6292 10908
rect 6292 10852 6296 10908
rect 6232 10848 6296 10852
rect 6312 10908 6376 10912
rect 6312 10852 6316 10908
rect 6316 10852 6372 10908
rect 6372 10852 6376 10908
rect 6312 10848 6376 10852
rect 6392 10908 6456 10912
rect 6392 10852 6396 10908
rect 6396 10852 6452 10908
rect 6452 10852 6456 10908
rect 6392 10848 6456 10852
rect 6472 10908 6536 10912
rect 6472 10852 6476 10908
rect 6476 10852 6532 10908
rect 6532 10852 6536 10908
rect 6472 10848 6536 10852
rect 6552 10908 6616 10912
rect 6552 10852 6556 10908
rect 6556 10852 6612 10908
rect 6612 10852 6616 10908
rect 6552 10848 6616 10852
rect 6632 10908 6696 10912
rect 6632 10852 6636 10908
rect 6636 10852 6692 10908
rect 6692 10852 6696 10908
rect 6632 10848 6696 10852
rect 9512 11452 9576 11456
rect 9512 11396 9516 11452
rect 9516 11396 9572 11452
rect 9572 11396 9576 11452
rect 9512 11392 9576 11396
rect 9592 11452 9656 11456
rect 9592 11396 9596 11452
rect 9596 11396 9652 11452
rect 9652 11396 9656 11452
rect 9592 11392 9656 11396
rect 9672 11452 9736 11456
rect 9672 11396 9676 11452
rect 9676 11396 9732 11452
rect 9732 11396 9736 11452
rect 9672 11392 9736 11396
rect 9752 11452 9816 11456
rect 9752 11396 9756 11452
rect 9756 11396 9812 11452
rect 9812 11396 9816 11452
rect 9752 11392 9816 11396
rect 9832 11452 9896 11456
rect 9832 11396 9836 11452
rect 9836 11396 9892 11452
rect 9892 11396 9896 11452
rect 9832 11392 9896 11396
rect 9912 11452 9976 11456
rect 9912 11396 9916 11452
rect 9916 11396 9972 11452
rect 9972 11396 9976 11452
rect 9912 11392 9976 11396
rect 9992 11452 10056 11456
rect 9992 11396 9996 11452
rect 9996 11396 10052 11452
rect 10052 11396 10056 11452
rect 9992 11392 10056 11396
rect 10072 11452 10136 11456
rect 10072 11396 10076 11452
rect 10076 11396 10132 11452
rect 10132 11396 10136 11452
rect 10072 11392 10136 11396
rect 10152 11452 10216 11456
rect 10152 11396 10156 11452
rect 10156 11396 10212 11452
rect 10212 11396 10216 11452
rect 10152 11392 10216 11396
rect 10232 11452 10296 11456
rect 10232 11396 10236 11452
rect 10236 11396 10292 11452
rect 10292 11396 10296 11452
rect 10232 11392 10296 11396
rect 10312 11452 10376 11456
rect 10312 11396 10316 11452
rect 10316 11396 10372 11452
rect 10372 11396 10376 11452
rect 10312 11392 10376 11396
rect 10392 11452 10456 11456
rect 10392 11396 10396 11452
rect 10396 11396 10452 11452
rect 10452 11396 10456 11452
rect 10392 11392 10456 11396
rect 10472 11452 10536 11456
rect 10472 11396 10476 11452
rect 10476 11396 10532 11452
rect 10532 11396 10536 11452
rect 10472 11392 10536 11396
rect 10552 11452 10616 11456
rect 10552 11396 10556 11452
rect 10556 11396 10612 11452
rect 10612 11396 10616 11452
rect 10552 11392 10616 11396
rect 10632 11452 10696 11456
rect 10632 11396 10636 11452
rect 10636 11396 10692 11452
rect 10692 11396 10696 11452
rect 10632 11392 10696 11396
rect 13512 13084 13576 13088
rect 13512 13028 13516 13084
rect 13516 13028 13572 13084
rect 13572 13028 13576 13084
rect 13512 13024 13576 13028
rect 13592 13084 13656 13088
rect 13592 13028 13596 13084
rect 13596 13028 13652 13084
rect 13652 13028 13656 13084
rect 13592 13024 13656 13028
rect 13672 13084 13736 13088
rect 13672 13028 13676 13084
rect 13676 13028 13732 13084
rect 13732 13028 13736 13084
rect 13672 13024 13736 13028
rect 13752 13084 13816 13088
rect 13752 13028 13756 13084
rect 13756 13028 13812 13084
rect 13812 13028 13816 13084
rect 13752 13024 13816 13028
rect 13832 13084 13896 13088
rect 13832 13028 13836 13084
rect 13836 13028 13892 13084
rect 13892 13028 13896 13084
rect 13832 13024 13896 13028
rect 13912 13084 13976 13088
rect 13912 13028 13916 13084
rect 13916 13028 13972 13084
rect 13972 13028 13976 13084
rect 13912 13024 13976 13028
rect 13992 13084 14056 13088
rect 13992 13028 13996 13084
rect 13996 13028 14052 13084
rect 14052 13028 14056 13084
rect 13992 13024 14056 13028
rect 14072 13084 14136 13088
rect 14072 13028 14076 13084
rect 14076 13028 14132 13084
rect 14132 13028 14136 13084
rect 14072 13024 14136 13028
rect 14152 13084 14216 13088
rect 14152 13028 14156 13084
rect 14156 13028 14212 13084
rect 14212 13028 14216 13084
rect 14152 13024 14216 13028
rect 14232 13084 14296 13088
rect 14232 13028 14236 13084
rect 14236 13028 14292 13084
rect 14292 13028 14296 13084
rect 14232 13024 14296 13028
rect 14312 13084 14376 13088
rect 14312 13028 14316 13084
rect 14316 13028 14372 13084
rect 14372 13028 14376 13084
rect 14312 13024 14376 13028
rect 14392 13084 14456 13088
rect 14392 13028 14396 13084
rect 14396 13028 14452 13084
rect 14452 13028 14456 13084
rect 14392 13024 14456 13028
rect 14472 13084 14536 13088
rect 14472 13028 14476 13084
rect 14476 13028 14532 13084
rect 14532 13028 14536 13084
rect 14472 13024 14536 13028
rect 14552 13084 14616 13088
rect 14552 13028 14556 13084
rect 14556 13028 14612 13084
rect 14612 13028 14616 13084
rect 14552 13024 14616 13028
rect 14632 13084 14696 13088
rect 14632 13028 14636 13084
rect 14636 13028 14692 13084
rect 14692 13028 14696 13084
rect 14632 13024 14696 13028
rect 17512 12540 17576 12544
rect 17512 12484 17516 12540
rect 17516 12484 17572 12540
rect 17572 12484 17576 12540
rect 17512 12480 17576 12484
rect 17592 12540 17656 12544
rect 17592 12484 17596 12540
rect 17596 12484 17652 12540
rect 17652 12484 17656 12540
rect 17592 12480 17656 12484
rect 17672 12540 17736 12544
rect 17672 12484 17676 12540
rect 17676 12484 17732 12540
rect 17732 12484 17736 12540
rect 17672 12480 17736 12484
rect 17752 12540 17816 12544
rect 17752 12484 17756 12540
rect 17756 12484 17812 12540
rect 17812 12484 17816 12540
rect 17752 12480 17816 12484
rect 17832 12540 17896 12544
rect 17832 12484 17836 12540
rect 17836 12484 17892 12540
rect 17892 12484 17896 12540
rect 17832 12480 17896 12484
rect 17912 12540 17976 12544
rect 17912 12484 17916 12540
rect 17916 12484 17972 12540
rect 17972 12484 17976 12540
rect 17912 12480 17976 12484
rect 17992 12540 18056 12544
rect 17992 12484 17996 12540
rect 17996 12484 18052 12540
rect 18052 12484 18056 12540
rect 17992 12480 18056 12484
rect 18072 12540 18136 12544
rect 18072 12484 18076 12540
rect 18076 12484 18132 12540
rect 18132 12484 18136 12540
rect 18072 12480 18136 12484
rect 18152 12540 18216 12544
rect 18152 12484 18156 12540
rect 18156 12484 18212 12540
rect 18212 12484 18216 12540
rect 18152 12480 18216 12484
rect 18232 12540 18296 12544
rect 18232 12484 18236 12540
rect 18236 12484 18292 12540
rect 18292 12484 18296 12540
rect 18232 12480 18296 12484
rect 18312 12540 18376 12544
rect 18312 12484 18316 12540
rect 18316 12484 18372 12540
rect 18372 12484 18376 12540
rect 18312 12480 18376 12484
rect 18392 12540 18456 12544
rect 18392 12484 18396 12540
rect 18396 12484 18452 12540
rect 18452 12484 18456 12540
rect 18392 12480 18456 12484
rect 18472 12540 18536 12544
rect 18472 12484 18476 12540
rect 18476 12484 18532 12540
rect 18532 12484 18536 12540
rect 18472 12480 18536 12484
rect 18552 12540 18616 12544
rect 18552 12484 18556 12540
rect 18556 12484 18612 12540
rect 18612 12484 18616 12540
rect 18552 12480 18616 12484
rect 18632 12540 18696 12544
rect 18632 12484 18636 12540
rect 18636 12484 18692 12540
rect 18692 12484 18696 12540
rect 18632 12480 18696 12484
rect 13512 11996 13576 12000
rect 13512 11940 13516 11996
rect 13516 11940 13572 11996
rect 13572 11940 13576 11996
rect 13512 11936 13576 11940
rect 13592 11996 13656 12000
rect 13592 11940 13596 11996
rect 13596 11940 13652 11996
rect 13652 11940 13656 11996
rect 13592 11936 13656 11940
rect 13672 11996 13736 12000
rect 13672 11940 13676 11996
rect 13676 11940 13732 11996
rect 13732 11940 13736 11996
rect 13672 11936 13736 11940
rect 13752 11996 13816 12000
rect 13752 11940 13756 11996
rect 13756 11940 13812 11996
rect 13812 11940 13816 11996
rect 13752 11936 13816 11940
rect 13832 11996 13896 12000
rect 13832 11940 13836 11996
rect 13836 11940 13892 11996
rect 13892 11940 13896 11996
rect 13832 11936 13896 11940
rect 13912 11996 13976 12000
rect 13912 11940 13916 11996
rect 13916 11940 13972 11996
rect 13972 11940 13976 11996
rect 13912 11936 13976 11940
rect 13992 11996 14056 12000
rect 13992 11940 13996 11996
rect 13996 11940 14052 11996
rect 14052 11940 14056 11996
rect 13992 11936 14056 11940
rect 14072 11996 14136 12000
rect 14072 11940 14076 11996
rect 14076 11940 14132 11996
rect 14132 11940 14136 11996
rect 14072 11936 14136 11940
rect 14152 11996 14216 12000
rect 14152 11940 14156 11996
rect 14156 11940 14212 11996
rect 14212 11940 14216 11996
rect 14152 11936 14216 11940
rect 14232 11996 14296 12000
rect 14232 11940 14236 11996
rect 14236 11940 14292 11996
rect 14292 11940 14296 11996
rect 14232 11936 14296 11940
rect 14312 11996 14376 12000
rect 14312 11940 14316 11996
rect 14316 11940 14372 11996
rect 14372 11940 14376 11996
rect 14312 11936 14376 11940
rect 14392 11996 14456 12000
rect 14392 11940 14396 11996
rect 14396 11940 14452 11996
rect 14452 11940 14456 11996
rect 14392 11936 14456 11940
rect 14472 11996 14536 12000
rect 14472 11940 14476 11996
rect 14476 11940 14532 11996
rect 14532 11940 14536 11996
rect 14472 11936 14536 11940
rect 14552 11996 14616 12000
rect 14552 11940 14556 11996
rect 14556 11940 14612 11996
rect 14612 11940 14616 11996
rect 14552 11936 14616 11940
rect 14632 11996 14696 12000
rect 14632 11940 14636 11996
rect 14636 11940 14692 11996
rect 14692 11940 14696 11996
rect 14632 11936 14696 11940
rect 18828 11596 18892 11660
rect 17512 11452 17576 11456
rect 17512 11396 17516 11452
rect 17516 11396 17572 11452
rect 17572 11396 17576 11452
rect 17512 11392 17576 11396
rect 17592 11452 17656 11456
rect 17592 11396 17596 11452
rect 17596 11396 17652 11452
rect 17652 11396 17656 11452
rect 17592 11392 17656 11396
rect 17672 11452 17736 11456
rect 17672 11396 17676 11452
rect 17676 11396 17732 11452
rect 17732 11396 17736 11452
rect 17672 11392 17736 11396
rect 17752 11452 17816 11456
rect 17752 11396 17756 11452
rect 17756 11396 17812 11452
rect 17812 11396 17816 11452
rect 17752 11392 17816 11396
rect 17832 11452 17896 11456
rect 17832 11396 17836 11452
rect 17836 11396 17892 11452
rect 17892 11396 17896 11452
rect 17832 11392 17896 11396
rect 17912 11452 17976 11456
rect 17912 11396 17916 11452
rect 17916 11396 17972 11452
rect 17972 11396 17976 11452
rect 17912 11392 17976 11396
rect 17992 11452 18056 11456
rect 17992 11396 17996 11452
rect 17996 11396 18052 11452
rect 18052 11396 18056 11452
rect 17992 11392 18056 11396
rect 18072 11452 18136 11456
rect 18072 11396 18076 11452
rect 18076 11396 18132 11452
rect 18132 11396 18136 11452
rect 18072 11392 18136 11396
rect 18152 11452 18216 11456
rect 18152 11396 18156 11452
rect 18156 11396 18212 11452
rect 18212 11396 18216 11452
rect 18152 11392 18216 11396
rect 18232 11452 18296 11456
rect 18232 11396 18236 11452
rect 18236 11396 18292 11452
rect 18292 11396 18296 11452
rect 18232 11392 18296 11396
rect 18312 11452 18376 11456
rect 18312 11396 18316 11452
rect 18316 11396 18372 11452
rect 18372 11396 18376 11452
rect 18312 11392 18376 11396
rect 18392 11452 18456 11456
rect 18392 11396 18396 11452
rect 18396 11396 18452 11452
rect 18452 11396 18456 11452
rect 18392 11392 18456 11396
rect 18472 11452 18536 11456
rect 18472 11396 18476 11452
rect 18476 11396 18532 11452
rect 18532 11396 18536 11452
rect 18472 11392 18536 11396
rect 18552 11452 18616 11456
rect 18552 11396 18556 11452
rect 18556 11396 18612 11452
rect 18612 11396 18616 11452
rect 18552 11392 18616 11396
rect 18632 11452 18696 11456
rect 18632 11396 18636 11452
rect 18636 11396 18692 11452
rect 18692 11396 18696 11452
rect 18632 11392 18696 11396
rect 13512 10908 13576 10912
rect 13512 10852 13516 10908
rect 13516 10852 13572 10908
rect 13572 10852 13576 10908
rect 13512 10848 13576 10852
rect 13592 10908 13656 10912
rect 13592 10852 13596 10908
rect 13596 10852 13652 10908
rect 13652 10852 13656 10908
rect 13592 10848 13656 10852
rect 13672 10908 13736 10912
rect 13672 10852 13676 10908
rect 13676 10852 13732 10908
rect 13732 10852 13736 10908
rect 13672 10848 13736 10852
rect 13752 10908 13816 10912
rect 13752 10852 13756 10908
rect 13756 10852 13812 10908
rect 13812 10852 13816 10908
rect 13752 10848 13816 10852
rect 13832 10908 13896 10912
rect 13832 10852 13836 10908
rect 13836 10852 13892 10908
rect 13892 10852 13896 10908
rect 13832 10848 13896 10852
rect 13912 10908 13976 10912
rect 13912 10852 13916 10908
rect 13916 10852 13972 10908
rect 13972 10852 13976 10908
rect 13912 10848 13976 10852
rect 13992 10908 14056 10912
rect 13992 10852 13996 10908
rect 13996 10852 14052 10908
rect 14052 10852 14056 10908
rect 13992 10848 14056 10852
rect 14072 10908 14136 10912
rect 14072 10852 14076 10908
rect 14076 10852 14132 10908
rect 14132 10852 14136 10908
rect 14072 10848 14136 10852
rect 14152 10908 14216 10912
rect 14152 10852 14156 10908
rect 14156 10852 14212 10908
rect 14212 10852 14216 10908
rect 14152 10848 14216 10852
rect 14232 10908 14296 10912
rect 14232 10852 14236 10908
rect 14236 10852 14292 10908
rect 14292 10852 14296 10908
rect 14232 10848 14296 10852
rect 14312 10908 14376 10912
rect 14312 10852 14316 10908
rect 14316 10852 14372 10908
rect 14372 10852 14376 10908
rect 14312 10848 14376 10852
rect 14392 10908 14456 10912
rect 14392 10852 14396 10908
rect 14396 10852 14452 10908
rect 14452 10852 14456 10908
rect 14392 10848 14456 10852
rect 14472 10908 14536 10912
rect 14472 10852 14476 10908
rect 14476 10852 14532 10908
rect 14532 10852 14536 10908
rect 14472 10848 14536 10852
rect 14552 10908 14616 10912
rect 14552 10852 14556 10908
rect 14556 10852 14612 10908
rect 14612 10852 14616 10908
rect 14552 10848 14616 10852
rect 14632 10908 14696 10912
rect 14632 10852 14636 10908
rect 14636 10852 14692 10908
rect 14692 10852 14696 10908
rect 14632 10848 14696 10852
rect 1512 10364 1576 10368
rect 1512 10308 1516 10364
rect 1516 10308 1572 10364
rect 1572 10308 1576 10364
rect 1512 10304 1576 10308
rect 1592 10364 1656 10368
rect 1592 10308 1596 10364
rect 1596 10308 1652 10364
rect 1652 10308 1656 10364
rect 1592 10304 1656 10308
rect 1672 10364 1736 10368
rect 1672 10308 1676 10364
rect 1676 10308 1732 10364
rect 1732 10308 1736 10364
rect 1672 10304 1736 10308
rect 1752 10364 1816 10368
rect 1752 10308 1756 10364
rect 1756 10308 1812 10364
rect 1812 10308 1816 10364
rect 1752 10304 1816 10308
rect 1832 10364 1896 10368
rect 1832 10308 1836 10364
rect 1836 10308 1892 10364
rect 1892 10308 1896 10364
rect 1832 10304 1896 10308
rect 1912 10364 1976 10368
rect 1912 10308 1916 10364
rect 1916 10308 1972 10364
rect 1972 10308 1976 10364
rect 1912 10304 1976 10308
rect 1992 10364 2056 10368
rect 1992 10308 1996 10364
rect 1996 10308 2052 10364
rect 2052 10308 2056 10364
rect 1992 10304 2056 10308
rect 2072 10364 2136 10368
rect 2072 10308 2076 10364
rect 2076 10308 2132 10364
rect 2132 10308 2136 10364
rect 2072 10304 2136 10308
rect 2152 10364 2216 10368
rect 2152 10308 2156 10364
rect 2156 10308 2212 10364
rect 2212 10308 2216 10364
rect 2152 10304 2216 10308
rect 2232 10364 2296 10368
rect 2232 10308 2236 10364
rect 2236 10308 2292 10364
rect 2292 10308 2296 10364
rect 2232 10304 2296 10308
rect 2312 10364 2376 10368
rect 2312 10308 2316 10364
rect 2316 10308 2372 10364
rect 2372 10308 2376 10364
rect 2312 10304 2376 10308
rect 2392 10364 2456 10368
rect 2392 10308 2396 10364
rect 2396 10308 2452 10364
rect 2452 10308 2456 10364
rect 2392 10304 2456 10308
rect 2472 10364 2536 10368
rect 2472 10308 2476 10364
rect 2476 10308 2532 10364
rect 2532 10308 2536 10364
rect 2472 10304 2536 10308
rect 2552 10364 2616 10368
rect 2552 10308 2556 10364
rect 2556 10308 2612 10364
rect 2612 10308 2616 10364
rect 2552 10304 2616 10308
rect 2632 10364 2696 10368
rect 2632 10308 2636 10364
rect 2636 10308 2692 10364
rect 2692 10308 2696 10364
rect 2632 10304 2696 10308
rect 9512 10364 9576 10368
rect 9512 10308 9516 10364
rect 9516 10308 9572 10364
rect 9572 10308 9576 10364
rect 9512 10304 9576 10308
rect 9592 10364 9656 10368
rect 9592 10308 9596 10364
rect 9596 10308 9652 10364
rect 9652 10308 9656 10364
rect 9592 10304 9656 10308
rect 9672 10364 9736 10368
rect 9672 10308 9676 10364
rect 9676 10308 9732 10364
rect 9732 10308 9736 10364
rect 9672 10304 9736 10308
rect 9752 10364 9816 10368
rect 9752 10308 9756 10364
rect 9756 10308 9812 10364
rect 9812 10308 9816 10364
rect 9752 10304 9816 10308
rect 9832 10364 9896 10368
rect 9832 10308 9836 10364
rect 9836 10308 9892 10364
rect 9892 10308 9896 10364
rect 9832 10304 9896 10308
rect 9912 10364 9976 10368
rect 9912 10308 9916 10364
rect 9916 10308 9972 10364
rect 9972 10308 9976 10364
rect 9912 10304 9976 10308
rect 9992 10364 10056 10368
rect 9992 10308 9996 10364
rect 9996 10308 10052 10364
rect 10052 10308 10056 10364
rect 9992 10304 10056 10308
rect 10072 10364 10136 10368
rect 10072 10308 10076 10364
rect 10076 10308 10132 10364
rect 10132 10308 10136 10364
rect 10072 10304 10136 10308
rect 10152 10364 10216 10368
rect 10152 10308 10156 10364
rect 10156 10308 10212 10364
rect 10212 10308 10216 10364
rect 10152 10304 10216 10308
rect 10232 10364 10296 10368
rect 10232 10308 10236 10364
rect 10236 10308 10292 10364
rect 10292 10308 10296 10364
rect 10232 10304 10296 10308
rect 10312 10364 10376 10368
rect 10312 10308 10316 10364
rect 10316 10308 10372 10364
rect 10372 10308 10376 10364
rect 10312 10304 10376 10308
rect 10392 10364 10456 10368
rect 10392 10308 10396 10364
rect 10396 10308 10452 10364
rect 10452 10308 10456 10364
rect 10392 10304 10456 10308
rect 10472 10364 10536 10368
rect 10472 10308 10476 10364
rect 10476 10308 10532 10364
rect 10532 10308 10536 10364
rect 10472 10304 10536 10308
rect 10552 10364 10616 10368
rect 10552 10308 10556 10364
rect 10556 10308 10612 10364
rect 10612 10308 10616 10364
rect 10552 10304 10616 10308
rect 10632 10364 10696 10368
rect 10632 10308 10636 10364
rect 10636 10308 10692 10364
rect 10692 10308 10696 10364
rect 10632 10304 10696 10308
rect 19012 10644 19076 10708
rect 17512 10364 17576 10368
rect 17512 10308 17516 10364
rect 17516 10308 17572 10364
rect 17572 10308 17576 10364
rect 17512 10304 17576 10308
rect 17592 10364 17656 10368
rect 17592 10308 17596 10364
rect 17596 10308 17652 10364
rect 17652 10308 17656 10364
rect 17592 10304 17656 10308
rect 17672 10364 17736 10368
rect 17672 10308 17676 10364
rect 17676 10308 17732 10364
rect 17732 10308 17736 10364
rect 17672 10304 17736 10308
rect 17752 10364 17816 10368
rect 17752 10308 17756 10364
rect 17756 10308 17812 10364
rect 17812 10308 17816 10364
rect 17752 10304 17816 10308
rect 17832 10364 17896 10368
rect 17832 10308 17836 10364
rect 17836 10308 17892 10364
rect 17892 10308 17896 10364
rect 17832 10304 17896 10308
rect 17912 10364 17976 10368
rect 17912 10308 17916 10364
rect 17916 10308 17972 10364
rect 17972 10308 17976 10364
rect 17912 10304 17976 10308
rect 17992 10364 18056 10368
rect 17992 10308 17996 10364
rect 17996 10308 18052 10364
rect 18052 10308 18056 10364
rect 17992 10304 18056 10308
rect 18072 10364 18136 10368
rect 18072 10308 18076 10364
rect 18076 10308 18132 10364
rect 18132 10308 18136 10364
rect 18072 10304 18136 10308
rect 18152 10364 18216 10368
rect 18152 10308 18156 10364
rect 18156 10308 18212 10364
rect 18212 10308 18216 10364
rect 18152 10304 18216 10308
rect 18232 10364 18296 10368
rect 18232 10308 18236 10364
rect 18236 10308 18292 10364
rect 18292 10308 18296 10364
rect 18232 10304 18296 10308
rect 18312 10364 18376 10368
rect 18312 10308 18316 10364
rect 18316 10308 18372 10364
rect 18372 10308 18376 10364
rect 18312 10304 18376 10308
rect 18392 10364 18456 10368
rect 18392 10308 18396 10364
rect 18396 10308 18452 10364
rect 18452 10308 18456 10364
rect 18392 10304 18456 10308
rect 18472 10364 18536 10368
rect 18472 10308 18476 10364
rect 18476 10308 18532 10364
rect 18532 10308 18536 10364
rect 18472 10304 18536 10308
rect 18552 10364 18616 10368
rect 18552 10308 18556 10364
rect 18556 10308 18612 10364
rect 18612 10308 18616 10364
rect 18552 10304 18616 10308
rect 18632 10364 18696 10368
rect 18632 10308 18636 10364
rect 18636 10308 18692 10364
rect 18692 10308 18696 10364
rect 18632 10304 18696 10308
rect 5512 9820 5576 9824
rect 5512 9764 5516 9820
rect 5516 9764 5572 9820
rect 5572 9764 5576 9820
rect 5512 9760 5576 9764
rect 5592 9820 5656 9824
rect 5592 9764 5596 9820
rect 5596 9764 5652 9820
rect 5652 9764 5656 9820
rect 5592 9760 5656 9764
rect 5672 9820 5736 9824
rect 5672 9764 5676 9820
rect 5676 9764 5732 9820
rect 5732 9764 5736 9820
rect 5672 9760 5736 9764
rect 5752 9820 5816 9824
rect 5752 9764 5756 9820
rect 5756 9764 5812 9820
rect 5812 9764 5816 9820
rect 5752 9760 5816 9764
rect 5832 9820 5896 9824
rect 5832 9764 5836 9820
rect 5836 9764 5892 9820
rect 5892 9764 5896 9820
rect 5832 9760 5896 9764
rect 5912 9820 5976 9824
rect 5912 9764 5916 9820
rect 5916 9764 5972 9820
rect 5972 9764 5976 9820
rect 5912 9760 5976 9764
rect 5992 9820 6056 9824
rect 5992 9764 5996 9820
rect 5996 9764 6052 9820
rect 6052 9764 6056 9820
rect 5992 9760 6056 9764
rect 6072 9820 6136 9824
rect 6072 9764 6076 9820
rect 6076 9764 6132 9820
rect 6132 9764 6136 9820
rect 6072 9760 6136 9764
rect 6152 9820 6216 9824
rect 6152 9764 6156 9820
rect 6156 9764 6212 9820
rect 6212 9764 6216 9820
rect 6152 9760 6216 9764
rect 6232 9820 6296 9824
rect 6232 9764 6236 9820
rect 6236 9764 6292 9820
rect 6292 9764 6296 9820
rect 6232 9760 6296 9764
rect 6312 9820 6376 9824
rect 6312 9764 6316 9820
rect 6316 9764 6372 9820
rect 6372 9764 6376 9820
rect 6312 9760 6376 9764
rect 6392 9820 6456 9824
rect 6392 9764 6396 9820
rect 6396 9764 6452 9820
rect 6452 9764 6456 9820
rect 6392 9760 6456 9764
rect 6472 9820 6536 9824
rect 6472 9764 6476 9820
rect 6476 9764 6532 9820
rect 6532 9764 6536 9820
rect 6472 9760 6536 9764
rect 6552 9820 6616 9824
rect 6552 9764 6556 9820
rect 6556 9764 6612 9820
rect 6612 9764 6616 9820
rect 6552 9760 6616 9764
rect 6632 9820 6696 9824
rect 6632 9764 6636 9820
rect 6636 9764 6692 9820
rect 6692 9764 6696 9820
rect 6632 9760 6696 9764
rect 13512 9820 13576 9824
rect 13512 9764 13516 9820
rect 13516 9764 13572 9820
rect 13572 9764 13576 9820
rect 13512 9760 13576 9764
rect 13592 9820 13656 9824
rect 13592 9764 13596 9820
rect 13596 9764 13652 9820
rect 13652 9764 13656 9820
rect 13592 9760 13656 9764
rect 13672 9820 13736 9824
rect 13672 9764 13676 9820
rect 13676 9764 13732 9820
rect 13732 9764 13736 9820
rect 13672 9760 13736 9764
rect 13752 9820 13816 9824
rect 13752 9764 13756 9820
rect 13756 9764 13812 9820
rect 13812 9764 13816 9820
rect 13752 9760 13816 9764
rect 13832 9820 13896 9824
rect 13832 9764 13836 9820
rect 13836 9764 13892 9820
rect 13892 9764 13896 9820
rect 13832 9760 13896 9764
rect 13912 9820 13976 9824
rect 13912 9764 13916 9820
rect 13916 9764 13972 9820
rect 13972 9764 13976 9820
rect 13912 9760 13976 9764
rect 13992 9820 14056 9824
rect 13992 9764 13996 9820
rect 13996 9764 14052 9820
rect 14052 9764 14056 9820
rect 13992 9760 14056 9764
rect 14072 9820 14136 9824
rect 14072 9764 14076 9820
rect 14076 9764 14132 9820
rect 14132 9764 14136 9820
rect 14072 9760 14136 9764
rect 14152 9820 14216 9824
rect 14152 9764 14156 9820
rect 14156 9764 14212 9820
rect 14212 9764 14216 9820
rect 14152 9760 14216 9764
rect 14232 9820 14296 9824
rect 14232 9764 14236 9820
rect 14236 9764 14292 9820
rect 14292 9764 14296 9820
rect 14232 9760 14296 9764
rect 14312 9820 14376 9824
rect 14312 9764 14316 9820
rect 14316 9764 14372 9820
rect 14372 9764 14376 9820
rect 14312 9760 14376 9764
rect 14392 9820 14456 9824
rect 14392 9764 14396 9820
rect 14396 9764 14452 9820
rect 14452 9764 14456 9820
rect 14392 9760 14456 9764
rect 14472 9820 14536 9824
rect 14472 9764 14476 9820
rect 14476 9764 14532 9820
rect 14532 9764 14536 9820
rect 14472 9760 14536 9764
rect 14552 9820 14616 9824
rect 14552 9764 14556 9820
rect 14556 9764 14612 9820
rect 14612 9764 14616 9820
rect 14552 9760 14616 9764
rect 14632 9820 14696 9824
rect 14632 9764 14636 9820
rect 14636 9764 14692 9820
rect 14692 9764 14696 9820
rect 14632 9760 14696 9764
rect 1512 9276 1576 9280
rect 1512 9220 1516 9276
rect 1516 9220 1572 9276
rect 1572 9220 1576 9276
rect 1512 9216 1576 9220
rect 1592 9276 1656 9280
rect 1592 9220 1596 9276
rect 1596 9220 1652 9276
rect 1652 9220 1656 9276
rect 1592 9216 1656 9220
rect 1672 9276 1736 9280
rect 1672 9220 1676 9276
rect 1676 9220 1732 9276
rect 1732 9220 1736 9276
rect 1672 9216 1736 9220
rect 1752 9276 1816 9280
rect 1752 9220 1756 9276
rect 1756 9220 1812 9276
rect 1812 9220 1816 9276
rect 1752 9216 1816 9220
rect 1832 9276 1896 9280
rect 1832 9220 1836 9276
rect 1836 9220 1892 9276
rect 1892 9220 1896 9276
rect 1832 9216 1896 9220
rect 1912 9276 1976 9280
rect 1912 9220 1916 9276
rect 1916 9220 1972 9276
rect 1972 9220 1976 9276
rect 1912 9216 1976 9220
rect 1992 9276 2056 9280
rect 1992 9220 1996 9276
rect 1996 9220 2052 9276
rect 2052 9220 2056 9276
rect 1992 9216 2056 9220
rect 2072 9276 2136 9280
rect 2072 9220 2076 9276
rect 2076 9220 2132 9276
rect 2132 9220 2136 9276
rect 2072 9216 2136 9220
rect 2152 9276 2216 9280
rect 2152 9220 2156 9276
rect 2156 9220 2212 9276
rect 2212 9220 2216 9276
rect 2152 9216 2216 9220
rect 2232 9276 2296 9280
rect 2232 9220 2236 9276
rect 2236 9220 2292 9276
rect 2292 9220 2296 9276
rect 2232 9216 2296 9220
rect 2312 9276 2376 9280
rect 2312 9220 2316 9276
rect 2316 9220 2372 9276
rect 2372 9220 2376 9276
rect 2312 9216 2376 9220
rect 2392 9276 2456 9280
rect 2392 9220 2396 9276
rect 2396 9220 2452 9276
rect 2452 9220 2456 9276
rect 2392 9216 2456 9220
rect 2472 9276 2536 9280
rect 2472 9220 2476 9276
rect 2476 9220 2532 9276
rect 2532 9220 2536 9276
rect 2472 9216 2536 9220
rect 2552 9276 2616 9280
rect 2552 9220 2556 9276
rect 2556 9220 2612 9276
rect 2612 9220 2616 9276
rect 2552 9216 2616 9220
rect 2632 9276 2696 9280
rect 2632 9220 2636 9276
rect 2636 9220 2692 9276
rect 2692 9220 2696 9276
rect 2632 9216 2696 9220
rect 9512 9276 9576 9280
rect 9512 9220 9516 9276
rect 9516 9220 9572 9276
rect 9572 9220 9576 9276
rect 9512 9216 9576 9220
rect 9592 9276 9656 9280
rect 9592 9220 9596 9276
rect 9596 9220 9652 9276
rect 9652 9220 9656 9276
rect 9592 9216 9656 9220
rect 9672 9276 9736 9280
rect 9672 9220 9676 9276
rect 9676 9220 9732 9276
rect 9732 9220 9736 9276
rect 9672 9216 9736 9220
rect 9752 9276 9816 9280
rect 9752 9220 9756 9276
rect 9756 9220 9812 9276
rect 9812 9220 9816 9276
rect 9752 9216 9816 9220
rect 9832 9276 9896 9280
rect 9832 9220 9836 9276
rect 9836 9220 9892 9276
rect 9892 9220 9896 9276
rect 9832 9216 9896 9220
rect 9912 9276 9976 9280
rect 9912 9220 9916 9276
rect 9916 9220 9972 9276
rect 9972 9220 9976 9276
rect 9912 9216 9976 9220
rect 9992 9276 10056 9280
rect 9992 9220 9996 9276
rect 9996 9220 10052 9276
rect 10052 9220 10056 9276
rect 9992 9216 10056 9220
rect 10072 9276 10136 9280
rect 10072 9220 10076 9276
rect 10076 9220 10132 9276
rect 10132 9220 10136 9276
rect 10072 9216 10136 9220
rect 10152 9276 10216 9280
rect 10152 9220 10156 9276
rect 10156 9220 10212 9276
rect 10212 9220 10216 9276
rect 10152 9216 10216 9220
rect 10232 9276 10296 9280
rect 10232 9220 10236 9276
rect 10236 9220 10292 9276
rect 10292 9220 10296 9276
rect 10232 9216 10296 9220
rect 10312 9276 10376 9280
rect 10312 9220 10316 9276
rect 10316 9220 10372 9276
rect 10372 9220 10376 9276
rect 10312 9216 10376 9220
rect 10392 9276 10456 9280
rect 10392 9220 10396 9276
rect 10396 9220 10452 9276
rect 10452 9220 10456 9276
rect 10392 9216 10456 9220
rect 10472 9276 10536 9280
rect 10472 9220 10476 9276
rect 10476 9220 10532 9276
rect 10532 9220 10536 9276
rect 10472 9216 10536 9220
rect 10552 9276 10616 9280
rect 10552 9220 10556 9276
rect 10556 9220 10612 9276
rect 10612 9220 10616 9276
rect 10552 9216 10616 9220
rect 10632 9276 10696 9280
rect 10632 9220 10636 9276
rect 10636 9220 10692 9276
rect 10692 9220 10696 9276
rect 10632 9216 10696 9220
rect 19196 9420 19260 9484
rect 17512 9276 17576 9280
rect 17512 9220 17516 9276
rect 17516 9220 17572 9276
rect 17572 9220 17576 9276
rect 17512 9216 17576 9220
rect 17592 9276 17656 9280
rect 17592 9220 17596 9276
rect 17596 9220 17652 9276
rect 17652 9220 17656 9276
rect 17592 9216 17656 9220
rect 17672 9276 17736 9280
rect 17672 9220 17676 9276
rect 17676 9220 17732 9276
rect 17732 9220 17736 9276
rect 17672 9216 17736 9220
rect 17752 9276 17816 9280
rect 17752 9220 17756 9276
rect 17756 9220 17812 9276
rect 17812 9220 17816 9276
rect 17752 9216 17816 9220
rect 17832 9276 17896 9280
rect 17832 9220 17836 9276
rect 17836 9220 17892 9276
rect 17892 9220 17896 9276
rect 17832 9216 17896 9220
rect 17912 9276 17976 9280
rect 17912 9220 17916 9276
rect 17916 9220 17972 9276
rect 17972 9220 17976 9276
rect 17912 9216 17976 9220
rect 17992 9276 18056 9280
rect 17992 9220 17996 9276
rect 17996 9220 18052 9276
rect 18052 9220 18056 9276
rect 17992 9216 18056 9220
rect 18072 9276 18136 9280
rect 18072 9220 18076 9276
rect 18076 9220 18132 9276
rect 18132 9220 18136 9276
rect 18072 9216 18136 9220
rect 18152 9276 18216 9280
rect 18152 9220 18156 9276
rect 18156 9220 18212 9276
rect 18212 9220 18216 9276
rect 18152 9216 18216 9220
rect 18232 9276 18296 9280
rect 18232 9220 18236 9276
rect 18236 9220 18292 9276
rect 18292 9220 18296 9276
rect 18232 9216 18296 9220
rect 18312 9276 18376 9280
rect 18312 9220 18316 9276
rect 18316 9220 18372 9276
rect 18372 9220 18376 9276
rect 18312 9216 18376 9220
rect 18392 9276 18456 9280
rect 18392 9220 18396 9276
rect 18396 9220 18452 9276
rect 18452 9220 18456 9276
rect 18392 9216 18456 9220
rect 18472 9276 18536 9280
rect 18472 9220 18476 9276
rect 18476 9220 18532 9276
rect 18532 9220 18536 9276
rect 18472 9216 18536 9220
rect 18552 9276 18616 9280
rect 18552 9220 18556 9276
rect 18556 9220 18612 9276
rect 18612 9220 18616 9276
rect 18552 9216 18616 9220
rect 18632 9276 18696 9280
rect 18632 9220 18636 9276
rect 18636 9220 18692 9276
rect 18692 9220 18696 9276
rect 18632 9216 18696 9220
rect 5512 8732 5576 8736
rect 5512 8676 5516 8732
rect 5516 8676 5572 8732
rect 5572 8676 5576 8732
rect 5512 8672 5576 8676
rect 5592 8732 5656 8736
rect 5592 8676 5596 8732
rect 5596 8676 5652 8732
rect 5652 8676 5656 8732
rect 5592 8672 5656 8676
rect 5672 8732 5736 8736
rect 5672 8676 5676 8732
rect 5676 8676 5732 8732
rect 5732 8676 5736 8732
rect 5672 8672 5736 8676
rect 5752 8732 5816 8736
rect 5752 8676 5756 8732
rect 5756 8676 5812 8732
rect 5812 8676 5816 8732
rect 5752 8672 5816 8676
rect 5832 8732 5896 8736
rect 5832 8676 5836 8732
rect 5836 8676 5892 8732
rect 5892 8676 5896 8732
rect 5832 8672 5896 8676
rect 5912 8732 5976 8736
rect 5912 8676 5916 8732
rect 5916 8676 5972 8732
rect 5972 8676 5976 8732
rect 5912 8672 5976 8676
rect 5992 8732 6056 8736
rect 5992 8676 5996 8732
rect 5996 8676 6052 8732
rect 6052 8676 6056 8732
rect 5992 8672 6056 8676
rect 6072 8732 6136 8736
rect 6072 8676 6076 8732
rect 6076 8676 6132 8732
rect 6132 8676 6136 8732
rect 6072 8672 6136 8676
rect 6152 8732 6216 8736
rect 6152 8676 6156 8732
rect 6156 8676 6212 8732
rect 6212 8676 6216 8732
rect 6152 8672 6216 8676
rect 6232 8732 6296 8736
rect 6232 8676 6236 8732
rect 6236 8676 6292 8732
rect 6292 8676 6296 8732
rect 6232 8672 6296 8676
rect 6312 8732 6376 8736
rect 6312 8676 6316 8732
rect 6316 8676 6372 8732
rect 6372 8676 6376 8732
rect 6312 8672 6376 8676
rect 6392 8732 6456 8736
rect 6392 8676 6396 8732
rect 6396 8676 6452 8732
rect 6452 8676 6456 8732
rect 6392 8672 6456 8676
rect 6472 8732 6536 8736
rect 6472 8676 6476 8732
rect 6476 8676 6532 8732
rect 6532 8676 6536 8732
rect 6472 8672 6536 8676
rect 6552 8732 6616 8736
rect 6552 8676 6556 8732
rect 6556 8676 6612 8732
rect 6612 8676 6616 8732
rect 6552 8672 6616 8676
rect 6632 8732 6696 8736
rect 6632 8676 6636 8732
rect 6636 8676 6692 8732
rect 6692 8676 6696 8732
rect 6632 8672 6696 8676
rect 13512 8732 13576 8736
rect 13512 8676 13516 8732
rect 13516 8676 13572 8732
rect 13572 8676 13576 8732
rect 13512 8672 13576 8676
rect 13592 8732 13656 8736
rect 13592 8676 13596 8732
rect 13596 8676 13652 8732
rect 13652 8676 13656 8732
rect 13592 8672 13656 8676
rect 13672 8732 13736 8736
rect 13672 8676 13676 8732
rect 13676 8676 13732 8732
rect 13732 8676 13736 8732
rect 13672 8672 13736 8676
rect 13752 8732 13816 8736
rect 13752 8676 13756 8732
rect 13756 8676 13812 8732
rect 13812 8676 13816 8732
rect 13752 8672 13816 8676
rect 13832 8732 13896 8736
rect 13832 8676 13836 8732
rect 13836 8676 13892 8732
rect 13892 8676 13896 8732
rect 13832 8672 13896 8676
rect 13912 8732 13976 8736
rect 13912 8676 13916 8732
rect 13916 8676 13972 8732
rect 13972 8676 13976 8732
rect 13912 8672 13976 8676
rect 13992 8732 14056 8736
rect 13992 8676 13996 8732
rect 13996 8676 14052 8732
rect 14052 8676 14056 8732
rect 13992 8672 14056 8676
rect 14072 8732 14136 8736
rect 14072 8676 14076 8732
rect 14076 8676 14132 8732
rect 14132 8676 14136 8732
rect 14072 8672 14136 8676
rect 14152 8732 14216 8736
rect 14152 8676 14156 8732
rect 14156 8676 14212 8732
rect 14212 8676 14216 8732
rect 14152 8672 14216 8676
rect 14232 8732 14296 8736
rect 14232 8676 14236 8732
rect 14236 8676 14292 8732
rect 14292 8676 14296 8732
rect 14232 8672 14296 8676
rect 14312 8732 14376 8736
rect 14312 8676 14316 8732
rect 14316 8676 14372 8732
rect 14372 8676 14376 8732
rect 14312 8672 14376 8676
rect 14392 8732 14456 8736
rect 14392 8676 14396 8732
rect 14396 8676 14452 8732
rect 14452 8676 14456 8732
rect 14392 8672 14456 8676
rect 14472 8732 14536 8736
rect 14472 8676 14476 8732
rect 14476 8676 14532 8732
rect 14532 8676 14536 8732
rect 14472 8672 14536 8676
rect 14552 8732 14616 8736
rect 14552 8676 14556 8732
rect 14556 8676 14612 8732
rect 14612 8676 14616 8732
rect 14552 8672 14616 8676
rect 14632 8732 14696 8736
rect 14632 8676 14636 8732
rect 14636 8676 14692 8732
rect 14692 8676 14696 8732
rect 14632 8672 14696 8676
rect 1512 8188 1576 8192
rect 1512 8132 1516 8188
rect 1516 8132 1572 8188
rect 1572 8132 1576 8188
rect 1512 8128 1576 8132
rect 1592 8188 1656 8192
rect 1592 8132 1596 8188
rect 1596 8132 1652 8188
rect 1652 8132 1656 8188
rect 1592 8128 1656 8132
rect 1672 8188 1736 8192
rect 1672 8132 1676 8188
rect 1676 8132 1732 8188
rect 1732 8132 1736 8188
rect 1672 8128 1736 8132
rect 1752 8188 1816 8192
rect 1752 8132 1756 8188
rect 1756 8132 1812 8188
rect 1812 8132 1816 8188
rect 1752 8128 1816 8132
rect 1832 8188 1896 8192
rect 1832 8132 1836 8188
rect 1836 8132 1892 8188
rect 1892 8132 1896 8188
rect 1832 8128 1896 8132
rect 1912 8188 1976 8192
rect 1912 8132 1916 8188
rect 1916 8132 1972 8188
rect 1972 8132 1976 8188
rect 1912 8128 1976 8132
rect 1992 8188 2056 8192
rect 1992 8132 1996 8188
rect 1996 8132 2052 8188
rect 2052 8132 2056 8188
rect 1992 8128 2056 8132
rect 2072 8188 2136 8192
rect 2072 8132 2076 8188
rect 2076 8132 2132 8188
rect 2132 8132 2136 8188
rect 2072 8128 2136 8132
rect 2152 8188 2216 8192
rect 2152 8132 2156 8188
rect 2156 8132 2212 8188
rect 2212 8132 2216 8188
rect 2152 8128 2216 8132
rect 2232 8188 2296 8192
rect 2232 8132 2236 8188
rect 2236 8132 2292 8188
rect 2292 8132 2296 8188
rect 2232 8128 2296 8132
rect 2312 8188 2376 8192
rect 2312 8132 2316 8188
rect 2316 8132 2372 8188
rect 2372 8132 2376 8188
rect 2312 8128 2376 8132
rect 2392 8188 2456 8192
rect 2392 8132 2396 8188
rect 2396 8132 2452 8188
rect 2452 8132 2456 8188
rect 2392 8128 2456 8132
rect 2472 8188 2536 8192
rect 2472 8132 2476 8188
rect 2476 8132 2532 8188
rect 2532 8132 2536 8188
rect 2472 8128 2536 8132
rect 2552 8188 2616 8192
rect 2552 8132 2556 8188
rect 2556 8132 2612 8188
rect 2612 8132 2616 8188
rect 2552 8128 2616 8132
rect 2632 8188 2696 8192
rect 2632 8132 2636 8188
rect 2636 8132 2692 8188
rect 2692 8132 2696 8188
rect 2632 8128 2696 8132
rect 9512 8188 9576 8192
rect 9512 8132 9516 8188
rect 9516 8132 9572 8188
rect 9572 8132 9576 8188
rect 9512 8128 9576 8132
rect 9592 8188 9656 8192
rect 9592 8132 9596 8188
rect 9596 8132 9652 8188
rect 9652 8132 9656 8188
rect 9592 8128 9656 8132
rect 9672 8188 9736 8192
rect 9672 8132 9676 8188
rect 9676 8132 9732 8188
rect 9732 8132 9736 8188
rect 9672 8128 9736 8132
rect 9752 8188 9816 8192
rect 9752 8132 9756 8188
rect 9756 8132 9812 8188
rect 9812 8132 9816 8188
rect 9752 8128 9816 8132
rect 9832 8188 9896 8192
rect 9832 8132 9836 8188
rect 9836 8132 9892 8188
rect 9892 8132 9896 8188
rect 9832 8128 9896 8132
rect 9912 8188 9976 8192
rect 9912 8132 9916 8188
rect 9916 8132 9972 8188
rect 9972 8132 9976 8188
rect 9912 8128 9976 8132
rect 9992 8188 10056 8192
rect 9992 8132 9996 8188
rect 9996 8132 10052 8188
rect 10052 8132 10056 8188
rect 9992 8128 10056 8132
rect 10072 8188 10136 8192
rect 10072 8132 10076 8188
rect 10076 8132 10132 8188
rect 10132 8132 10136 8188
rect 10072 8128 10136 8132
rect 10152 8188 10216 8192
rect 10152 8132 10156 8188
rect 10156 8132 10212 8188
rect 10212 8132 10216 8188
rect 10152 8128 10216 8132
rect 10232 8188 10296 8192
rect 10232 8132 10236 8188
rect 10236 8132 10292 8188
rect 10292 8132 10296 8188
rect 10232 8128 10296 8132
rect 10312 8188 10376 8192
rect 10312 8132 10316 8188
rect 10316 8132 10372 8188
rect 10372 8132 10376 8188
rect 10312 8128 10376 8132
rect 10392 8188 10456 8192
rect 10392 8132 10396 8188
rect 10396 8132 10452 8188
rect 10452 8132 10456 8188
rect 10392 8128 10456 8132
rect 10472 8188 10536 8192
rect 10472 8132 10476 8188
rect 10476 8132 10532 8188
rect 10532 8132 10536 8188
rect 10472 8128 10536 8132
rect 10552 8188 10616 8192
rect 10552 8132 10556 8188
rect 10556 8132 10612 8188
rect 10612 8132 10616 8188
rect 10552 8128 10616 8132
rect 10632 8188 10696 8192
rect 10632 8132 10636 8188
rect 10636 8132 10692 8188
rect 10692 8132 10696 8188
rect 10632 8128 10696 8132
rect 17512 8188 17576 8192
rect 17512 8132 17516 8188
rect 17516 8132 17572 8188
rect 17572 8132 17576 8188
rect 17512 8128 17576 8132
rect 17592 8188 17656 8192
rect 17592 8132 17596 8188
rect 17596 8132 17652 8188
rect 17652 8132 17656 8188
rect 17592 8128 17656 8132
rect 17672 8188 17736 8192
rect 17672 8132 17676 8188
rect 17676 8132 17732 8188
rect 17732 8132 17736 8188
rect 17672 8128 17736 8132
rect 17752 8188 17816 8192
rect 17752 8132 17756 8188
rect 17756 8132 17812 8188
rect 17812 8132 17816 8188
rect 17752 8128 17816 8132
rect 17832 8188 17896 8192
rect 17832 8132 17836 8188
rect 17836 8132 17892 8188
rect 17892 8132 17896 8188
rect 17832 8128 17896 8132
rect 17912 8188 17976 8192
rect 17912 8132 17916 8188
rect 17916 8132 17972 8188
rect 17972 8132 17976 8188
rect 17912 8128 17976 8132
rect 17992 8188 18056 8192
rect 17992 8132 17996 8188
rect 17996 8132 18052 8188
rect 18052 8132 18056 8188
rect 17992 8128 18056 8132
rect 18072 8188 18136 8192
rect 18072 8132 18076 8188
rect 18076 8132 18132 8188
rect 18132 8132 18136 8188
rect 18072 8128 18136 8132
rect 18152 8188 18216 8192
rect 18152 8132 18156 8188
rect 18156 8132 18212 8188
rect 18212 8132 18216 8188
rect 18152 8128 18216 8132
rect 18232 8188 18296 8192
rect 18232 8132 18236 8188
rect 18236 8132 18292 8188
rect 18292 8132 18296 8188
rect 18232 8128 18296 8132
rect 18312 8188 18376 8192
rect 18312 8132 18316 8188
rect 18316 8132 18372 8188
rect 18372 8132 18376 8188
rect 18312 8128 18376 8132
rect 18392 8188 18456 8192
rect 18392 8132 18396 8188
rect 18396 8132 18452 8188
rect 18452 8132 18456 8188
rect 18392 8128 18456 8132
rect 18472 8188 18536 8192
rect 18472 8132 18476 8188
rect 18476 8132 18532 8188
rect 18532 8132 18536 8188
rect 18472 8128 18536 8132
rect 18552 8188 18616 8192
rect 18552 8132 18556 8188
rect 18556 8132 18612 8188
rect 18612 8132 18616 8188
rect 18552 8128 18616 8132
rect 18632 8188 18696 8192
rect 18632 8132 18636 8188
rect 18636 8132 18692 8188
rect 18692 8132 18696 8188
rect 18632 8128 18696 8132
rect 5512 7644 5576 7648
rect 5512 7588 5516 7644
rect 5516 7588 5572 7644
rect 5572 7588 5576 7644
rect 5512 7584 5576 7588
rect 5592 7644 5656 7648
rect 5592 7588 5596 7644
rect 5596 7588 5652 7644
rect 5652 7588 5656 7644
rect 5592 7584 5656 7588
rect 5672 7644 5736 7648
rect 5672 7588 5676 7644
rect 5676 7588 5732 7644
rect 5732 7588 5736 7644
rect 5672 7584 5736 7588
rect 5752 7644 5816 7648
rect 5752 7588 5756 7644
rect 5756 7588 5812 7644
rect 5812 7588 5816 7644
rect 5752 7584 5816 7588
rect 5832 7644 5896 7648
rect 5832 7588 5836 7644
rect 5836 7588 5892 7644
rect 5892 7588 5896 7644
rect 5832 7584 5896 7588
rect 5912 7644 5976 7648
rect 5912 7588 5916 7644
rect 5916 7588 5972 7644
rect 5972 7588 5976 7644
rect 5912 7584 5976 7588
rect 5992 7644 6056 7648
rect 5992 7588 5996 7644
rect 5996 7588 6052 7644
rect 6052 7588 6056 7644
rect 5992 7584 6056 7588
rect 6072 7644 6136 7648
rect 6072 7588 6076 7644
rect 6076 7588 6132 7644
rect 6132 7588 6136 7644
rect 6072 7584 6136 7588
rect 6152 7644 6216 7648
rect 6152 7588 6156 7644
rect 6156 7588 6212 7644
rect 6212 7588 6216 7644
rect 6152 7584 6216 7588
rect 6232 7644 6296 7648
rect 6232 7588 6236 7644
rect 6236 7588 6292 7644
rect 6292 7588 6296 7644
rect 6232 7584 6296 7588
rect 6312 7644 6376 7648
rect 6312 7588 6316 7644
rect 6316 7588 6372 7644
rect 6372 7588 6376 7644
rect 6312 7584 6376 7588
rect 6392 7644 6456 7648
rect 6392 7588 6396 7644
rect 6396 7588 6452 7644
rect 6452 7588 6456 7644
rect 6392 7584 6456 7588
rect 6472 7644 6536 7648
rect 6472 7588 6476 7644
rect 6476 7588 6532 7644
rect 6532 7588 6536 7644
rect 6472 7584 6536 7588
rect 6552 7644 6616 7648
rect 6552 7588 6556 7644
rect 6556 7588 6612 7644
rect 6612 7588 6616 7644
rect 6552 7584 6616 7588
rect 6632 7644 6696 7648
rect 6632 7588 6636 7644
rect 6636 7588 6692 7644
rect 6692 7588 6696 7644
rect 6632 7584 6696 7588
rect 13512 7644 13576 7648
rect 13512 7588 13516 7644
rect 13516 7588 13572 7644
rect 13572 7588 13576 7644
rect 13512 7584 13576 7588
rect 13592 7644 13656 7648
rect 13592 7588 13596 7644
rect 13596 7588 13652 7644
rect 13652 7588 13656 7644
rect 13592 7584 13656 7588
rect 13672 7644 13736 7648
rect 13672 7588 13676 7644
rect 13676 7588 13732 7644
rect 13732 7588 13736 7644
rect 13672 7584 13736 7588
rect 13752 7644 13816 7648
rect 13752 7588 13756 7644
rect 13756 7588 13812 7644
rect 13812 7588 13816 7644
rect 13752 7584 13816 7588
rect 13832 7644 13896 7648
rect 13832 7588 13836 7644
rect 13836 7588 13892 7644
rect 13892 7588 13896 7644
rect 13832 7584 13896 7588
rect 13912 7644 13976 7648
rect 13912 7588 13916 7644
rect 13916 7588 13972 7644
rect 13972 7588 13976 7644
rect 13912 7584 13976 7588
rect 13992 7644 14056 7648
rect 13992 7588 13996 7644
rect 13996 7588 14052 7644
rect 14052 7588 14056 7644
rect 13992 7584 14056 7588
rect 14072 7644 14136 7648
rect 14072 7588 14076 7644
rect 14076 7588 14132 7644
rect 14132 7588 14136 7644
rect 14072 7584 14136 7588
rect 14152 7644 14216 7648
rect 14152 7588 14156 7644
rect 14156 7588 14212 7644
rect 14212 7588 14216 7644
rect 14152 7584 14216 7588
rect 14232 7644 14296 7648
rect 14232 7588 14236 7644
rect 14236 7588 14292 7644
rect 14292 7588 14296 7644
rect 14232 7584 14296 7588
rect 14312 7644 14376 7648
rect 14312 7588 14316 7644
rect 14316 7588 14372 7644
rect 14372 7588 14376 7644
rect 14312 7584 14376 7588
rect 14392 7644 14456 7648
rect 14392 7588 14396 7644
rect 14396 7588 14452 7644
rect 14452 7588 14456 7644
rect 14392 7584 14456 7588
rect 14472 7644 14536 7648
rect 14472 7588 14476 7644
rect 14476 7588 14532 7644
rect 14532 7588 14536 7644
rect 14472 7584 14536 7588
rect 14552 7644 14616 7648
rect 14552 7588 14556 7644
rect 14556 7588 14612 7644
rect 14612 7588 14616 7644
rect 14552 7584 14616 7588
rect 14632 7644 14696 7648
rect 14632 7588 14636 7644
rect 14636 7588 14692 7644
rect 14692 7588 14696 7644
rect 14632 7584 14696 7588
rect 1512 7100 1576 7104
rect 1512 7044 1516 7100
rect 1516 7044 1572 7100
rect 1572 7044 1576 7100
rect 1512 7040 1576 7044
rect 1592 7100 1656 7104
rect 1592 7044 1596 7100
rect 1596 7044 1652 7100
rect 1652 7044 1656 7100
rect 1592 7040 1656 7044
rect 1672 7100 1736 7104
rect 1672 7044 1676 7100
rect 1676 7044 1732 7100
rect 1732 7044 1736 7100
rect 1672 7040 1736 7044
rect 1752 7100 1816 7104
rect 1752 7044 1756 7100
rect 1756 7044 1812 7100
rect 1812 7044 1816 7100
rect 1752 7040 1816 7044
rect 1832 7100 1896 7104
rect 1832 7044 1836 7100
rect 1836 7044 1892 7100
rect 1892 7044 1896 7100
rect 1832 7040 1896 7044
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 2312 7100 2376 7104
rect 2312 7044 2316 7100
rect 2316 7044 2372 7100
rect 2372 7044 2376 7100
rect 2312 7040 2376 7044
rect 2392 7100 2456 7104
rect 2392 7044 2396 7100
rect 2396 7044 2452 7100
rect 2452 7044 2456 7100
rect 2392 7040 2456 7044
rect 2472 7100 2536 7104
rect 2472 7044 2476 7100
rect 2476 7044 2532 7100
rect 2532 7044 2536 7100
rect 2472 7040 2536 7044
rect 2552 7100 2616 7104
rect 2552 7044 2556 7100
rect 2556 7044 2612 7100
rect 2612 7044 2616 7100
rect 2552 7040 2616 7044
rect 2632 7100 2696 7104
rect 2632 7044 2636 7100
rect 2636 7044 2692 7100
rect 2692 7044 2696 7100
rect 2632 7040 2696 7044
rect 9512 7100 9576 7104
rect 9512 7044 9516 7100
rect 9516 7044 9572 7100
rect 9572 7044 9576 7100
rect 9512 7040 9576 7044
rect 9592 7100 9656 7104
rect 9592 7044 9596 7100
rect 9596 7044 9652 7100
rect 9652 7044 9656 7100
rect 9592 7040 9656 7044
rect 9672 7100 9736 7104
rect 9672 7044 9676 7100
rect 9676 7044 9732 7100
rect 9732 7044 9736 7100
rect 9672 7040 9736 7044
rect 9752 7100 9816 7104
rect 9752 7044 9756 7100
rect 9756 7044 9812 7100
rect 9812 7044 9816 7100
rect 9752 7040 9816 7044
rect 9832 7100 9896 7104
rect 9832 7044 9836 7100
rect 9836 7044 9892 7100
rect 9892 7044 9896 7100
rect 9832 7040 9896 7044
rect 9912 7100 9976 7104
rect 9912 7044 9916 7100
rect 9916 7044 9972 7100
rect 9972 7044 9976 7100
rect 9912 7040 9976 7044
rect 9992 7100 10056 7104
rect 9992 7044 9996 7100
rect 9996 7044 10052 7100
rect 10052 7044 10056 7100
rect 9992 7040 10056 7044
rect 10072 7100 10136 7104
rect 10072 7044 10076 7100
rect 10076 7044 10132 7100
rect 10132 7044 10136 7100
rect 10072 7040 10136 7044
rect 10152 7100 10216 7104
rect 10152 7044 10156 7100
rect 10156 7044 10212 7100
rect 10212 7044 10216 7100
rect 10152 7040 10216 7044
rect 10232 7100 10296 7104
rect 10232 7044 10236 7100
rect 10236 7044 10292 7100
rect 10292 7044 10296 7100
rect 10232 7040 10296 7044
rect 10312 7100 10376 7104
rect 10312 7044 10316 7100
rect 10316 7044 10372 7100
rect 10372 7044 10376 7100
rect 10312 7040 10376 7044
rect 10392 7100 10456 7104
rect 10392 7044 10396 7100
rect 10396 7044 10452 7100
rect 10452 7044 10456 7100
rect 10392 7040 10456 7044
rect 10472 7100 10536 7104
rect 10472 7044 10476 7100
rect 10476 7044 10532 7100
rect 10532 7044 10536 7100
rect 10472 7040 10536 7044
rect 10552 7100 10616 7104
rect 10552 7044 10556 7100
rect 10556 7044 10612 7100
rect 10612 7044 10616 7100
rect 10552 7040 10616 7044
rect 10632 7100 10696 7104
rect 10632 7044 10636 7100
rect 10636 7044 10692 7100
rect 10692 7044 10696 7100
rect 10632 7040 10696 7044
rect 17512 7100 17576 7104
rect 17512 7044 17516 7100
rect 17516 7044 17572 7100
rect 17572 7044 17576 7100
rect 17512 7040 17576 7044
rect 17592 7100 17656 7104
rect 17592 7044 17596 7100
rect 17596 7044 17652 7100
rect 17652 7044 17656 7100
rect 17592 7040 17656 7044
rect 17672 7100 17736 7104
rect 17672 7044 17676 7100
rect 17676 7044 17732 7100
rect 17732 7044 17736 7100
rect 17672 7040 17736 7044
rect 17752 7100 17816 7104
rect 17752 7044 17756 7100
rect 17756 7044 17812 7100
rect 17812 7044 17816 7100
rect 17752 7040 17816 7044
rect 17832 7100 17896 7104
rect 17832 7044 17836 7100
rect 17836 7044 17892 7100
rect 17892 7044 17896 7100
rect 17832 7040 17896 7044
rect 17912 7100 17976 7104
rect 17912 7044 17916 7100
rect 17916 7044 17972 7100
rect 17972 7044 17976 7100
rect 17912 7040 17976 7044
rect 17992 7100 18056 7104
rect 17992 7044 17996 7100
rect 17996 7044 18052 7100
rect 18052 7044 18056 7100
rect 17992 7040 18056 7044
rect 18072 7100 18136 7104
rect 18072 7044 18076 7100
rect 18076 7044 18132 7100
rect 18132 7044 18136 7100
rect 18072 7040 18136 7044
rect 18152 7100 18216 7104
rect 18152 7044 18156 7100
rect 18156 7044 18212 7100
rect 18212 7044 18216 7100
rect 18152 7040 18216 7044
rect 18232 7100 18296 7104
rect 18232 7044 18236 7100
rect 18236 7044 18292 7100
rect 18292 7044 18296 7100
rect 18232 7040 18296 7044
rect 18312 7100 18376 7104
rect 18312 7044 18316 7100
rect 18316 7044 18372 7100
rect 18372 7044 18376 7100
rect 18312 7040 18376 7044
rect 18392 7100 18456 7104
rect 18392 7044 18396 7100
rect 18396 7044 18452 7100
rect 18452 7044 18456 7100
rect 18392 7040 18456 7044
rect 18472 7100 18536 7104
rect 18472 7044 18476 7100
rect 18476 7044 18532 7100
rect 18532 7044 18536 7100
rect 18472 7040 18536 7044
rect 18552 7100 18616 7104
rect 18552 7044 18556 7100
rect 18556 7044 18612 7100
rect 18612 7044 18616 7100
rect 18552 7040 18616 7044
rect 18632 7100 18696 7104
rect 18632 7044 18636 7100
rect 18636 7044 18692 7100
rect 18692 7044 18696 7100
rect 18632 7040 18696 7044
rect 5512 6556 5576 6560
rect 5512 6500 5516 6556
rect 5516 6500 5572 6556
rect 5572 6500 5576 6556
rect 5512 6496 5576 6500
rect 5592 6556 5656 6560
rect 5592 6500 5596 6556
rect 5596 6500 5652 6556
rect 5652 6500 5656 6556
rect 5592 6496 5656 6500
rect 5672 6556 5736 6560
rect 5672 6500 5676 6556
rect 5676 6500 5732 6556
rect 5732 6500 5736 6556
rect 5672 6496 5736 6500
rect 5752 6556 5816 6560
rect 5752 6500 5756 6556
rect 5756 6500 5812 6556
rect 5812 6500 5816 6556
rect 5752 6496 5816 6500
rect 5832 6556 5896 6560
rect 5832 6500 5836 6556
rect 5836 6500 5892 6556
rect 5892 6500 5896 6556
rect 5832 6496 5896 6500
rect 5912 6556 5976 6560
rect 5912 6500 5916 6556
rect 5916 6500 5972 6556
rect 5972 6500 5976 6556
rect 5912 6496 5976 6500
rect 5992 6556 6056 6560
rect 5992 6500 5996 6556
rect 5996 6500 6052 6556
rect 6052 6500 6056 6556
rect 5992 6496 6056 6500
rect 6072 6556 6136 6560
rect 6072 6500 6076 6556
rect 6076 6500 6132 6556
rect 6132 6500 6136 6556
rect 6072 6496 6136 6500
rect 6152 6556 6216 6560
rect 6152 6500 6156 6556
rect 6156 6500 6212 6556
rect 6212 6500 6216 6556
rect 6152 6496 6216 6500
rect 6232 6556 6296 6560
rect 6232 6500 6236 6556
rect 6236 6500 6292 6556
rect 6292 6500 6296 6556
rect 6232 6496 6296 6500
rect 6312 6556 6376 6560
rect 6312 6500 6316 6556
rect 6316 6500 6372 6556
rect 6372 6500 6376 6556
rect 6312 6496 6376 6500
rect 6392 6556 6456 6560
rect 6392 6500 6396 6556
rect 6396 6500 6452 6556
rect 6452 6500 6456 6556
rect 6392 6496 6456 6500
rect 6472 6556 6536 6560
rect 6472 6500 6476 6556
rect 6476 6500 6532 6556
rect 6532 6500 6536 6556
rect 6472 6496 6536 6500
rect 6552 6556 6616 6560
rect 6552 6500 6556 6556
rect 6556 6500 6612 6556
rect 6612 6500 6616 6556
rect 6552 6496 6616 6500
rect 6632 6556 6696 6560
rect 6632 6500 6636 6556
rect 6636 6500 6692 6556
rect 6692 6500 6696 6556
rect 6632 6496 6696 6500
rect 13512 6556 13576 6560
rect 13512 6500 13516 6556
rect 13516 6500 13572 6556
rect 13572 6500 13576 6556
rect 13512 6496 13576 6500
rect 13592 6556 13656 6560
rect 13592 6500 13596 6556
rect 13596 6500 13652 6556
rect 13652 6500 13656 6556
rect 13592 6496 13656 6500
rect 13672 6556 13736 6560
rect 13672 6500 13676 6556
rect 13676 6500 13732 6556
rect 13732 6500 13736 6556
rect 13672 6496 13736 6500
rect 13752 6556 13816 6560
rect 13752 6500 13756 6556
rect 13756 6500 13812 6556
rect 13812 6500 13816 6556
rect 13752 6496 13816 6500
rect 13832 6556 13896 6560
rect 13832 6500 13836 6556
rect 13836 6500 13892 6556
rect 13892 6500 13896 6556
rect 13832 6496 13896 6500
rect 13912 6556 13976 6560
rect 13912 6500 13916 6556
rect 13916 6500 13972 6556
rect 13972 6500 13976 6556
rect 13912 6496 13976 6500
rect 13992 6556 14056 6560
rect 13992 6500 13996 6556
rect 13996 6500 14052 6556
rect 14052 6500 14056 6556
rect 13992 6496 14056 6500
rect 14072 6556 14136 6560
rect 14072 6500 14076 6556
rect 14076 6500 14132 6556
rect 14132 6500 14136 6556
rect 14072 6496 14136 6500
rect 14152 6556 14216 6560
rect 14152 6500 14156 6556
rect 14156 6500 14212 6556
rect 14212 6500 14216 6556
rect 14152 6496 14216 6500
rect 14232 6556 14296 6560
rect 14232 6500 14236 6556
rect 14236 6500 14292 6556
rect 14292 6500 14296 6556
rect 14232 6496 14296 6500
rect 14312 6556 14376 6560
rect 14312 6500 14316 6556
rect 14316 6500 14372 6556
rect 14372 6500 14376 6556
rect 14312 6496 14376 6500
rect 14392 6556 14456 6560
rect 14392 6500 14396 6556
rect 14396 6500 14452 6556
rect 14452 6500 14456 6556
rect 14392 6496 14456 6500
rect 14472 6556 14536 6560
rect 14472 6500 14476 6556
rect 14476 6500 14532 6556
rect 14532 6500 14536 6556
rect 14472 6496 14536 6500
rect 14552 6556 14616 6560
rect 14552 6500 14556 6556
rect 14556 6500 14612 6556
rect 14612 6500 14616 6556
rect 14552 6496 14616 6500
rect 14632 6556 14696 6560
rect 14632 6500 14636 6556
rect 14636 6500 14692 6556
rect 14692 6500 14696 6556
rect 14632 6496 14696 6500
rect 1512 6012 1576 6016
rect 1512 5956 1516 6012
rect 1516 5956 1572 6012
rect 1572 5956 1576 6012
rect 1512 5952 1576 5956
rect 1592 6012 1656 6016
rect 1592 5956 1596 6012
rect 1596 5956 1652 6012
rect 1652 5956 1656 6012
rect 1592 5952 1656 5956
rect 1672 6012 1736 6016
rect 1672 5956 1676 6012
rect 1676 5956 1732 6012
rect 1732 5956 1736 6012
rect 1672 5952 1736 5956
rect 1752 6012 1816 6016
rect 1752 5956 1756 6012
rect 1756 5956 1812 6012
rect 1812 5956 1816 6012
rect 1752 5952 1816 5956
rect 1832 6012 1896 6016
rect 1832 5956 1836 6012
rect 1836 5956 1892 6012
rect 1892 5956 1896 6012
rect 1832 5952 1896 5956
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 2312 6012 2376 6016
rect 2312 5956 2316 6012
rect 2316 5956 2372 6012
rect 2372 5956 2376 6012
rect 2312 5952 2376 5956
rect 2392 6012 2456 6016
rect 2392 5956 2396 6012
rect 2396 5956 2452 6012
rect 2452 5956 2456 6012
rect 2392 5952 2456 5956
rect 2472 6012 2536 6016
rect 2472 5956 2476 6012
rect 2476 5956 2532 6012
rect 2532 5956 2536 6012
rect 2472 5952 2536 5956
rect 2552 6012 2616 6016
rect 2552 5956 2556 6012
rect 2556 5956 2612 6012
rect 2612 5956 2616 6012
rect 2552 5952 2616 5956
rect 2632 6012 2696 6016
rect 2632 5956 2636 6012
rect 2636 5956 2692 6012
rect 2692 5956 2696 6012
rect 2632 5952 2696 5956
rect 9512 6012 9576 6016
rect 9512 5956 9516 6012
rect 9516 5956 9572 6012
rect 9572 5956 9576 6012
rect 9512 5952 9576 5956
rect 9592 6012 9656 6016
rect 9592 5956 9596 6012
rect 9596 5956 9652 6012
rect 9652 5956 9656 6012
rect 9592 5952 9656 5956
rect 9672 6012 9736 6016
rect 9672 5956 9676 6012
rect 9676 5956 9732 6012
rect 9732 5956 9736 6012
rect 9672 5952 9736 5956
rect 9752 6012 9816 6016
rect 9752 5956 9756 6012
rect 9756 5956 9812 6012
rect 9812 5956 9816 6012
rect 9752 5952 9816 5956
rect 9832 6012 9896 6016
rect 9832 5956 9836 6012
rect 9836 5956 9892 6012
rect 9892 5956 9896 6012
rect 9832 5952 9896 5956
rect 9912 6012 9976 6016
rect 9912 5956 9916 6012
rect 9916 5956 9972 6012
rect 9972 5956 9976 6012
rect 9912 5952 9976 5956
rect 9992 6012 10056 6016
rect 9992 5956 9996 6012
rect 9996 5956 10052 6012
rect 10052 5956 10056 6012
rect 9992 5952 10056 5956
rect 10072 6012 10136 6016
rect 10072 5956 10076 6012
rect 10076 5956 10132 6012
rect 10132 5956 10136 6012
rect 10072 5952 10136 5956
rect 10152 6012 10216 6016
rect 10152 5956 10156 6012
rect 10156 5956 10212 6012
rect 10212 5956 10216 6012
rect 10152 5952 10216 5956
rect 10232 6012 10296 6016
rect 10232 5956 10236 6012
rect 10236 5956 10292 6012
rect 10292 5956 10296 6012
rect 10232 5952 10296 5956
rect 10312 6012 10376 6016
rect 10312 5956 10316 6012
rect 10316 5956 10372 6012
rect 10372 5956 10376 6012
rect 10312 5952 10376 5956
rect 10392 6012 10456 6016
rect 10392 5956 10396 6012
rect 10396 5956 10452 6012
rect 10452 5956 10456 6012
rect 10392 5952 10456 5956
rect 10472 6012 10536 6016
rect 10472 5956 10476 6012
rect 10476 5956 10532 6012
rect 10532 5956 10536 6012
rect 10472 5952 10536 5956
rect 10552 6012 10616 6016
rect 10552 5956 10556 6012
rect 10556 5956 10612 6012
rect 10612 5956 10616 6012
rect 10552 5952 10616 5956
rect 10632 6012 10696 6016
rect 10632 5956 10636 6012
rect 10636 5956 10692 6012
rect 10692 5956 10696 6012
rect 10632 5952 10696 5956
rect 17512 6012 17576 6016
rect 17512 5956 17516 6012
rect 17516 5956 17572 6012
rect 17572 5956 17576 6012
rect 17512 5952 17576 5956
rect 17592 6012 17656 6016
rect 17592 5956 17596 6012
rect 17596 5956 17652 6012
rect 17652 5956 17656 6012
rect 17592 5952 17656 5956
rect 17672 6012 17736 6016
rect 17672 5956 17676 6012
rect 17676 5956 17732 6012
rect 17732 5956 17736 6012
rect 17672 5952 17736 5956
rect 17752 6012 17816 6016
rect 17752 5956 17756 6012
rect 17756 5956 17812 6012
rect 17812 5956 17816 6012
rect 17752 5952 17816 5956
rect 17832 6012 17896 6016
rect 17832 5956 17836 6012
rect 17836 5956 17892 6012
rect 17892 5956 17896 6012
rect 17832 5952 17896 5956
rect 17912 6012 17976 6016
rect 17912 5956 17916 6012
rect 17916 5956 17972 6012
rect 17972 5956 17976 6012
rect 17912 5952 17976 5956
rect 17992 6012 18056 6016
rect 17992 5956 17996 6012
rect 17996 5956 18052 6012
rect 18052 5956 18056 6012
rect 17992 5952 18056 5956
rect 18072 6012 18136 6016
rect 18072 5956 18076 6012
rect 18076 5956 18132 6012
rect 18132 5956 18136 6012
rect 18072 5952 18136 5956
rect 18152 6012 18216 6016
rect 18152 5956 18156 6012
rect 18156 5956 18212 6012
rect 18212 5956 18216 6012
rect 18152 5952 18216 5956
rect 18232 6012 18296 6016
rect 18232 5956 18236 6012
rect 18236 5956 18292 6012
rect 18292 5956 18296 6012
rect 18232 5952 18296 5956
rect 18312 6012 18376 6016
rect 18312 5956 18316 6012
rect 18316 5956 18372 6012
rect 18372 5956 18376 6012
rect 18312 5952 18376 5956
rect 18392 6012 18456 6016
rect 18392 5956 18396 6012
rect 18396 5956 18452 6012
rect 18452 5956 18456 6012
rect 18392 5952 18456 5956
rect 18472 6012 18536 6016
rect 18472 5956 18476 6012
rect 18476 5956 18532 6012
rect 18532 5956 18536 6012
rect 18472 5952 18536 5956
rect 18552 6012 18616 6016
rect 18552 5956 18556 6012
rect 18556 5956 18612 6012
rect 18612 5956 18616 6012
rect 18552 5952 18616 5956
rect 18632 6012 18696 6016
rect 18632 5956 18636 6012
rect 18636 5956 18692 6012
rect 18692 5956 18696 6012
rect 18632 5952 18696 5956
rect 5512 5468 5576 5472
rect 5512 5412 5516 5468
rect 5516 5412 5572 5468
rect 5572 5412 5576 5468
rect 5512 5408 5576 5412
rect 5592 5468 5656 5472
rect 5592 5412 5596 5468
rect 5596 5412 5652 5468
rect 5652 5412 5656 5468
rect 5592 5408 5656 5412
rect 5672 5468 5736 5472
rect 5672 5412 5676 5468
rect 5676 5412 5732 5468
rect 5732 5412 5736 5468
rect 5672 5408 5736 5412
rect 5752 5468 5816 5472
rect 5752 5412 5756 5468
rect 5756 5412 5812 5468
rect 5812 5412 5816 5468
rect 5752 5408 5816 5412
rect 5832 5468 5896 5472
rect 5832 5412 5836 5468
rect 5836 5412 5892 5468
rect 5892 5412 5896 5468
rect 5832 5408 5896 5412
rect 5912 5468 5976 5472
rect 5912 5412 5916 5468
rect 5916 5412 5972 5468
rect 5972 5412 5976 5468
rect 5912 5408 5976 5412
rect 5992 5468 6056 5472
rect 5992 5412 5996 5468
rect 5996 5412 6052 5468
rect 6052 5412 6056 5468
rect 5992 5408 6056 5412
rect 6072 5468 6136 5472
rect 6072 5412 6076 5468
rect 6076 5412 6132 5468
rect 6132 5412 6136 5468
rect 6072 5408 6136 5412
rect 6152 5468 6216 5472
rect 6152 5412 6156 5468
rect 6156 5412 6212 5468
rect 6212 5412 6216 5468
rect 6152 5408 6216 5412
rect 6232 5468 6296 5472
rect 6232 5412 6236 5468
rect 6236 5412 6292 5468
rect 6292 5412 6296 5468
rect 6232 5408 6296 5412
rect 6312 5468 6376 5472
rect 6312 5412 6316 5468
rect 6316 5412 6372 5468
rect 6372 5412 6376 5468
rect 6312 5408 6376 5412
rect 6392 5468 6456 5472
rect 6392 5412 6396 5468
rect 6396 5412 6452 5468
rect 6452 5412 6456 5468
rect 6392 5408 6456 5412
rect 6472 5468 6536 5472
rect 6472 5412 6476 5468
rect 6476 5412 6532 5468
rect 6532 5412 6536 5468
rect 6472 5408 6536 5412
rect 6552 5468 6616 5472
rect 6552 5412 6556 5468
rect 6556 5412 6612 5468
rect 6612 5412 6616 5468
rect 6552 5408 6616 5412
rect 6632 5468 6696 5472
rect 6632 5412 6636 5468
rect 6636 5412 6692 5468
rect 6692 5412 6696 5468
rect 6632 5408 6696 5412
rect 13512 5468 13576 5472
rect 13512 5412 13516 5468
rect 13516 5412 13572 5468
rect 13572 5412 13576 5468
rect 13512 5408 13576 5412
rect 13592 5468 13656 5472
rect 13592 5412 13596 5468
rect 13596 5412 13652 5468
rect 13652 5412 13656 5468
rect 13592 5408 13656 5412
rect 13672 5468 13736 5472
rect 13672 5412 13676 5468
rect 13676 5412 13732 5468
rect 13732 5412 13736 5468
rect 13672 5408 13736 5412
rect 13752 5468 13816 5472
rect 13752 5412 13756 5468
rect 13756 5412 13812 5468
rect 13812 5412 13816 5468
rect 13752 5408 13816 5412
rect 13832 5468 13896 5472
rect 13832 5412 13836 5468
rect 13836 5412 13892 5468
rect 13892 5412 13896 5468
rect 13832 5408 13896 5412
rect 13912 5468 13976 5472
rect 13912 5412 13916 5468
rect 13916 5412 13972 5468
rect 13972 5412 13976 5468
rect 13912 5408 13976 5412
rect 13992 5468 14056 5472
rect 13992 5412 13996 5468
rect 13996 5412 14052 5468
rect 14052 5412 14056 5468
rect 13992 5408 14056 5412
rect 14072 5468 14136 5472
rect 14072 5412 14076 5468
rect 14076 5412 14132 5468
rect 14132 5412 14136 5468
rect 14072 5408 14136 5412
rect 14152 5468 14216 5472
rect 14152 5412 14156 5468
rect 14156 5412 14212 5468
rect 14212 5412 14216 5468
rect 14152 5408 14216 5412
rect 14232 5468 14296 5472
rect 14232 5412 14236 5468
rect 14236 5412 14292 5468
rect 14292 5412 14296 5468
rect 14232 5408 14296 5412
rect 14312 5468 14376 5472
rect 14312 5412 14316 5468
rect 14316 5412 14372 5468
rect 14372 5412 14376 5468
rect 14312 5408 14376 5412
rect 14392 5468 14456 5472
rect 14392 5412 14396 5468
rect 14396 5412 14452 5468
rect 14452 5412 14456 5468
rect 14392 5408 14456 5412
rect 14472 5468 14536 5472
rect 14472 5412 14476 5468
rect 14476 5412 14532 5468
rect 14532 5412 14536 5468
rect 14472 5408 14536 5412
rect 14552 5468 14616 5472
rect 14552 5412 14556 5468
rect 14556 5412 14612 5468
rect 14612 5412 14616 5468
rect 14552 5408 14616 5412
rect 14632 5468 14696 5472
rect 14632 5412 14636 5468
rect 14636 5412 14692 5468
rect 14692 5412 14696 5468
rect 14632 5408 14696 5412
rect 18828 5068 18892 5132
rect 1512 4924 1576 4928
rect 1512 4868 1516 4924
rect 1516 4868 1572 4924
rect 1572 4868 1576 4924
rect 1512 4864 1576 4868
rect 1592 4924 1656 4928
rect 1592 4868 1596 4924
rect 1596 4868 1652 4924
rect 1652 4868 1656 4924
rect 1592 4864 1656 4868
rect 1672 4924 1736 4928
rect 1672 4868 1676 4924
rect 1676 4868 1732 4924
rect 1732 4868 1736 4924
rect 1672 4864 1736 4868
rect 1752 4924 1816 4928
rect 1752 4868 1756 4924
rect 1756 4868 1812 4924
rect 1812 4868 1816 4924
rect 1752 4864 1816 4868
rect 1832 4924 1896 4928
rect 1832 4868 1836 4924
rect 1836 4868 1892 4924
rect 1892 4868 1896 4924
rect 1832 4864 1896 4868
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 2312 4924 2376 4928
rect 2312 4868 2316 4924
rect 2316 4868 2372 4924
rect 2372 4868 2376 4924
rect 2312 4864 2376 4868
rect 2392 4924 2456 4928
rect 2392 4868 2396 4924
rect 2396 4868 2452 4924
rect 2452 4868 2456 4924
rect 2392 4864 2456 4868
rect 2472 4924 2536 4928
rect 2472 4868 2476 4924
rect 2476 4868 2532 4924
rect 2532 4868 2536 4924
rect 2472 4864 2536 4868
rect 2552 4924 2616 4928
rect 2552 4868 2556 4924
rect 2556 4868 2612 4924
rect 2612 4868 2616 4924
rect 2552 4864 2616 4868
rect 2632 4924 2696 4928
rect 2632 4868 2636 4924
rect 2636 4868 2692 4924
rect 2692 4868 2696 4924
rect 2632 4864 2696 4868
rect 9512 4924 9576 4928
rect 9512 4868 9516 4924
rect 9516 4868 9572 4924
rect 9572 4868 9576 4924
rect 9512 4864 9576 4868
rect 9592 4924 9656 4928
rect 9592 4868 9596 4924
rect 9596 4868 9652 4924
rect 9652 4868 9656 4924
rect 9592 4864 9656 4868
rect 9672 4924 9736 4928
rect 9672 4868 9676 4924
rect 9676 4868 9732 4924
rect 9732 4868 9736 4924
rect 9672 4864 9736 4868
rect 9752 4924 9816 4928
rect 9752 4868 9756 4924
rect 9756 4868 9812 4924
rect 9812 4868 9816 4924
rect 9752 4864 9816 4868
rect 9832 4924 9896 4928
rect 9832 4868 9836 4924
rect 9836 4868 9892 4924
rect 9892 4868 9896 4924
rect 9832 4864 9896 4868
rect 9912 4924 9976 4928
rect 9912 4868 9916 4924
rect 9916 4868 9972 4924
rect 9972 4868 9976 4924
rect 9912 4864 9976 4868
rect 9992 4924 10056 4928
rect 9992 4868 9996 4924
rect 9996 4868 10052 4924
rect 10052 4868 10056 4924
rect 9992 4864 10056 4868
rect 10072 4924 10136 4928
rect 10072 4868 10076 4924
rect 10076 4868 10132 4924
rect 10132 4868 10136 4924
rect 10072 4864 10136 4868
rect 10152 4924 10216 4928
rect 10152 4868 10156 4924
rect 10156 4868 10212 4924
rect 10212 4868 10216 4924
rect 10152 4864 10216 4868
rect 10232 4924 10296 4928
rect 10232 4868 10236 4924
rect 10236 4868 10292 4924
rect 10292 4868 10296 4924
rect 10232 4864 10296 4868
rect 10312 4924 10376 4928
rect 10312 4868 10316 4924
rect 10316 4868 10372 4924
rect 10372 4868 10376 4924
rect 10312 4864 10376 4868
rect 10392 4924 10456 4928
rect 10392 4868 10396 4924
rect 10396 4868 10452 4924
rect 10452 4868 10456 4924
rect 10392 4864 10456 4868
rect 10472 4924 10536 4928
rect 10472 4868 10476 4924
rect 10476 4868 10532 4924
rect 10532 4868 10536 4924
rect 10472 4864 10536 4868
rect 10552 4924 10616 4928
rect 10552 4868 10556 4924
rect 10556 4868 10612 4924
rect 10612 4868 10616 4924
rect 10552 4864 10616 4868
rect 10632 4924 10696 4928
rect 10632 4868 10636 4924
rect 10636 4868 10692 4924
rect 10692 4868 10696 4924
rect 10632 4864 10696 4868
rect 17512 4924 17576 4928
rect 17512 4868 17516 4924
rect 17516 4868 17572 4924
rect 17572 4868 17576 4924
rect 17512 4864 17576 4868
rect 17592 4924 17656 4928
rect 17592 4868 17596 4924
rect 17596 4868 17652 4924
rect 17652 4868 17656 4924
rect 17592 4864 17656 4868
rect 17672 4924 17736 4928
rect 17672 4868 17676 4924
rect 17676 4868 17732 4924
rect 17732 4868 17736 4924
rect 17672 4864 17736 4868
rect 17752 4924 17816 4928
rect 17752 4868 17756 4924
rect 17756 4868 17812 4924
rect 17812 4868 17816 4924
rect 17752 4864 17816 4868
rect 17832 4924 17896 4928
rect 17832 4868 17836 4924
rect 17836 4868 17892 4924
rect 17892 4868 17896 4924
rect 17832 4864 17896 4868
rect 17912 4924 17976 4928
rect 17912 4868 17916 4924
rect 17916 4868 17972 4924
rect 17972 4868 17976 4924
rect 17912 4864 17976 4868
rect 17992 4924 18056 4928
rect 17992 4868 17996 4924
rect 17996 4868 18052 4924
rect 18052 4868 18056 4924
rect 17992 4864 18056 4868
rect 18072 4924 18136 4928
rect 18072 4868 18076 4924
rect 18076 4868 18132 4924
rect 18132 4868 18136 4924
rect 18072 4864 18136 4868
rect 18152 4924 18216 4928
rect 18152 4868 18156 4924
rect 18156 4868 18212 4924
rect 18212 4868 18216 4924
rect 18152 4864 18216 4868
rect 18232 4924 18296 4928
rect 18232 4868 18236 4924
rect 18236 4868 18292 4924
rect 18292 4868 18296 4924
rect 18232 4864 18296 4868
rect 18312 4924 18376 4928
rect 18312 4868 18316 4924
rect 18316 4868 18372 4924
rect 18372 4868 18376 4924
rect 18312 4864 18376 4868
rect 18392 4924 18456 4928
rect 18392 4868 18396 4924
rect 18396 4868 18452 4924
rect 18452 4868 18456 4924
rect 18392 4864 18456 4868
rect 18472 4924 18536 4928
rect 18472 4868 18476 4924
rect 18476 4868 18532 4924
rect 18532 4868 18536 4924
rect 18472 4864 18536 4868
rect 18552 4924 18616 4928
rect 18552 4868 18556 4924
rect 18556 4868 18612 4924
rect 18612 4868 18616 4924
rect 18552 4864 18616 4868
rect 18632 4924 18696 4928
rect 18632 4868 18636 4924
rect 18636 4868 18692 4924
rect 18692 4868 18696 4924
rect 18632 4864 18696 4868
rect 19196 4524 19260 4588
rect 5512 4380 5576 4384
rect 5512 4324 5516 4380
rect 5516 4324 5572 4380
rect 5572 4324 5576 4380
rect 5512 4320 5576 4324
rect 5592 4380 5656 4384
rect 5592 4324 5596 4380
rect 5596 4324 5652 4380
rect 5652 4324 5656 4380
rect 5592 4320 5656 4324
rect 5672 4380 5736 4384
rect 5672 4324 5676 4380
rect 5676 4324 5732 4380
rect 5732 4324 5736 4380
rect 5672 4320 5736 4324
rect 5752 4380 5816 4384
rect 5752 4324 5756 4380
rect 5756 4324 5812 4380
rect 5812 4324 5816 4380
rect 5752 4320 5816 4324
rect 5832 4380 5896 4384
rect 5832 4324 5836 4380
rect 5836 4324 5892 4380
rect 5892 4324 5896 4380
rect 5832 4320 5896 4324
rect 5912 4380 5976 4384
rect 5912 4324 5916 4380
rect 5916 4324 5972 4380
rect 5972 4324 5976 4380
rect 5912 4320 5976 4324
rect 5992 4380 6056 4384
rect 5992 4324 5996 4380
rect 5996 4324 6052 4380
rect 6052 4324 6056 4380
rect 5992 4320 6056 4324
rect 6072 4380 6136 4384
rect 6072 4324 6076 4380
rect 6076 4324 6132 4380
rect 6132 4324 6136 4380
rect 6072 4320 6136 4324
rect 6152 4380 6216 4384
rect 6152 4324 6156 4380
rect 6156 4324 6212 4380
rect 6212 4324 6216 4380
rect 6152 4320 6216 4324
rect 6232 4380 6296 4384
rect 6232 4324 6236 4380
rect 6236 4324 6292 4380
rect 6292 4324 6296 4380
rect 6232 4320 6296 4324
rect 6312 4380 6376 4384
rect 6312 4324 6316 4380
rect 6316 4324 6372 4380
rect 6372 4324 6376 4380
rect 6312 4320 6376 4324
rect 6392 4380 6456 4384
rect 6392 4324 6396 4380
rect 6396 4324 6452 4380
rect 6452 4324 6456 4380
rect 6392 4320 6456 4324
rect 6472 4380 6536 4384
rect 6472 4324 6476 4380
rect 6476 4324 6532 4380
rect 6532 4324 6536 4380
rect 6472 4320 6536 4324
rect 6552 4380 6616 4384
rect 6552 4324 6556 4380
rect 6556 4324 6612 4380
rect 6612 4324 6616 4380
rect 6552 4320 6616 4324
rect 6632 4380 6696 4384
rect 6632 4324 6636 4380
rect 6636 4324 6692 4380
rect 6692 4324 6696 4380
rect 6632 4320 6696 4324
rect 13512 4380 13576 4384
rect 13512 4324 13516 4380
rect 13516 4324 13572 4380
rect 13572 4324 13576 4380
rect 13512 4320 13576 4324
rect 13592 4380 13656 4384
rect 13592 4324 13596 4380
rect 13596 4324 13652 4380
rect 13652 4324 13656 4380
rect 13592 4320 13656 4324
rect 13672 4380 13736 4384
rect 13672 4324 13676 4380
rect 13676 4324 13732 4380
rect 13732 4324 13736 4380
rect 13672 4320 13736 4324
rect 13752 4380 13816 4384
rect 13752 4324 13756 4380
rect 13756 4324 13812 4380
rect 13812 4324 13816 4380
rect 13752 4320 13816 4324
rect 13832 4380 13896 4384
rect 13832 4324 13836 4380
rect 13836 4324 13892 4380
rect 13892 4324 13896 4380
rect 13832 4320 13896 4324
rect 13912 4380 13976 4384
rect 13912 4324 13916 4380
rect 13916 4324 13972 4380
rect 13972 4324 13976 4380
rect 13912 4320 13976 4324
rect 13992 4380 14056 4384
rect 13992 4324 13996 4380
rect 13996 4324 14052 4380
rect 14052 4324 14056 4380
rect 13992 4320 14056 4324
rect 14072 4380 14136 4384
rect 14072 4324 14076 4380
rect 14076 4324 14132 4380
rect 14132 4324 14136 4380
rect 14072 4320 14136 4324
rect 14152 4380 14216 4384
rect 14152 4324 14156 4380
rect 14156 4324 14212 4380
rect 14212 4324 14216 4380
rect 14152 4320 14216 4324
rect 14232 4380 14296 4384
rect 14232 4324 14236 4380
rect 14236 4324 14292 4380
rect 14292 4324 14296 4380
rect 14232 4320 14296 4324
rect 14312 4380 14376 4384
rect 14312 4324 14316 4380
rect 14316 4324 14372 4380
rect 14372 4324 14376 4380
rect 14312 4320 14376 4324
rect 14392 4380 14456 4384
rect 14392 4324 14396 4380
rect 14396 4324 14452 4380
rect 14452 4324 14456 4380
rect 14392 4320 14456 4324
rect 14472 4380 14536 4384
rect 14472 4324 14476 4380
rect 14476 4324 14532 4380
rect 14532 4324 14536 4380
rect 14472 4320 14536 4324
rect 14552 4380 14616 4384
rect 14552 4324 14556 4380
rect 14556 4324 14612 4380
rect 14612 4324 14616 4380
rect 14552 4320 14616 4324
rect 14632 4380 14696 4384
rect 14632 4324 14636 4380
rect 14636 4324 14692 4380
rect 14692 4324 14696 4380
rect 14632 4320 14696 4324
rect 19012 4116 19076 4180
rect 1512 3836 1576 3840
rect 1512 3780 1516 3836
rect 1516 3780 1572 3836
rect 1572 3780 1576 3836
rect 1512 3776 1576 3780
rect 1592 3836 1656 3840
rect 1592 3780 1596 3836
rect 1596 3780 1652 3836
rect 1652 3780 1656 3836
rect 1592 3776 1656 3780
rect 1672 3836 1736 3840
rect 1672 3780 1676 3836
rect 1676 3780 1732 3836
rect 1732 3780 1736 3836
rect 1672 3776 1736 3780
rect 1752 3836 1816 3840
rect 1752 3780 1756 3836
rect 1756 3780 1812 3836
rect 1812 3780 1816 3836
rect 1752 3776 1816 3780
rect 1832 3836 1896 3840
rect 1832 3780 1836 3836
rect 1836 3780 1892 3836
rect 1892 3780 1896 3836
rect 1832 3776 1896 3780
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 2312 3836 2376 3840
rect 2312 3780 2316 3836
rect 2316 3780 2372 3836
rect 2372 3780 2376 3836
rect 2312 3776 2376 3780
rect 2392 3836 2456 3840
rect 2392 3780 2396 3836
rect 2396 3780 2452 3836
rect 2452 3780 2456 3836
rect 2392 3776 2456 3780
rect 2472 3836 2536 3840
rect 2472 3780 2476 3836
rect 2476 3780 2532 3836
rect 2532 3780 2536 3836
rect 2472 3776 2536 3780
rect 2552 3836 2616 3840
rect 2552 3780 2556 3836
rect 2556 3780 2612 3836
rect 2612 3780 2616 3836
rect 2552 3776 2616 3780
rect 2632 3836 2696 3840
rect 2632 3780 2636 3836
rect 2636 3780 2692 3836
rect 2692 3780 2696 3836
rect 2632 3776 2696 3780
rect 9512 3836 9576 3840
rect 9512 3780 9516 3836
rect 9516 3780 9572 3836
rect 9572 3780 9576 3836
rect 9512 3776 9576 3780
rect 9592 3836 9656 3840
rect 9592 3780 9596 3836
rect 9596 3780 9652 3836
rect 9652 3780 9656 3836
rect 9592 3776 9656 3780
rect 9672 3836 9736 3840
rect 9672 3780 9676 3836
rect 9676 3780 9732 3836
rect 9732 3780 9736 3836
rect 9672 3776 9736 3780
rect 9752 3836 9816 3840
rect 9752 3780 9756 3836
rect 9756 3780 9812 3836
rect 9812 3780 9816 3836
rect 9752 3776 9816 3780
rect 9832 3836 9896 3840
rect 9832 3780 9836 3836
rect 9836 3780 9892 3836
rect 9892 3780 9896 3836
rect 9832 3776 9896 3780
rect 9912 3836 9976 3840
rect 9912 3780 9916 3836
rect 9916 3780 9972 3836
rect 9972 3780 9976 3836
rect 9912 3776 9976 3780
rect 9992 3836 10056 3840
rect 9992 3780 9996 3836
rect 9996 3780 10052 3836
rect 10052 3780 10056 3836
rect 9992 3776 10056 3780
rect 10072 3836 10136 3840
rect 10072 3780 10076 3836
rect 10076 3780 10132 3836
rect 10132 3780 10136 3836
rect 10072 3776 10136 3780
rect 10152 3836 10216 3840
rect 10152 3780 10156 3836
rect 10156 3780 10212 3836
rect 10212 3780 10216 3836
rect 10152 3776 10216 3780
rect 10232 3836 10296 3840
rect 10232 3780 10236 3836
rect 10236 3780 10292 3836
rect 10292 3780 10296 3836
rect 10232 3776 10296 3780
rect 10312 3836 10376 3840
rect 10312 3780 10316 3836
rect 10316 3780 10372 3836
rect 10372 3780 10376 3836
rect 10312 3776 10376 3780
rect 10392 3836 10456 3840
rect 10392 3780 10396 3836
rect 10396 3780 10452 3836
rect 10452 3780 10456 3836
rect 10392 3776 10456 3780
rect 10472 3836 10536 3840
rect 10472 3780 10476 3836
rect 10476 3780 10532 3836
rect 10532 3780 10536 3836
rect 10472 3776 10536 3780
rect 10552 3836 10616 3840
rect 10552 3780 10556 3836
rect 10556 3780 10612 3836
rect 10612 3780 10616 3836
rect 10552 3776 10616 3780
rect 10632 3836 10696 3840
rect 10632 3780 10636 3836
rect 10636 3780 10692 3836
rect 10692 3780 10696 3836
rect 10632 3776 10696 3780
rect 17512 3836 17576 3840
rect 17512 3780 17516 3836
rect 17516 3780 17572 3836
rect 17572 3780 17576 3836
rect 17512 3776 17576 3780
rect 17592 3836 17656 3840
rect 17592 3780 17596 3836
rect 17596 3780 17652 3836
rect 17652 3780 17656 3836
rect 17592 3776 17656 3780
rect 17672 3836 17736 3840
rect 17672 3780 17676 3836
rect 17676 3780 17732 3836
rect 17732 3780 17736 3836
rect 17672 3776 17736 3780
rect 17752 3836 17816 3840
rect 17752 3780 17756 3836
rect 17756 3780 17812 3836
rect 17812 3780 17816 3836
rect 17752 3776 17816 3780
rect 17832 3836 17896 3840
rect 17832 3780 17836 3836
rect 17836 3780 17892 3836
rect 17892 3780 17896 3836
rect 17832 3776 17896 3780
rect 17912 3836 17976 3840
rect 17912 3780 17916 3836
rect 17916 3780 17972 3836
rect 17972 3780 17976 3836
rect 17912 3776 17976 3780
rect 17992 3836 18056 3840
rect 17992 3780 17996 3836
rect 17996 3780 18052 3836
rect 18052 3780 18056 3836
rect 17992 3776 18056 3780
rect 18072 3836 18136 3840
rect 18072 3780 18076 3836
rect 18076 3780 18132 3836
rect 18132 3780 18136 3836
rect 18072 3776 18136 3780
rect 18152 3836 18216 3840
rect 18152 3780 18156 3836
rect 18156 3780 18212 3836
rect 18212 3780 18216 3836
rect 18152 3776 18216 3780
rect 18232 3836 18296 3840
rect 18232 3780 18236 3836
rect 18236 3780 18292 3836
rect 18292 3780 18296 3836
rect 18232 3776 18296 3780
rect 18312 3836 18376 3840
rect 18312 3780 18316 3836
rect 18316 3780 18372 3836
rect 18372 3780 18376 3836
rect 18312 3776 18376 3780
rect 18392 3836 18456 3840
rect 18392 3780 18396 3836
rect 18396 3780 18452 3836
rect 18452 3780 18456 3836
rect 18392 3776 18456 3780
rect 18472 3836 18536 3840
rect 18472 3780 18476 3836
rect 18476 3780 18532 3836
rect 18532 3780 18536 3836
rect 18472 3776 18536 3780
rect 18552 3836 18616 3840
rect 18552 3780 18556 3836
rect 18556 3780 18612 3836
rect 18612 3780 18616 3836
rect 18552 3776 18616 3780
rect 18632 3836 18696 3840
rect 18632 3780 18636 3836
rect 18636 3780 18692 3836
rect 18692 3780 18696 3836
rect 18632 3776 18696 3780
rect 5512 3292 5576 3296
rect 5512 3236 5516 3292
rect 5516 3236 5572 3292
rect 5572 3236 5576 3292
rect 5512 3232 5576 3236
rect 5592 3292 5656 3296
rect 5592 3236 5596 3292
rect 5596 3236 5652 3292
rect 5652 3236 5656 3292
rect 5592 3232 5656 3236
rect 5672 3292 5736 3296
rect 5672 3236 5676 3292
rect 5676 3236 5732 3292
rect 5732 3236 5736 3292
rect 5672 3232 5736 3236
rect 5752 3292 5816 3296
rect 5752 3236 5756 3292
rect 5756 3236 5812 3292
rect 5812 3236 5816 3292
rect 5752 3232 5816 3236
rect 5832 3292 5896 3296
rect 5832 3236 5836 3292
rect 5836 3236 5892 3292
rect 5892 3236 5896 3292
rect 5832 3232 5896 3236
rect 5912 3292 5976 3296
rect 5912 3236 5916 3292
rect 5916 3236 5972 3292
rect 5972 3236 5976 3292
rect 5912 3232 5976 3236
rect 5992 3292 6056 3296
rect 5992 3236 5996 3292
rect 5996 3236 6052 3292
rect 6052 3236 6056 3292
rect 5992 3232 6056 3236
rect 6072 3292 6136 3296
rect 6072 3236 6076 3292
rect 6076 3236 6132 3292
rect 6132 3236 6136 3292
rect 6072 3232 6136 3236
rect 6152 3292 6216 3296
rect 6152 3236 6156 3292
rect 6156 3236 6212 3292
rect 6212 3236 6216 3292
rect 6152 3232 6216 3236
rect 6232 3292 6296 3296
rect 6232 3236 6236 3292
rect 6236 3236 6292 3292
rect 6292 3236 6296 3292
rect 6232 3232 6296 3236
rect 6312 3292 6376 3296
rect 6312 3236 6316 3292
rect 6316 3236 6372 3292
rect 6372 3236 6376 3292
rect 6312 3232 6376 3236
rect 6392 3292 6456 3296
rect 6392 3236 6396 3292
rect 6396 3236 6452 3292
rect 6452 3236 6456 3292
rect 6392 3232 6456 3236
rect 6472 3292 6536 3296
rect 6472 3236 6476 3292
rect 6476 3236 6532 3292
rect 6532 3236 6536 3292
rect 6472 3232 6536 3236
rect 6552 3292 6616 3296
rect 6552 3236 6556 3292
rect 6556 3236 6612 3292
rect 6612 3236 6616 3292
rect 6552 3232 6616 3236
rect 6632 3292 6696 3296
rect 6632 3236 6636 3292
rect 6636 3236 6692 3292
rect 6692 3236 6696 3292
rect 6632 3232 6696 3236
rect 13512 3292 13576 3296
rect 13512 3236 13516 3292
rect 13516 3236 13572 3292
rect 13572 3236 13576 3292
rect 13512 3232 13576 3236
rect 13592 3292 13656 3296
rect 13592 3236 13596 3292
rect 13596 3236 13652 3292
rect 13652 3236 13656 3292
rect 13592 3232 13656 3236
rect 13672 3292 13736 3296
rect 13672 3236 13676 3292
rect 13676 3236 13732 3292
rect 13732 3236 13736 3292
rect 13672 3232 13736 3236
rect 13752 3292 13816 3296
rect 13752 3236 13756 3292
rect 13756 3236 13812 3292
rect 13812 3236 13816 3292
rect 13752 3232 13816 3236
rect 13832 3292 13896 3296
rect 13832 3236 13836 3292
rect 13836 3236 13892 3292
rect 13892 3236 13896 3292
rect 13832 3232 13896 3236
rect 13912 3292 13976 3296
rect 13912 3236 13916 3292
rect 13916 3236 13972 3292
rect 13972 3236 13976 3292
rect 13912 3232 13976 3236
rect 13992 3292 14056 3296
rect 13992 3236 13996 3292
rect 13996 3236 14052 3292
rect 14052 3236 14056 3292
rect 13992 3232 14056 3236
rect 14072 3292 14136 3296
rect 14072 3236 14076 3292
rect 14076 3236 14132 3292
rect 14132 3236 14136 3292
rect 14072 3232 14136 3236
rect 14152 3292 14216 3296
rect 14152 3236 14156 3292
rect 14156 3236 14212 3292
rect 14212 3236 14216 3292
rect 14152 3232 14216 3236
rect 14232 3292 14296 3296
rect 14232 3236 14236 3292
rect 14236 3236 14292 3292
rect 14292 3236 14296 3292
rect 14232 3232 14296 3236
rect 14312 3292 14376 3296
rect 14312 3236 14316 3292
rect 14316 3236 14372 3292
rect 14372 3236 14376 3292
rect 14312 3232 14376 3236
rect 14392 3292 14456 3296
rect 14392 3236 14396 3292
rect 14396 3236 14452 3292
rect 14452 3236 14456 3292
rect 14392 3232 14456 3236
rect 14472 3292 14536 3296
rect 14472 3236 14476 3292
rect 14476 3236 14532 3292
rect 14532 3236 14536 3292
rect 14472 3232 14536 3236
rect 14552 3292 14616 3296
rect 14552 3236 14556 3292
rect 14556 3236 14612 3292
rect 14612 3236 14616 3292
rect 14552 3232 14616 3236
rect 14632 3292 14696 3296
rect 14632 3236 14636 3292
rect 14636 3236 14692 3292
rect 14692 3236 14696 3292
rect 14632 3232 14696 3236
rect 1512 2748 1576 2752
rect 1512 2692 1516 2748
rect 1516 2692 1572 2748
rect 1572 2692 1576 2748
rect 1512 2688 1576 2692
rect 1592 2748 1656 2752
rect 1592 2692 1596 2748
rect 1596 2692 1652 2748
rect 1652 2692 1656 2748
rect 1592 2688 1656 2692
rect 1672 2748 1736 2752
rect 1672 2692 1676 2748
rect 1676 2692 1732 2748
rect 1732 2692 1736 2748
rect 1672 2688 1736 2692
rect 1752 2748 1816 2752
rect 1752 2692 1756 2748
rect 1756 2692 1812 2748
rect 1812 2692 1816 2748
rect 1752 2688 1816 2692
rect 1832 2748 1896 2752
rect 1832 2692 1836 2748
rect 1836 2692 1892 2748
rect 1892 2692 1896 2748
rect 1832 2688 1896 2692
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 2312 2748 2376 2752
rect 2312 2692 2316 2748
rect 2316 2692 2372 2748
rect 2372 2692 2376 2748
rect 2312 2688 2376 2692
rect 2392 2748 2456 2752
rect 2392 2692 2396 2748
rect 2396 2692 2452 2748
rect 2452 2692 2456 2748
rect 2392 2688 2456 2692
rect 2472 2748 2536 2752
rect 2472 2692 2476 2748
rect 2476 2692 2532 2748
rect 2532 2692 2536 2748
rect 2472 2688 2536 2692
rect 2552 2748 2616 2752
rect 2552 2692 2556 2748
rect 2556 2692 2612 2748
rect 2612 2692 2616 2748
rect 2552 2688 2616 2692
rect 2632 2748 2696 2752
rect 2632 2692 2636 2748
rect 2636 2692 2692 2748
rect 2692 2692 2696 2748
rect 2632 2688 2696 2692
rect 9512 2748 9576 2752
rect 9512 2692 9516 2748
rect 9516 2692 9572 2748
rect 9572 2692 9576 2748
rect 9512 2688 9576 2692
rect 9592 2748 9656 2752
rect 9592 2692 9596 2748
rect 9596 2692 9652 2748
rect 9652 2692 9656 2748
rect 9592 2688 9656 2692
rect 9672 2748 9736 2752
rect 9672 2692 9676 2748
rect 9676 2692 9732 2748
rect 9732 2692 9736 2748
rect 9672 2688 9736 2692
rect 9752 2748 9816 2752
rect 9752 2692 9756 2748
rect 9756 2692 9812 2748
rect 9812 2692 9816 2748
rect 9752 2688 9816 2692
rect 9832 2748 9896 2752
rect 9832 2692 9836 2748
rect 9836 2692 9892 2748
rect 9892 2692 9896 2748
rect 9832 2688 9896 2692
rect 9912 2748 9976 2752
rect 9912 2692 9916 2748
rect 9916 2692 9972 2748
rect 9972 2692 9976 2748
rect 9912 2688 9976 2692
rect 9992 2748 10056 2752
rect 9992 2692 9996 2748
rect 9996 2692 10052 2748
rect 10052 2692 10056 2748
rect 9992 2688 10056 2692
rect 10072 2748 10136 2752
rect 10072 2692 10076 2748
rect 10076 2692 10132 2748
rect 10132 2692 10136 2748
rect 10072 2688 10136 2692
rect 10152 2748 10216 2752
rect 10152 2692 10156 2748
rect 10156 2692 10212 2748
rect 10212 2692 10216 2748
rect 10152 2688 10216 2692
rect 10232 2748 10296 2752
rect 10232 2692 10236 2748
rect 10236 2692 10292 2748
rect 10292 2692 10296 2748
rect 10232 2688 10296 2692
rect 10312 2748 10376 2752
rect 10312 2692 10316 2748
rect 10316 2692 10372 2748
rect 10372 2692 10376 2748
rect 10312 2688 10376 2692
rect 10392 2748 10456 2752
rect 10392 2692 10396 2748
rect 10396 2692 10452 2748
rect 10452 2692 10456 2748
rect 10392 2688 10456 2692
rect 10472 2748 10536 2752
rect 10472 2692 10476 2748
rect 10476 2692 10532 2748
rect 10532 2692 10536 2748
rect 10472 2688 10536 2692
rect 10552 2748 10616 2752
rect 10552 2692 10556 2748
rect 10556 2692 10612 2748
rect 10612 2692 10616 2748
rect 10552 2688 10616 2692
rect 10632 2748 10696 2752
rect 10632 2692 10636 2748
rect 10636 2692 10692 2748
rect 10692 2692 10696 2748
rect 10632 2688 10696 2692
rect 17512 2748 17576 2752
rect 17512 2692 17516 2748
rect 17516 2692 17572 2748
rect 17572 2692 17576 2748
rect 17512 2688 17576 2692
rect 17592 2748 17656 2752
rect 17592 2692 17596 2748
rect 17596 2692 17652 2748
rect 17652 2692 17656 2748
rect 17592 2688 17656 2692
rect 17672 2748 17736 2752
rect 17672 2692 17676 2748
rect 17676 2692 17732 2748
rect 17732 2692 17736 2748
rect 17672 2688 17736 2692
rect 17752 2748 17816 2752
rect 17752 2692 17756 2748
rect 17756 2692 17812 2748
rect 17812 2692 17816 2748
rect 17752 2688 17816 2692
rect 17832 2748 17896 2752
rect 17832 2692 17836 2748
rect 17836 2692 17892 2748
rect 17892 2692 17896 2748
rect 17832 2688 17896 2692
rect 17912 2748 17976 2752
rect 17912 2692 17916 2748
rect 17916 2692 17972 2748
rect 17972 2692 17976 2748
rect 17912 2688 17976 2692
rect 17992 2748 18056 2752
rect 17992 2692 17996 2748
rect 17996 2692 18052 2748
rect 18052 2692 18056 2748
rect 17992 2688 18056 2692
rect 18072 2748 18136 2752
rect 18072 2692 18076 2748
rect 18076 2692 18132 2748
rect 18132 2692 18136 2748
rect 18072 2688 18136 2692
rect 18152 2748 18216 2752
rect 18152 2692 18156 2748
rect 18156 2692 18212 2748
rect 18212 2692 18216 2748
rect 18152 2688 18216 2692
rect 18232 2748 18296 2752
rect 18232 2692 18236 2748
rect 18236 2692 18292 2748
rect 18292 2692 18296 2748
rect 18232 2688 18296 2692
rect 18312 2748 18376 2752
rect 18312 2692 18316 2748
rect 18316 2692 18372 2748
rect 18372 2692 18376 2748
rect 18312 2688 18376 2692
rect 18392 2748 18456 2752
rect 18392 2692 18396 2748
rect 18396 2692 18452 2748
rect 18452 2692 18456 2748
rect 18392 2688 18456 2692
rect 18472 2748 18536 2752
rect 18472 2692 18476 2748
rect 18476 2692 18532 2748
rect 18532 2692 18536 2748
rect 18472 2688 18536 2692
rect 18552 2748 18616 2752
rect 18552 2692 18556 2748
rect 18556 2692 18612 2748
rect 18612 2692 18616 2748
rect 18552 2688 18616 2692
rect 18632 2748 18696 2752
rect 18632 2692 18636 2748
rect 18636 2692 18692 2748
rect 18692 2692 18696 2748
rect 18632 2688 18696 2692
rect 5512 2204 5576 2208
rect 5512 2148 5516 2204
rect 5516 2148 5572 2204
rect 5572 2148 5576 2204
rect 5512 2144 5576 2148
rect 5592 2204 5656 2208
rect 5592 2148 5596 2204
rect 5596 2148 5652 2204
rect 5652 2148 5656 2204
rect 5592 2144 5656 2148
rect 5672 2204 5736 2208
rect 5672 2148 5676 2204
rect 5676 2148 5732 2204
rect 5732 2148 5736 2204
rect 5672 2144 5736 2148
rect 5752 2204 5816 2208
rect 5752 2148 5756 2204
rect 5756 2148 5812 2204
rect 5812 2148 5816 2204
rect 5752 2144 5816 2148
rect 5832 2204 5896 2208
rect 5832 2148 5836 2204
rect 5836 2148 5892 2204
rect 5892 2148 5896 2204
rect 5832 2144 5896 2148
rect 5912 2204 5976 2208
rect 5912 2148 5916 2204
rect 5916 2148 5972 2204
rect 5972 2148 5976 2204
rect 5912 2144 5976 2148
rect 5992 2204 6056 2208
rect 5992 2148 5996 2204
rect 5996 2148 6052 2204
rect 6052 2148 6056 2204
rect 5992 2144 6056 2148
rect 6072 2204 6136 2208
rect 6072 2148 6076 2204
rect 6076 2148 6132 2204
rect 6132 2148 6136 2204
rect 6072 2144 6136 2148
rect 6152 2204 6216 2208
rect 6152 2148 6156 2204
rect 6156 2148 6212 2204
rect 6212 2148 6216 2204
rect 6152 2144 6216 2148
rect 6232 2204 6296 2208
rect 6232 2148 6236 2204
rect 6236 2148 6292 2204
rect 6292 2148 6296 2204
rect 6232 2144 6296 2148
rect 6312 2204 6376 2208
rect 6312 2148 6316 2204
rect 6316 2148 6372 2204
rect 6372 2148 6376 2204
rect 6312 2144 6376 2148
rect 6392 2204 6456 2208
rect 6392 2148 6396 2204
rect 6396 2148 6452 2204
rect 6452 2148 6456 2204
rect 6392 2144 6456 2148
rect 6472 2204 6536 2208
rect 6472 2148 6476 2204
rect 6476 2148 6532 2204
rect 6532 2148 6536 2204
rect 6472 2144 6536 2148
rect 6552 2204 6616 2208
rect 6552 2148 6556 2204
rect 6556 2148 6612 2204
rect 6612 2148 6616 2204
rect 6552 2144 6616 2148
rect 6632 2204 6696 2208
rect 6632 2148 6636 2204
rect 6636 2148 6692 2204
rect 6692 2148 6696 2204
rect 6632 2144 6696 2148
rect 13512 2204 13576 2208
rect 13512 2148 13516 2204
rect 13516 2148 13572 2204
rect 13572 2148 13576 2204
rect 13512 2144 13576 2148
rect 13592 2204 13656 2208
rect 13592 2148 13596 2204
rect 13596 2148 13652 2204
rect 13652 2148 13656 2204
rect 13592 2144 13656 2148
rect 13672 2204 13736 2208
rect 13672 2148 13676 2204
rect 13676 2148 13732 2204
rect 13732 2148 13736 2204
rect 13672 2144 13736 2148
rect 13752 2204 13816 2208
rect 13752 2148 13756 2204
rect 13756 2148 13812 2204
rect 13812 2148 13816 2204
rect 13752 2144 13816 2148
rect 13832 2204 13896 2208
rect 13832 2148 13836 2204
rect 13836 2148 13892 2204
rect 13892 2148 13896 2204
rect 13832 2144 13896 2148
rect 13912 2204 13976 2208
rect 13912 2148 13916 2204
rect 13916 2148 13972 2204
rect 13972 2148 13976 2204
rect 13912 2144 13976 2148
rect 13992 2204 14056 2208
rect 13992 2148 13996 2204
rect 13996 2148 14052 2204
rect 14052 2148 14056 2204
rect 13992 2144 14056 2148
rect 14072 2204 14136 2208
rect 14072 2148 14076 2204
rect 14076 2148 14132 2204
rect 14132 2148 14136 2204
rect 14072 2144 14136 2148
rect 14152 2204 14216 2208
rect 14152 2148 14156 2204
rect 14156 2148 14212 2204
rect 14212 2148 14216 2204
rect 14152 2144 14216 2148
rect 14232 2204 14296 2208
rect 14232 2148 14236 2204
rect 14236 2148 14292 2204
rect 14292 2148 14296 2204
rect 14232 2144 14296 2148
rect 14312 2204 14376 2208
rect 14312 2148 14316 2204
rect 14316 2148 14372 2204
rect 14372 2148 14376 2204
rect 14312 2144 14376 2148
rect 14392 2204 14456 2208
rect 14392 2148 14396 2204
rect 14396 2148 14452 2204
rect 14452 2148 14456 2204
rect 14392 2144 14456 2148
rect 14472 2204 14536 2208
rect 14472 2148 14476 2204
rect 14476 2148 14532 2204
rect 14532 2148 14536 2204
rect 14472 2144 14536 2148
rect 14552 2204 14616 2208
rect 14552 2148 14556 2204
rect 14556 2148 14612 2204
rect 14612 2148 14616 2204
rect 14552 2144 14616 2148
rect 14632 2204 14696 2208
rect 14632 2148 14636 2204
rect 14636 2148 14692 2204
rect 14692 2148 14696 2204
rect 14632 2144 14696 2148
<< metal4 >>
rect 1484 16896 2724 17456
rect 1484 16832 1512 16896
rect 1576 16832 1592 16896
rect 1656 16832 1672 16896
rect 1736 16832 1752 16896
rect 1816 16832 1832 16896
rect 1896 16832 1912 16896
rect 1976 16832 1992 16896
rect 2056 16832 2072 16896
rect 2136 16832 2152 16896
rect 2216 16832 2232 16896
rect 2296 16832 2312 16896
rect 2376 16832 2392 16896
rect 2456 16832 2472 16896
rect 2536 16832 2552 16896
rect 2616 16832 2632 16896
rect 2696 16832 2724 16896
rect 1484 15808 2724 16832
rect 1484 15744 1512 15808
rect 1576 15744 1592 15808
rect 1656 15744 1672 15808
rect 1736 15744 1752 15808
rect 1816 15744 1832 15808
rect 1896 15744 1912 15808
rect 1976 15744 1992 15808
rect 2056 15744 2072 15808
rect 2136 15744 2152 15808
rect 2216 15744 2232 15808
rect 2296 15744 2312 15808
rect 2376 15744 2392 15808
rect 2456 15744 2472 15808
rect 2536 15744 2552 15808
rect 2616 15744 2632 15808
rect 2696 15744 2724 15808
rect 1484 14720 2724 15744
rect 1484 14656 1512 14720
rect 1576 14656 1592 14720
rect 1656 14656 1672 14720
rect 1736 14656 1752 14720
rect 1816 14656 1832 14720
rect 1896 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2312 14720
rect 2376 14656 2392 14720
rect 2456 14656 2472 14720
rect 2536 14656 2552 14720
rect 2616 14656 2632 14720
rect 2696 14656 2724 14720
rect 1484 13632 2724 14656
rect 1484 13568 1512 13632
rect 1576 13568 1592 13632
rect 1656 13568 1672 13632
rect 1736 13568 1752 13632
rect 1816 13568 1832 13632
rect 1896 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2312 13632
rect 2376 13568 2392 13632
rect 2456 13568 2472 13632
rect 2536 13568 2552 13632
rect 2616 13568 2632 13632
rect 2696 13568 2724 13632
rect 1484 12544 2724 13568
rect 1484 12480 1512 12544
rect 1576 12480 1592 12544
rect 1656 12480 1672 12544
rect 1736 12480 1752 12544
rect 1816 12480 1832 12544
rect 1896 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2312 12544
rect 2376 12480 2392 12544
rect 2456 12480 2472 12544
rect 2536 12480 2552 12544
rect 2616 12480 2632 12544
rect 2696 12480 2724 12544
rect 1484 11456 2724 12480
rect 1484 11392 1512 11456
rect 1576 11392 1592 11456
rect 1656 11392 1672 11456
rect 1736 11392 1752 11456
rect 1816 11392 1832 11456
rect 1896 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2312 11456
rect 2376 11392 2392 11456
rect 2456 11392 2472 11456
rect 2536 11392 2552 11456
rect 2616 11392 2632 11456
rect 2696 11392 2724 11456
rect 1484 10368 2724 11392
rect 1484 10304 1512 10368
rect 1576 10304 1592 10368
rect 1656 10304 1672 10368
rect 1736 10304 1752 10368
rect 1816 10304 1832 10368
rect 1896 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2312 10368
rect 2376 10304 2392 10368
rect 2456 10304 2472 10368
rect 2536 10304 2552 10368
rect 2616 10304 2632 10368
rect 2696 10304 2724 10368
rect 1484 9280 2724 10304
rect 1484 9216 1512 9280
rect 1576 9216 1592 9280
rect 1656 9216 1672 9280
rect 1736 9216 1752 9280
rect 1816 9216 1832 9280
rect 1896 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2312 9280
rect 2376 9216 2392 9280
rect 2456 9216 2472 9280
rect 2536 9216 2552 9280
rect 2616 9216 2632 9280
rect 2696 9216 2724 9280
rect 1484 8192 2724 9216
rect 1484 8128 1512 8192
rect 1576 8128 1592 8192
rect 1656 8128 1672 8192
rect 1736 8128 1752 8192
rect 1816 8128 1832 8192
rect 1896 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2312 8192
rect 2376 8128 2392 8192
rect 2456 8128 2472 8192
rect 2536 8128 2552 8192
rect 2616 8128 2632 8192
rect 2696 8128 2724 8192
rect 1484 7104 2724 8128
rect 1484 7040 1512 7104
rect 1576 7040 1592 7104
rect 1656 7040 1672 7104
rect 1736 7040 1752 7104
rect 1816 7040 1832 7104
rect 1896 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2312 7104
rect 2376 7040 2392 7104
rect 2456 7040 2472 7104
rect 2536 7040 2552 7104
rect 2616 7040 2632 7104
rect 2696 7040 2724 7104
rect 1484 6016 2724 7040
rect 1484 5952 1512 6016
rect 1576 5952 1592 6016
rect 1656 5952 1672 6016
rect 1736 5952 1752 6016
rect 1816 5952 1832 6016
rect 1896 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2312 6016
rect 2376 5952 2392 6016
rect 2456 5952 2472 6016
rect 2536 5952 2552 6016
rect 2616 5952 2632 6016
rect 2696 5952 2724 6016
rect 1484 4928 2724 5952
rect 1484 4864 1512 4928
rect 1576 4864 1592 4928
rect 1656 4864 1672 4928
rect 1736 4864 1752 4928
rect 1816 4864 1832 4928
rect 1896 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2312 4928
rect 2376 4864 2392 4928
rect 2456 4864 2472 4928
rect 2536 4864 2552 4928
rect 2616 4864 2632 4928
rect 2696 4864 2724 4928
rect 1484 3840 2724 4864
rect 1484 3776 1512 3840
rect 1576 3776 1592 3840
rect 1656 3776 1672 3840
rect 1736 3776 1752 3840
rect 1816 3776 1832 3840
rect 1896 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2312 3840
rect 2376 3776 2392 3840
rect 2456 3776 2472 3840
rect 2536 3776 2552 3840
rect 2616 3776 2632 3840
rect 2696 3776 2724 3840
rect 1484 2752 2724 3776
rect 1484 2688 1512 2752
rect 1576 2688 1592 2752
rect 1656 2688 1672 2752
rect 1736 2688 1752 2752
rect 1816 2688 1832 2752
rect 1896 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2312 2752
rect 2376 2688 2392 2752
rect 2456 2688 2472 2752
rect 2536 2688 2552 2752
rect 2616 2688 2632 2752
rect 2696 2688 2724 2752
rect 1484 2128 2724 2688
rect 5484 17440 6724 17456
rect 5484 17376 5512 17440
rect 5576 17376 5592 17440
rect 5656 17376 5672 17440
rect 5736 17376 5752 17440
rect 5816 17376 5832 17440
rect 5896 17376 5912 17440
rect 5976 17376 5992 17440
rect 6056 17376 6072 17440
rect 6136 17376 6152 17440
rect 6216 17376 6232 17440
rect 6296 17376 6312 17440
rect 6376 17376 6392 17440
rect 6456 17376 6472 17440
rect 6536 17376 6552 17440
rect 6616 17376 6632 17440
rect 6696 17376 6724 17440
rect 5484 16352 6724 17376
rect 5484 16288 5512 16352
rect 5576 16288 5592 16352
rect 5656 16288 5672 16352
rect 5736 16288 5752 16352
rect 5816 16288 5832 16352
rect 5896 16288 5912 16352
rect 5976 16288 5992 16352
rect 6056 16288 6072 16352
rect 6136 16288 6152 16352
rect 6216 16288 6232 16352
rect 6296 16288 6312 16352
rect 6376 16288 6392 16352
rect 6456 16288 6472 16352
rect 6536 16288 6552 16352
rect 6616 16288 6632 16352
rect 6696 16288 6724 16352
rect 5484 15264 6724 16288
rect 5484 15200 5512 15264
rect 5576 15200 5592 15264
rect 5656 15200 5672 15264
rect 5736 15200 5752 15264
rect 5816 15200 5832 15264
rect 5896 15200 5912 15264
rect 5976 15200 5992 15264
rect 6056 15200 6072 15264
rect 6136 15200 6152 15264
rect 6216 15200 6232 15264
rect 6296 15200 6312 15264
rect 6376 15200 6392 15264
rect 6456 15200 6472 15264
rect 6536 15200 6552 15264
rect 6616 15200 6632 15264
rect 6696 15200 6724 15264
rect 5484 14176 6724 15200
rect 5484 14112 5512 14176
rect 5576 14112 5592 14176
rect 5656 14112 5672 14176
rect 5736 14112 5752 14176
rect 5816 14112 5832 14176
rect 5896 14112 5912 14176
rect 5976 14112 5992 14176
rect 6056 14112 6072 14176
rect 6136 14112 6152 14176
rect 6216 14112 6232 14176
rect 6296 14112 6312 14176
rect 6376 14112 6392 14176
rect 6456 14112 6472 14176
rect 6536 14112 6552 14176
rect 6616 14112 6632 14176
rect 6696 14112 6724 14176
rect 5484 13088 6724 14112
rect 5484 13024 5512 13088
rect 5576 13024 5592 13088
rect 5656 13024 5672 13088
rect 5736 13024 5752 13088
rect 5816 13024 5832 13088
rect 5896 13024 5912 13088
rect 5976 13024 5992 13088
rect 6056 13024 6072 13088
rect 6136 13024 6152 13088
rect 6216 13024 6232 13088
rect 6296 13024 6312 13088
rect 6376 13024 6392 13088
rect 6456 13024 6472 13088
rect 6536 13024 6552 13088
rect 6616 13024 6632 13088
rect 6696 13024 6724 13088
rect 5484 12000 6724 13024
rect 5484 11936 5512 12000
rect 5576 11936 5592 12000
rect 5656 11936 5672 12000
rect 5736 11936 5752 12000
rect 5816 11936 5832 12000
rect 5896 11936 5912 12000
rect 5976 11936 5992 12000
rect 6056 11936 6072 12000
rect 6136 11936 6152 12000
rect 6216 11936 6232 12000
rect 6296 11936 6312 12000
rect 6376 11936 6392 12000
rect 6456 11936 6472 12000
rect 6536 11936 6552 12000
rect 6616 11936 6632 12000
rect 6696 11936 6724 12000
rect 5484 10912 6724 11936
rect 5484 10848 5512 10912
rect 5576 10848 5592 10912
rect 5656 10848 5672 10912
rect 5736 10848 5752 10912
rect 5816 10848 5832 10912
rect 5896 10848 5912 10912
rect 5976 10848 5992 10912
rect 6056 10848 6072 10912
rect 6136 10848 6152 10912
rect 6216 10848 6232 10912
rect 6296 10848 6312 10912
rect 6376 10848 6392 10912
rect 6456 10848 6472 10912
rect 6536 10848 6552 10912
rect 6616 10848 6632 10912
rect 6696 10848 6724 10912
rect 5484 9824 6724 10848
rect 5484 9760 5512 9824
rect 5576 9760 5592 9824
rect 5656 9760 5672 9824
rect 5736 9760 5752 9824
rect 5816 9760 5832 9824
rect 5896 9760 5912 9824
rect 5976 9760 5992 9824
rect 6056 9760 6072 9824
rect 6136 9760 6152 9824
rect 6216 9760 6232 9824
rect 6296 9760 6312 9824
rect 6376 9760 6392 9824
rect 6456 9760 6472 9824
rect 6536 9760 6552 9824
rect 6616 9760 6632 9824
rect 6696 9760 6724 9824
rect 5484 8736 6724 9760
rect 5484 8672 5512 8736
rect 5576 8672 5592 8736
rect 5656 8672 5672 8736
rect 5736 8672 5752 8736
rect 5816 8672 5832 8736
rect 5896 8672 5912 8736
rect 5976 8672 5992 8736
rect 6056 8672 6072 8736
rect 6136 8672 6152 8736
rect 6216 8672 6232 8736
rect 6296 8672 6312 8736
rect 6376 8672 6392 8736
rect 6456 8672 6472 8736
rect 6536 8672 6552 8736
rect 6616 8672 6632 8736
rect 6696 8672 6724 8736
rect 5484 7648 6724 8672
rect 5484 7584 5512 7648
rect 5576 7584 5592 7648
rect 5656 7584 5672 7648
rect 5736 7584 5752 7648
rect 5816 7584 5832 7648
rect 5896 7584 5912 7648
rect 5976 7584 5992 7648
rect 6056 7584 6072 7648
rect 6136 7584 6152 7648
rect 6216 7584 6232 7648
rect 6296 7584 6312 7648
rect 6376 7584 6392 7648
rect 6456 7584 6472 7648
rect 6536 7584 6552 7648
rect 6616 7584 6632 7648
rect 6696 7584 6724 7648
rect 5484 6560 6724 7584
rect 5484 6496 5512 6560
rect 5576 6496 5592 6560
rect 5656 6496 5672 6560
rect 5736 6496 5752 6560
rect 5816 6496 5832 6560
rect 5896 6496 5912 6560
rect 5976 6496 5992 6560
rect 6056 6496 6072 6560
rect 6136 6496 6152 6560
rect 6216 6496 6232 6560
rect 6296 6496 6312 6560
rect 6376 6496 6392 6560
rect 6456 6496 6472 6560
rect 6536 6496 6552 6560
rect 6616 6496 6632 6560
rect 6696 6496 6724 6560
rect 5484 5472 6724 6496
rect 5484 5408 5512 5472
rect 5576 5408 5592 5472
rect 5656 5408 5672 5472
rect 5736 5408 5752 5472
rect 5816 5408 5832 5472
rect 5896 5408 5912 5472
rect 5976 5408 5992 5472
rect 6056 5408 6072 5472
rect 6136 5408 6152 5472
rect 6216 5408 6232 5472
rect 6296 5408 6312 5472
rect 6376 5408 6392 5472
rect 6456 5408 6472 5472
rect 6536 5408 6552 5472
rect 6616 5408 6632 5472
rect 6696 5408 6724 5472
rect 5484 4384 6724 5408
rect 5484 4320 5512 4384
rect 5576 4320 5592 4384
rect 5656 4320 5672 4384
rect 5736 4320 5752 4384
rect 5816 4320 5832 4384
rect 5896 4320 5912 4384
rect 5976 4320 5992 4384
rect 6056 4320 6072 4384
rect 6136 4320 6152 4384
rect 6216 4320 6232 4384
rect 6296 4320 6312 4384
rect 6376 4320 6392 4384
rect 6456 4320 6472 4384
rect 6536 4320 6552 4384
rect 6616 4320 6632 4384
rect 6696 4320 6724 4384
rect 5484 3296 6724 4320
rect 5484 3232 5512 3296
rect 5576 3232 5592 3296
rect 5656 3232 5672 3296
rect 5736 3232 5752 3296
rect 5816 3232 5832 3296
rect 5896 3232 5912 3296
rect 5976 3232 5992 3296
rect 6056 3232 6072 3296
rect 6136 3232 6152 3296
rect 6216 3232 6232 3296
rect 6296 3232 6312 3296
rect 6376 3232 6392 3296
rect 6456 3232 6472 3296
rect 6536 3232 6552 3296
rect 6616 3232 6632 3296
rect 6696 3232 6724 3296
rect 5484 2208 6724 3232
rect 5484 2144 5512 2208
rect 5576 2144 5592 2208
rect 5656 2144 5672 2208
rect 5736 2144 5752 2208
rect 5816 2144 5832 2208
rect 5896 2144 5912 2208
rect 5976 2144 5992 2208
rect 6056 2144 6072 2208
rect 6136 2144 6152 2208
rect 6216 2144 6232 2208
rect 6296 2144 6312 2208
rect 6376 2144 6392 2208
rect 6456 2144 6472 2208
rect 6536 2144 6552 2208
rect 6616 2144 6632 2208
rect 6696 2144 6724 2208
rect 5484 2128 6724 2144
rect 9484 16896 10724 17456
rect 9484 16832 9512 16896
rect 9576 16832 9592 16896
rect 9656 16832 9672 16896
rect 9736 16832 9752 16896
rect 9816 16832 9832 16896
rect 9896 16832 9912 16896
rect 9976 16832 9992 16896
rect 10056 16832 10072 16896
rect 10136 16832 10152 16896
rect 10216 16832 10232 16896
rect 10296 16832 10312 16896
rect 10376 16832 10392 16896
rect 10456 16832 10472 16896
rect 10536 16832 10552 16896
rect 10616 16832 10632 16896
rect 10696 16832 10724 16896
rect 9484 15808 10724 16832
rect 9484 15744 9512 15808
rect 9576 15744 9592 15808
rect 9656 15744 9672 15808
rect 9736 15744 9752 15808
rect 9816 15744 9832 15808
rect 9896 15744 9912 15808
rect 9976 15744 9992 15808
rect 10056 15744 10072 15808
rect 10136 15744 10152 15808
rect 10216 15744 10232 15808
rect 10296 15744 10312 15808
rect 10376 15744 10392 15808
rect 10456 15744 10472 15808
rect 10536 15744 10552 15808
rect 10616 15744 10632 15808
rect 10696 15744 10724 15808
rect 9484 14720 10724 15744
rect 9484 14656 9512 14720
rect 9576 14656 9592 14720
rect 9656 14656 9672 14720
rect 9736 14656 9752 14720
rect 9816 14656 9832 14720
rect 9896 14656 9912 14720
rect 9976 14656 9992 14720
rect 10056 14656 10072 14720
rect 10136 14656 10152 14720
rect 10216 14656 10232 14720
rect 10296 14656 10312 14720
rect 10376 14656 10392 14720
rect 10456 14656 10472 14720
rect 10536 14656 10552 14720
rect 10616 14656 10632 14720
rect 10696 14656 10724 14720
rect 9484 13632 10724 14656
rect 9484 13568 9512 13632
rect 9576 13568 9592 13632
rect 9656 13568 9672 13632
rect 9736 13568 9752 13632
rect 9816 13568 9832 13632
rect 9896 13568 9912 13632
rect 9976 13568 9992 13632
rect 10056 13568 10072 13632
rect 10136 13568 10152 13632
rect 10216 13568 10232 13632
rect 10296 13568 10312 13632
rect 10376 13568 10392 13632
rect 10456 13568 10472 13632
rect 10536 13568 10552 13632
rect 10616 13568 10632 13632
rect 10696 13568 10724 13632
rect 9484 12544 10724 13568
rect 9484 12480 9512 12544
rect 9576 12480 9592 12544
rect 9656 12480 9672 12544
rect 9736 12480 9752 12544
rect 9816 12480 9832 12544
rect 9896 12480 9912 12544
rect 9976 12480 9992 12544
rect 10056 12480 10072 12544
rect 10136 12480 10152 12544
rect 10216 12480 10232 12544
rect 10296 12480 10312 12544
rect 10376 12480 10392 12544
rect 10456 12480 10472 12544
rect 10536 12480 10552 12544
rect 10616 12480 10632 12544
rect 10696 12480 10724 12544
rect 9484 11456 10724 12480
rect 9484 11392 9512 11456
rect 9576 11392 9592 11456
rect 9656 11392 9672 11456
rect 9736 11392 9752 11456
rect 9816 11392 9832 11456
rect 9896 11392 9912 11456
rect 9976 11392 9992 11456
rect 10056 11392 10072 11456
rect 10136 11392 10152 11456
rect 10216 11392 10232 11456
rect 10296 11392 10312 11456
rect 10376 11392 10392 11456
rect 10456 11392 10472 11456
rect 10536 11392 10552 11456
rect 10616 11392 10632 11456
rect 10696 11392 10724 11456
rect 9484 10368 10724 11392
rect 9484 10304 9512 10368
rect 9576 10304 9592 10368
rect 9656 10304 9672 10368
rect 9736 10304 9752 10368
rect 9816 10304 9832 10368
rect 9896 10304 9912 10368
rect 9976 10304 9992 10368
rect 10056 10304 10072 10368
rect 10136 10304 10152 10368
rect 10216 10304 10232 10368
rect 10296 10304 10312 10368
rect 10376 10304 10392 10368
rect 10456 10304 10472 10368
rect 10536 10304 10552 10368
rect 10616 10304 10632 10368
rect 10696 10304 10724 10368
rect 9484 9280 10724 10304
rect 9484 9216 9512 9280
rect 9576 9216 9592 9280
rect 9656 9216 9672 9280
rect 9736 9216 9752 9280
rect 9816 9216 9832 9280
rect 9896 9216 9912 9280
rect 9976 9216 9992 9280
rect 10056 9216 10072 9280
rect 10136 9216 10152 9280
rect 10216 9216 10232 9280
rect 10296 9216 10312 9280
rect 10376 9216 10392 9280
rect 10456 9216 10472 9280
rect 10536 9216 10552 9280
rect 10616 9216 10632 9280
rect 10696 9216 10724 9280
rect 9484 8192 10724 9216
rect 9484 8128 9512 8192
rect 9576 8128 9592 8192
rect 9656 8128 9672 8192
rect 9736 8128 9752 8192
rect 9816 8128 9832 8192
rect 9896 8128 9912 8192
rect 9976 8128 9992 8192
rect 10056 8128 10072 8192
rect 10136 8128 10152 8192
rect 10216 8128 10232 8192
rect 10296 8128 10312 8192
rect 10376 8128 10392 8192
rect 10456 8128 10472 8192
rect 10536 8128 10552 8192
rect 10616 8128 10632 8192
rect 10696 8128 10724 8192
rect 9484 7104 10724 8128
rect 9484 7040 9512 7104
rect 9576 7040 9592 7104
rect 9656 7040 9672 7104
rect 9736 7040 9752 7104
rect 9816 7040 9832 7104
rect 9896 7040 9912 7104
rect 9976 7040 9992 7104
rect 10056 7040 10072 7104
rect 10136 7040 10152 7104
rect 10216 7040 10232 7104
rect 10296 7040 10312 7104
rect 10376 7040 10392 7104
rect 10456 7040 10472 7104
rect 10536 7040 10552 7104
rect 10616 7040 10632 7104
rect 10696 7040 10724 7104
rect 9484 6016 10724 7040
rect 9484 5952 9512 6016
rect 9576 5952 9592 6016
rect 9656 5952 9672 6016
rect 9736 5952 9752 6016
rect 9816 5952 9832 6016
rect 9896 5952 9912 6016
rect 9976 5952 9992 6016
rect 10056 5952 10072 6016
rect 10136 5952 10152 6016
rect 10216 5952 10232 6016
rect 10296 5952 10312 6016
rect 10376 5952 10392 6016
rect 10456 5952 10472 6016
rect 10536 5952 10552 6016
rect 10616 5952 10632 6016
rect 10696 5952 10724 6016
rect 9484 4928 10724 5952
rect 9484 4864 9512 4928
rect 9576 4864 9592 4928
rect 9656 4864 9672 4928
rect 9736 4864 9752 4928
rect 9816 4864 9832 4928
rect 9896 4864 9912 4928
rect 9976 4864 9992 4928
rect 10056 4864 10072 4928
rect 10136 4864 10152 4928
rect 10216 4864 10232 4928
rect 10296 4864 10312 4928
rect 10376 4864 10392 4928
rect 10456 4864 10472 4928
rect 10536 4864 10552 4928
rect 10616 4864 10632 4928
rect 10696 4864 10724 4928
rect 9484 3840 10724 4864
rect 9484 3776 9512 3840
rect 9576 3776 9592 3840
rect 9656 3776 9672 3840
rect 9736 3776 9752 3840
rect 9816 3776 9832 3840
rect 9896 3776 9912 3840
rect 9976 3776 9992 3840
rect 10056 3776 10072 3840
rect 10136 3776 10152 3840
rect 10216 3776 10232 3840
rect 10296 3776 10312 3840
rect 10376 3776 10392 3840
rect 10456 3776 10472 3840
rect 10536 3776 10552 3840
rect 10616 3776 10632 3840
rect 10696 3776 10724 3840
rect 9484 2752 10724 3776
rect 9484 2688 9512 2752
rect 9576 2688 9592 2752
rect 9656 2688 9672 2752
rect 9736 2688 9752 2752
rect 9816 2688 9832 2752
rect 9896 2688 9912 2752
rect 9976 2688 9992 2752
rect 10056 2688 10072 2752
rect 10136 2688 10152 2752
rect 10216 2688 10232 2752
rect 10296 2688 10312 2752
rect 10376 2688 10392 2752
rect 10456 2688 10472 2752
rect 10536 2688 10552 2752
rect 10616 2688 10632 2752
rect 10696 2688 10724 2752
rect 9484 2128 10724 2688
rect 13484 17440 14724 17456
rect 13484 17376 13512 17440
rect 13576 17376 13592 17440
rect 13656 17376 13672 17440
rect 13736 17376 13752 17440
rect 13816 17376 13832 17440
rect 13896 17376 13912 17440
rect 13976 17376 13992 17440
rect 14056 17376 14072 17440
rect 14136 17376 14152 17440
rect 14216 17376 14232 17440
rect 14296 17376 14312 17440
rect 14376 17376 14392 17440
rect 14456 17376 14472 17440
rect 14536 17376 14552 17440
rect 14616 17376 14632 17440
rect 14696 17376 14724 17440
rect 13484 16352 14724 17376
rect 13484 16288 13512 16352
rect 13576 16288 13592 16352
rect 13656 16288 13672 16352
rect 13736 16288 13752 16352
rect 13816 16288 13832 16352
rect 13896 16288 13912 16352
rect 13976 16288 13992 16352
rect 14056 16288 14072 16352
rect 14136 16288 14152 16352
rect 14216 16288 14232 16352
rect 14296 16288 14312 16352
rect 14376 16288 14392 16352
rect 14456 16288 14472 16352
rect 14536 16288 14552 16352
rect 14616 16288 14632 16352
rect 14696 16288 14724 16352
rect 13484 15264 14724 16288
rect 13484 15200 13512 15264
rect 13576 15200 13592 15264
rect 13656 15200 13672 15264
rect 13736 15200 13752 15264
rect 13816 15200 13832 15264
rect 13896 15200 13912 15264
rect 13976 15200 13992 15264
rect 14056 15200 14072 15264
rect 14136 15200 14152 15264
rect 14216 15200 14232 15264
rect 14296 15200 14312 15264
rect 14376 15200 14392 15264
rect 14456 15200 14472 15264
rect 14536 15200 14552 15264
rect 14616 15200 14632 15264
rect 14696 15200 14724 15264
rect 13484 14176 14724 15200
rect 13484 14112 13512 14176
rect 13576 14112 13592 14176
rect 13656 14112 13672 14176
rect 13736 14112 13752 14176
rect 13816 14112 13832 14176
rect 13896 14112 13912 14176
rect 13976 14112 13992 14176
rect 14056 14112 14072 14176
rect 14136 14112 14152 14176
rect 14216 14112 14232 14176
rect 14296 14112 14312 14176
rect 14376 14112 14392 14176
rect 14456 14112 14472 14176
rect 14536 14112 14552 14176
rect 14616 14112 14632 14176
rect 14696 14112 14724 14176
rect 13484 13088 14724 14112
rect 13484 13024 13512 13088
rect 13576 13024 13592 13088
rect 13656 13024 13672 13088
rect 13736 13024 13752 13088
rect 13816 13024 13832 13088
rect 13896 13024 13912 13088
rect 13976 13024 13992 13088
rect 14056 13024 14072 13088
rect 14136 13024 14152 13088
rect 14216 13024 14232 13088
rect 14296 13024 14312 13088
rect 14376 13024 14392 13088
rect 14456 13024 14472 13088
rect 14536 13024 14552 13088
rect 14616 13024 14632 13088
rect 14696 13024 14724 13088
rect 13484 12000 14724 13024
rect 13484 11936 13512 12000
rect 13576 11936 13592 12000
rect 13656 11936 13672 12000
rect 13736 11936 13752 12000
rect 13816 11936 13832 12000
rect 13896 11936 13912 12000
rect 13976 11936 13992 12000
rect 14056 11936 14072 12000
rect 14136 11936 14152 12000
rect 14216 11936 14232 12000
rect 14296 11936 14312 12000
rect 14376 11936 14392 12000
rect 14456 11936 14472 12000
rect 14536 11936 14552 12000
rect 14616 11936 14632 12000
rect 14696 11936 14724 12000
rect 13484 10912 14724 11936
rect 13484 10848 13512 10912
rect 13576 10848 13592 10912
rect 13656 10848 13672 10912
rect 13736 10848 13752 10912
rect 13816 10848 13832 10912
rect 13896 10848 13912 10912
rect 13976 10848 13992 10912
rect 14056 10848 14072 10912
rect 14136 10848 14152 10912
rect 14216 10848 14232 10912
rect 14296 10848 14312 10912
rect 14376 10848 14392 10912
rect 14456 10848 14472 10912
rect 14536 10848 14552 10912
rect 14616 10848 14632 10912
rect 14696 10848 14724 10912
rect 13484 9824 14724 10848
rect 13484 9760 13512 9824
rect 13576 9760 13592 9824
rect 13656 9760 13672 9824
rect 13736 9760 13752 9824
rect 13816 9760 13832 9824
rect 13896 9760 13912 9824
rect 13976 9760 13992 9824
rect 14056 9760 14072 9824
rect 14136 9760 14152 9824
rect 14216 9760 14232 9824
rect 14296 9760 14312 9824
rect 14376 9760 14392 9824
rect 14456 9760 14472 9824
rect 14536 9760 14552 9824
rect 14616 9760 14632 9824
rect 14696 9760 14724 9824
rect 13484 8736 14724 9760
rect 13484 8672 13512 8736
rect 13576 8672 13592 8736
rect 13656 8672 13672 8736
rect 13736 8672 13752 8736
rect 13816 8672 13832 8736
rect 13896 8672 13912 8736
rect 13976 8672 13992 8736
rect 14056 8672 14072 8736
rect 14136 8672 14152 8736
rect 14216 8672 14232 8736
rect 14296 8672 14312 8736
rect 14376 8672 14392 8736
rect 14456 8672 14472 8736
rect 14536 8672 14552 8736
rect 14616 8672 14632 8736
rect 14696 8672 14724 8736
rect 13484 7648 14724 8672
rect 13484 7584 13512 7648
rect 13576 7584 13592 7648
rect 13656 7584 13672 7648
rect 13736 7584 13752 7648
rect 13816 7584 13832 7648
rect 13896 7584 13912 7648
rect 13976 7584 13992 7648
rect 14056 7584 14072 7648
rect 14136 7584 14152 7648
rect 14216 7584 14232 7648
rect 14296 7584 14312 7648
rect 14376 7584 14392 7648
rect 14456 7584 14472 7648
rect 14536 7584 14552 7648
rect 14616 7584 14632 7648
rect 14696 7584 14724 7648
rect 13484 6560 14724 7584
rect 13484 6496 13512 6560
rect 13576 6496 13592 6560
rect 13656 6496 13672 6560
rect 13736 6496 13752 6560
rect 13816 6496 13832 6560
rect 13896 6496 13912 6560
rect 13976 6496 13992 6560
rect 14056 6496 14072 6560
rect 14136 6496 14152 6560
rect 14216 6496 14232 6560
rect 14296 6496 14312 6560
rect 14376 6496 14392 6560
rect 14456 6496 14472 6560
rect 14536 6496 14552 6560
rect 14616 6496 14632 6560
rect 14696 6496 14724 6560
rect 13484 5472 14724 6496
rect 13484 5408 13512 5472
rect 13576 5408 13592 5472
rect 13656 5408 13672 5472
rect 13736 5408 13752 5472
rect 13816 5408 13832 5472
rect 13896 5408 13912 5472
rect 13976 5408 13992 5472
rect 14056 5408 14072 5472
rect 14136 5408 14152 5472
rect 14216 5408 14232 5472
rect 14296 5408 14312 5472
rect 14376 5408 14392 5472
rect 14456 5408 14472 5472
rect 14536 5408 14552 5472
rect 14616 5408 14632 5472
rect 14696 5408 14724 5472
rect 13484 4384 14724 5408
rect 13484 4320 13512 4384
rect 13576 4320 13592 4384
rect 13656 4320 13672 4384
rect 13736 4320 13752 4384
rect 13816 4320 13832 4384
rect 13896 4320 13912 4384
rect 13976 4320 13992 4384
rect 14056 4320 14072 4384
rect 14136 4320 14152 4384
rect 14216 4320 14232 4384
rect 14296 4320 14312 4384
rect 14376 4320 14392 4384
rect 14456 4320 14472 4384
rect 14536 4320 14552 4384
rect 14616 4320 14632 4384
rect 14696 4320 14724 4384
rect 13484 3296 14724 4320
rect 13484 3232 13512 3296
rect 13576 3232 13592 3296
rect 13656 3232 13672 3296
rect 13736 3232 13752 3296
rect 13816 3232 13832 3296
rect 13896 3232 13912 3296
rect 13976 3232 13992 3296
rect 14056 3232 14072 3296
rect 14136 3232 14152 3296
rect 14216 3232 14232 3296
rect 14296 3232 14312 3296
rect 14376 3232 14392 3296
rect 14456 3232 14472 3296
rect 14536 3232 14552 3296
rect 14616 3232 14632 3296
rect 14696 3232 14724 3296
rect 13484 2208 14724 3232
rect 13484 2144 13512 2208
rect 13576 2144 13592 2208
rect 13656 2144 13672 2208
rect 13736 2144 13752 2208
rect 13816 2144 13832 2208
rect 13896 2144 13912 2208
rect 13976 2144 13992 2208
rect 14056 2144 14072 2208
rect 14136 2144 14152 2208
rect 14216 2144 14232 2208
rect 14296 2144 14312 2208
rect 14376 2144 14392 2208
rect 14456 2144 14472 2208
rect 14536 2144 14552 2208
rect 14616 2144 14632 2208
rect 14696 2144 14724 2208
rect 13484 2128 14724 2144
rect 17484 16896 18724 17456
rect 17484 16832 17512 16896
rect 17576 16832 17592 16896
rect 17656 16832 17672 16896
rect 17736 16832 17752 16896
rect 17816 16832 17832 16896
rect 17896 16832 17912 16896
rect 17976 16832 17992 16896
rect 18056 16832 18072 16896
rect 18136 16832 18152 16896
rect 18216 16832 18232 16896
rect 18296 16832 18312 16896
rect 18376 16832 18392 16896
rect 18456 16832 18472 16896
rect 18536 16832 18552 16896
rect 18616 16832 18632 16896
rect 18696 16832 18724 16896
rect 17484 15808 18724 16832
rect 17484 15744 17512 15808
rect 17576 15744 17592 15808
rect 17656 15744 17672 15808
rect 17736 15744 17752 15808
rect 17816 15744 17832 15808
rect 17896 15744 17912 15808
rect 17976 15744 17992 15808
rect 18056 15744 18072 15808
rect 18136 15744 18152 15808
rect 18216 15744 18232 15808
rect 18296 15744 18312 15808
rect 18376 15744 18392 15808
rect 18456 15744 18472 15808
rect 18536 15744 18552 15808
rect 18616 15744 18632 15808
rect 18696 15744 18724 15808
rect 17484 14720 18724 15744
rect 17484 14656 17512 14720
rect 17576 14656 17592 14720
rect 17656 14656 17672 14720
rect 17736 14656 17752 14720
rect 17816 14656 17832 14720
rect 17896 14656 17912 14720
rect 17976 14656 17992 14720
rect 18056 14656 18072 14720
rect 18136 14656 18152 14720
rect 18216 14656 18232 14720
rect 18296 14656 18312 14720
rect 18376 14656 18392 14720
rect 18456 14656 18472 14720
rect 18536 14656 18552 14720
rect 18616 14656 18632 14720
rect 18696 14656 18724 14720
rect 17484 13632 18724 14656
rect 17484 13568 17512 13632
rect 17576 13568 17592 13632
rect 17656 13568 17672 13632
rect 17736 13568 17752 13632
rect 17816 13568 17832 13632
rect 17896 13568 17912 13632
rect 17976 13568 17992 13632
rect 18056 13568 18072 13632
rect 18136 13568 18152 13632
rect 18216 13568 18232 13632
rect 18296 13568 18312 13632
rect 18376 13568 18392 13632
rect 18456 13568 18472 13632
rect 18536 13568 18552 13632
rect 18616 13568 18632 13632
rect 18696 13568 18724 13632
rect 17484 12544 18724 13568
rect 17484 12480 17512 12544
rect 17576 12480 17592 12544
rect 17656 12480 17672 12544
rect 17736 12480 17752 12544
rect 17816 12480 17832 12544
rect 17896 12480 17912 12544
rect 17976 12480 17992 12544
rect 18056 12480 18072 12544
rect 18136 12480 18152 12544
rect 18216 12480 18232 12544
rect 18296 12480 18312 12544
rect 18376 12480 18392 12544
rect 18456 12480 18472 12544
rect 18536 12480 18552 12544
rect 18616 12480 18632 12544
rect 18696 12480 18724 12544
rect 17484 11456 18724 12480
rect 18827 11660 18893 11661
rect 18827 11596 18828 11660
rect 18892 11596 18893 11660
rect 18827 11595 18893 11596
rect 17484 11392 17512 11456
rect 17576 11392 17592 11456
rect 17656 11392 17672 11456
rect 17736 11392 17752 11456
rect 17816 11392 17832 11456
rect 17896 11392 17912 11456
rect 17976 11392 17992 11456
rect 18056 11392 18072 11456
rect 18136 11392 18152 11456
rect 18216 11392 18232 11456
rect 18296 11392 18312 11456
rect 18376 11392 18392 11456
rect 18456 11392 18472 11456
rect 18536 11392 18552 11456
rect 18616 11392 18632 11456
rect 18696 11392 18724 11456
rect 17484 10368 18724 11392
rect 17484 10304 17512 10368
rect 17576 10304 17592 10368
rect 17656 10304 17672 10368
rect 17736 10304 17752 10368
rect 17816 10304 17832 10368
rect 17896 10304 17912 10368
rect 17976 10304 17992 10368
rect 18056 10304 18072 10368
rect 18136 10304 18152 10368
rect 18216 10304 18232 10368
rect 18296 10304 18312 10368
rect 18376 10304 18392 10368
rect 18456 10304 18472 10368
rect 18536 10304 18552 10368
rect 18616 10304 18632 10368
rect 18696 10304 18724 10368
rect 17484 9280 18724 10304
rect 17484 9216 17512 9280
rect 17576 9216 17592 9280
rect 17656 9216 17672 9280
rect 17736 9216 17752 9280
rect 17816 9216 17832 9280
rect 17896 9216 17912 9280
rect 17976 9216 17992 9280
rect 18056 9216 18072 9280
rect 18136 9216 18152 9280
rect 18216 9216 18232 9280
rect 18296 9216 18312 9280
rect 18376 9216 18392 9280
rect 18456 9216 18472 9280
rect 18536 9216 18552 9280
rect 18616 9216 18632 9280
rect 18696 9216 18724 9280
rect 17484 8192 18724 9216
rect 17484 8128 17512 8192
rect 17576 8128 17592 8192
rect 17656 8128 17672 8192
rect 17736 8128 17752 8192
rect 17816 8128 17832 8192
rect 17896 8128 17912 8192
rect 17976 8128 17992 8192
rect 18056 8128 18072 8192
rect 18136 8128 18152 8192
rect 18216 8128 18232 8192
rect 18296 8128 18312 8192
rect 18376 8128 18392 8192
rect 18456 8128 18472 8192
rect 18536 8128 18552 8192
rect 18616 8128 18632 8192
rect 18696 8128 18724 8192
rect 17484 7104 18724 8128
rect 17484 7040 17512 7104
rect 17576 7040 17592 7104
rect 17656 7040 17672 7104
rect 17736 7040 17752 7104
rect 17816 7040 17832 7104
rect 17896 7040 17912 7104
rect 17976 7040 17992 7104
rect 18056 7040 18072 7104
rect 18136 7040 18152 7104
rect 18216 7040 18232 7104
rect 18296 7040 18312 7104
rect 18376 7040 18392 7104
rect 18456 7040 18472 7104
rect 18536 7040 18552 7104
rect 18616 7040 18632 7104
rect 18696 7040 18724 7104
rect 17484 6016 18724 7040
rect 17484 5952 17512 6016
rect 17576 5952 17592 6016
rect 17656 5952 17672 6016
rect 17736 5952 17752 6016
rect 17816 5952 17832 6016
rect 17896 5952 17912 6016
rect 17976 5952 17992 6016
rect 18056 5952 18072 6016
rect 18136 5952 18152 6016
rect 18216 5952 18232 6016
rect 18296 5952 18312 6016
rect 18376 5952 18392 6016
rect 18456 5952 18472 6016
rect 18536 5952 18552 6016
rect 18616 5952 18632 6016
rect 18696 5952 18724 6016
rect 17484 4928 18724 5952
rect 18830 5133 18890 11595
rect 19011 10708 19077 10709
rect 19011 10644 19012 10708
rect 19076 10644 19077 10708
rect 19011 10643 19077 10644
rect 18827 5132 18893 5133
rect 18827 5068 18828 5132
rect 18892 5068 18893 5132
rect 18827 5067 18893 5068
rect 17484 4864 17512 4928
rect 17576 4864 17592 4928
rect 17656 4864 17672 4928
rect 17736 4864 17752 4928
rect 17816 4864 17832 4928
rect 17896 4864 17912 4928
rect 17976 4864 17992 4928
rect 18056 4864 18072 4928
rect 18136 4864 18152 4928
rect 18216 4864 18232 4928
rect 18296 4864 18312 4928
rect 18376 4864 18392 4928
rect 18456 4864 18472 4928
rect 18536 4864 18552 4928
rect 18616 4864 18632 4928
rect 18696 4864 18724 4928
rect 17484 3840 18724 4864
rect 19014 4181 19074 10643
rect 19195 9484 19261 9485
rect 19195 9420 19196 9484
rect 19260 9420 19261 9484
rect 19195 9419 19261 9420
rect 19198 4589 19258 9419
rect 19195 4588 19261 4589
rect 19195 4524 19196 4588
rect 19260 4524 19261 4588
rect 19195 4523 19261 4524
rect 19011 4180 19077 4181
rect 19011 4116 19012 4180
rect 19076 4116 19077 4180
rect 19011 4115 19077 4116
rect 17484 3776 17512 3840
rect 17576 3776 17592 3840
rect 17656 3776 17672 3840
rect 17736 3776 17752 3840
rect 17816 3776 17832 3840
rect 17896 3776 17912 3840
rect 17976 3776 17992 3840
rect 18056 3776 18072 3840
rect 18136 3776 18152 3840
rect 18216 3776 18232 3840
rect 18296 3776 18312 3840
rect 18376 3776 18392 3840
rect 18456 3776 18472 3840
rect 18536 3776 18552 3840
rect 18616 3776 18632 3840
rect 18696 3776 18724 3840
rect 17484 2752 18724 3776
rect 17484 2688 17512 2752
rect 17576 2688 17592 2752
rect 17656 2688 17672 2752
rect 17736 2688 17752 2752
rect 17816 2688 17832 2752
rect 17896 2688 17912 2752
rect 17976 2688 17992 2752
rect 18056 2688 18072 2752
rect 18136 2688 18152 2752
rect 18216 2688 18232 2752
rect 18296 2688 18312 2752
rect 18376 2688 18392 2752
rect 18456 2688 18472 2752
rect 18536 2688 18552 2752
rect 18616 2688 18632 2752
rect 18696 2688 18724 2752
rect 17484 2128 18724 2688
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1676037725
transform 1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1676037725
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1676037725
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1676037725
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1676037725
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123
timestamp 1676037725
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_178
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1676037725
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_12
timestamp 1676037725
transform 1 0 2208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1676037725
transform 1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1676037725
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1676037725
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_72
timestamp 1676037725
transform 1 0 7728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_83
timestamp 1676037725
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_128
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1676037725
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1676037725
transform 1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1676037725
transform 1 0 2208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_16
timestamp 1676037725
transform 1 0 2576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1676037725
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_49
timestamp 1676037725
transform 1 0 5612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1676037725
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_96
timestamp 1676037725
transform 1 0 9936 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_102
timestamp 1676037725
transform 1 0 10488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_113
timestamp 1676037725
transform 1 0 11500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_150
timestamp 1676037725
transform 1 0 14904 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_154
timestamp 1676037725
transform 1 0 15272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_176
timestamp 1676037725
transform 1 0 17296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp 1676037725
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1676037725
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_16
timestamp 1676037725
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 1676037725
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_35
timestamp 1676037725
transform 1 0 4324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_66
timestamp 1676037725
transform 1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_70
timestamp 1676037725
transform 1 0 7544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_78
timestamp 1676037725
transform 1 0 8280 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_84
timestamp 1676037725
transform 1 0 8832 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1676037725
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_123
timestamp 1676037725
transform 1 0 12420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_144
timestamp 1676037725
transform 1 0 14352 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp 1676037725
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_186
timestamp 1676037725
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_12
timestamp 1676037725
transform 1 0 2208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_16
timestamp 1676037725
transform 1 0 2576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1676037725
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_49
timestamp 1676037725
transform 1 0 5612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1676037725
transform 1 0 6716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1676037725
transform 1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1676037725
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1676037725
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1676037725
transform 1 0 11684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1676037725
transform 1 0 12880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_151
timestamp 1676037725
transform 1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_176
timestamp 1676037725
transform 1 0 17296 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_187
timestamp 1676037725
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1676037725
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1676037725
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 1676037725
transform 1 0 3956 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_35
timestamp 1676037725
transform 1 0 4324 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1676037725
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp 1676037725
transform 1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_70
timestamp 1676037725
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_78
timestamp 1676037725
transform 1 0 8280 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_84
timestamp 1676037725
transform 1 0 8832 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1676037725
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_136
timestamp 1676037725
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1676037725
transform 1 0 17480 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1676037725
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_12
timestamp 1676037725
transform 1 0 2208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_16
timestamp 1676037725
transform 1 0 2576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1676037725
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_49
timestamp 1676037725
transform 1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_61
timestamp 1676037725
transform 1 0 6716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_68
timestamp 1676037725
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1676037725
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_90
timestamp 1676037725
transform 1 0 9384 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_98
timestamp 1676037725
transform 1 0 10120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_120
timestamp 1676037725
transform 1 0 12144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_150
timestamp 1676037725
transform 1 0 14904 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_175
timestamp 1676037725
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1676037725
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_16
timestamp 1676037725
transform 1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp 1676037725
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_35
timestamp 1676037725
transform 1 0 4324 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1676037725
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp 1676037725
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1676037725
transform 1 0 7544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_78
timestamp 1676037725
transform 1 0 8280 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_84
timestamp 1676037725
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_103
timestamp 1676037725
transform 1 0 10580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1676037725
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_151
timestamp 1676037725
transform 1 0 14996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1676037725
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1676037725
transform 1 0 18400 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1676037725
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_16
timestamp 1676037725
transform 1 0 2576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1676037725
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_49
timestamp 1676037725
transform 1 0 5612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1676037725
transform 1 0 6716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_68
timestamp 1676037725
transform 1 0 7360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1676037725
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_90
timestamp 1676037725
transform 1 0 9384 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_115
timestamp 1676037725
transform 1 0 11684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1676037725
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1676037725
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_164
timestamp 1676037725
transform 1 0 16192 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_172
timestamp 1676037725
transform 1 0 16928 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1676037725
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1676037725
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_31
timestamp 1676037725
transform 1 0 3956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_35
timestamp 1676037725
transform 1 0 4324 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_43
timestamp 1676037725
transform 1 0 5060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1676037725
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_66
timestamp 1676037725
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_70
timestamp 1676037725
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_78
timestamp 1676037725
transform 1 0 8280 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_84
timestamp 1676037725
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1676037725
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1676037725
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_141
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1676037725
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1676037725
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_16
timestamp 1676037725
transform 1 0 2576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1676037725
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_49
timestamp 1676037725
transform 1 0 5612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_61
timestamp 1676037725
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1676037725
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1676037725
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_90
timestamp 1676037725
transform 1 0 9384 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_99
timestamp 1676037725
transform 1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1676037725
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_150
timestamp 1676037725
transform 1 0 14904 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_156
timestamp 1676037725
transform 1 0 15456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_187
timestamp 1676037725
transform 1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_9
timestamp 1676037725
transform 1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_16
timestamp 1676037725
transform 1 0 2576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_31
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1676037725
transform 1 0 4324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1676037725
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1676037725
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_70
timestamp 1676037725
transform 1 0 7544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_78
timestamp 1676037725
transform 1 0 8280 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_84
timestamp 1676037725
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1676037725
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_123
timestamp 1676037725
transform 1 0 12420 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1676037725
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1676037725
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1676037725
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_187
timestamp 1676037725
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_12
timestamp 1676037725
transform 1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_16
timestamp 1676037725
transform 1 0 2576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1676037725
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_49
timestamp 1676037725
transform 1 0 5612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_61
timestamp 1676037725
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_68
timestamp 1676037725
transform 1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1676037725
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_90
timestamp 1676037725
transform 1 0 9384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1676037725
transform 1 0 10488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1676037725
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1676037725
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_164
timestamp 1676037725
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1676037725
transform 1 0 17020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_187
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_9
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_16
timestamp 1676037725
transform 1 0 2576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_31
timestamp 1676037725
transform 1 0 3956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1676037725
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_66
timestamp 1676037725
transform 1 0 7176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_70
timestamp 1676037725
transform 1 0 7544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_78
timestamp 1676037725
transform 1 0 8280 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_84
timestamp 1676037725
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1676037725
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_124
timestamp 1676037725
transform 1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1676037725
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1676037725
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1676037725
transform 1 0 17480 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_12
timestamp 1676037725
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_16
timestamp 1676037725
transform 1 0 2576 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1676037725
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_49
timestamp 1676037725
transform 1 0 5612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1676037725
transform 1 0 6716 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_68
timestamp 1676037725
transform 1 0 7360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1676037725
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_90
timestamp 1676037725
transform 1 0 9384 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_99
timestamp 1676037725
transform 1 0 10212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_116
timestamp 1676037725
transform 1 0 11776 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_124
timestamp 1676037725
transform 1 0 12512 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_148
timestamp 1676037725
transform 1 0 14720 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1676037725
transform 1 0 18400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_10
timestamp 1676037725
transform 1 0 2024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_38
timestamp 1676037725
transform 1 0 4600 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_44
timestamp 1676037725
transform 1 0 5152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_86
timestamp 1676037725
transform 1 0 9016 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_94
timestamp 1676037725
transform 1 0 9752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1676037725
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_127
timestamp 1676037725
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_144
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1676037725
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1676037725
transform 1 0 17388 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_186
timestamp 1676037725
transform 1 0 18216 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1676037725
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_40
timestamp 1676037725
transform 1 0 4784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_48
timestamp 1676037725
transform 1 0 5520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_62
timestamp 1676037725
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1676037725
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_108
timestamp 1676037725
transform 1 0 11040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_119
timestamp 1676037725
transform 1 0 12052 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_158
timestamp 1676037725
transform 1 0 15640 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1676037725
transform 1 0 16836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_180
timestamp 1676037725
transform 1 0 17664 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1676037725
transform 1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_20
timestamp 1676037725
transform 1 0 2944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_28
timestamp 1676037725
transform 1 0 3680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1676037725
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_67
timestamp 1676037725
transform 1 0 7268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_71
timestamp 1676037725
transform 1 0 7636 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_95
timestamp 1676037725
transform 1 0 9844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1676037725
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_129
timestamp 1676037725
transform 1 0 12972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1676037725
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1676037725
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1676037725
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_180
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_186
timestamp 1676037725
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1676037725
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_57
timestamp 1676037725
transform 1 0 6348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_66
timestamp 1676037725
transform 1 0 7176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_96
timestamp 1676037725
transform 1 0 9936 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1676037725
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_118
timestamp 1676037725
transform 1 0 11960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1676037725
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1676037725
transform 1 0 14720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1676037725
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_161
timestamp 1676037725
transform 1 0 15916 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1676037725
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_185
timestamp 1676037725
transform 1 0 18124 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_16
timestamp 1676037725
transform 1 0 2576 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_24
timestamp 1676037725
transform 1 0 3312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_36
timestamp 1676037725
transform 1 0 4416 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_42
timestamp 1676037725
transform 1 0 4968 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1676037725
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_67
timestamp 1676037725
transform 1 0 7268 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_78
timestamp 1676037725
transform 1 0 8280 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_84
timestamp 1676037725
transform 1 0 8832 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1676037725
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1676037725
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_128
timestamp 1676037725
transform 1 0 12880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_139
timestamp 1676037725
transform 1 0 13892 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_148
timestamp 1676037725
transform 1 0 14720 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_157
timestamp 1676037725
transform 1 0 15548 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_176 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17296 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp 1676037725
transform 1 0 18400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_10
timestamp 1676037725
transform 1 0 2024 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1676037725
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_39
timestamp 1676037725
transform 1 0 4692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_48
timestamp 1676037725
transform 1 0 5520 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1676037725
transform 1 0 6532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1676037725
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1676037725
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1676037725
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_113
timestamp 1676037725
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_130
timestamp 1676037725
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_148
timestamp 1676037725
transform 1 0 14720 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp 1676037725
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_164
timestamp 1676037725
transform 1 0 16192 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_170
timestamp 1676037725
transform 1 0 16744 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_182
timestamp 1676037725
transform 1 0 17848 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 1676037725
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_26
timestamp 1676037725
transform 1 0 3496 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1676037725
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_66
timestamp 1676037725
transform 1 0 7176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_76
timestamp 1676037725
transform 1 0 8096 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1676037725
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_94
timestamp 1676037725
transform 1 0 9752 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_103
timestamp 1676037725
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_120
timestamp 1676037725
transform 1 0 12144 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_129
timestamp 1676037725
transform 1 0 12972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_133
timestamp 1676037725
transform 1 0 13340 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_139
timestamp 1676037725
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_148
timestamp 1676037725
transform 1 0 14720 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1676037725
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1676037725
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1676037725
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1676037725
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_52
timestamp 1676037725
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_63
timestamp 1676037725
transform 1 0 6900 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1676037725
transform 1 0 7636 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1676037725
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_92
timestamp 1676037725
transform 1 0 9568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1676037725
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_103
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_129
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_14
timestamp 1676037725
transform 1 0 2392 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_22
timestamp 1676037725
transform 1 0 3128 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_32
timestamp 1676037725
transform 1 0 4048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_43
timestamp 1676037725
transform 1 0 5060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1676037725
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_65
timestamp 1676037725
transform 1 0 7084 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_74
timestamp 1676037725
transform 1 0 7912 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_83
timestamp 1676037725
transform 1 0 8740 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_92
timestamp 1676037725
transform 1 0 9568 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1676037725
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_13
timestamp 1676037725
transform 1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1676037725
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_38
timestamp 1676037725
transform 1 0 4600 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_50
timestamp 1676037725
transform 1 0 5704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_59
timestamp 1676037725
transform 1 0 6532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_68
timestamp 1676037725
transform 1 0 7360 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_92
timestamp 1676037725
transform 1 0 9568 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_104
timestamp 1676037725
transform 1 0 10672 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_116
timestamp 1676037725
transform 1 0 11776 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_128
timestamp 1676037725
transform 1 0 12880 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_18
timestamp 1676037725
transform 1 0 2760 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_24
timestamp 1676037725
transform 1 0 3312 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1676037725
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_42
timestamp 1676037725
transform 1 0 4968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_46
timestamp 1676037725
transform 1 0 5336 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1676037725
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_64
timestamp 1676037725
transform 1 0 6992 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_73
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_85
timestamp 1676037725
transform 1 0 8924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_97
timestamp 1676037725
transform 1 0 10028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1676037725
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_189
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_10
timestamp 1676037725
transform 1 0 2024 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_36
timestamp 1676037725
transform 1 0 4416 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_44
timestamp 1676037725
transform 1 0 5152 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_50
timestamp 1676037725
transform 1 0 5704 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_71
timestamp 1676037725
transform 1 0 7636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_17
timestamp 1676037725
transform 1 0 2668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1676037725
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1676037725
transform 1 0 3772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_36
timestamp 1676037725
transform 1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1676037725
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1676037725
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_153
timestamp 1676037725
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1676037725
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1676037725
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10212 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1676037725
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1676037725
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1676037725
transform -1 0 11224 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12052 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _181_
timestamp 1676037725
transform 1 0 14904 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _182_
timestamp 1676037725
transform 1 0 12052 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _183_
timestamp 1676037725
transform 1 0 13248 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 1676037725
transform 1 0 12512 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1676037725
transform 1 0 17296 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 1676037725
transform 1 0 17480 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18216 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13800 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14996 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _195_
timestamp 1676037725
transform 1 0 17664 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _196_
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _197_
timestamp 1676037725
transform 1 0 17020 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _198_
timestamp 1676037725
transform -1 0 18216 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15364 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _201_
timestamp 1676037725
transform 1 0 8464 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _202_
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _203_
timestamp 1676037725
transform -1 0 8740 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _204_
timestamp 1676037725
transform -1 0 13892 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _205_
timestamp 1676037725
transform -1 0 14352 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _206_
timestamp 1676037725
transform 1 0 14260 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _207_
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _208_
timestamp 1676037725
transform 1 0 17848 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _209_
timestamp 1676037725
transform 1 0 5244 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _210_
timestamp 1676037725
transform -1 0 12972 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _211_
timestamp 1676037725
transform 1 0 15088 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _212_
timestamp 1676037725
transform 1 0 7360 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _215_
timestamp 1676037725
transform 1 0 12788 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _216_
timestamp 1676037725
transform 1 0 17848 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _217_
timestamp 1676037725
transform -1 0 14720 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _218_
timestamp 1676037725
transform -1 0 11132 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _219_
timestamp 1676037725
transform -1 0 11224 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__o211ai_2  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _221_
timestamp 1676037725
transform 1 0 17848 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _222_
timestamp 1676037725
transform -1 0 14720 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _223_
timestamp 1676037725
transform -1 0 17480 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _224_
timestamp 1676037725
transform -1 0 9660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _225_
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_2  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9936 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _227_
timestamp 1676037725
transform -1 0 18308 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _228_
timestamp 1676037725
transform -1 0 9568 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_2  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8372 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _230_
timestamp 1676037725
transform -1 0 9568 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _231_
timestamp 1676037725
transform -1 0 6992 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _232_
timestamp 1676037725
transform -1 0 6532 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _234_
timestamp 1676037725
transform 1 0 6256 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _235_
timestamp 1676037725
transform -1 0 6072 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__o2bb2a_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9936 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_2  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7360 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8556 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _239_
timestamp 1676037725
transform -1 0 18308 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _240_
timestamp 1676037725
transform 1 0 8924 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _241_
timestamp 1676037725
transform -1 0 11132 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _242_
timestamp 1676037725
transform 1 0 9844 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_2  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10488 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _245_
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _246_
timestamp 1676037725
transform -1 0 12144 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _247_
timestamp 1676037725
transform 1 0 11408 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _249_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_2  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and4_2  _252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17572 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _253_
timestamp 1676037725
transform -1 0 13064 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _254_
timestamp 1676037725
transform -1 0 9568 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _255_
timestamp 1676037725
transform -1 0 10028 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _256_
timestamp 1676037725
transform -1 0 5520 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _257_
timestamp 1676037725
transform 1 0 9292 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _260_
timestamp 1676037725
transform -1 0 18216 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12144 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _262_
timestamp 1676037725
transform 1 0 9752 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _263_
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _264_
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _265_
timestamp 1676037725
transform -1 0 12236 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _266_
timestamp 1676037725
transform 1 0 12328 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _267_
timestamp 1676037725
transform -1 0 14168 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _268_
timestamp 1676037725
transform 1 0 10396 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _270_
timestamp 1676037725
transform 1 0 12052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11040 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _272_
timestamp 1676037725
transform 1 0 9568 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9844 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _274_
timestamp 1676037725
transform -1 0 8372 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _275_
timestamp 1676037725
transform 1 0 9752 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _276_
timestamp 1676037725
transform 1 0 10212 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _277_
timestamp 1676037725
transform 1 0 10580 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp 1676037725
transform -1 0 12512 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _279_
timestamp 1676037725
transform 1 0 12604 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _280_
timestamp 1676037725
transform 1 0 3404 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _281_
timestamp 1676037725
transform -1 0 4048 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _282_
timestamp 1676037725
transform -1 0 7176 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _283_
timestamp 1676037725
transform -1 0 5888 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _284_
timestamp 1676037725
transform -1 0 13524 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _285_
timestamp 1676037725
transform 1 0 5888 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _286_
timestamp 1676037725
transform -1 0 2024 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _287_
timestamp 1676037725
transform -1 0 13524 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _288_
timestamp 1676037725
transform 1 0 14904 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _289_
timestamp 1676037725
transform -1 0 3036 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _290_
timestamp 1676037725
transform -1 0 2760 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _291_
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _292_
timestamp 1676037725
transform -1 0 3312 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _293_
timestamp 1676037725
transform -1 0 4416 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _294_
timestamp 1676037725
transform -1 0 3496 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _295_
timestamp 1676037725
transform -1 0 2024 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _296_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _297_
timestamp 1676037725
transform -1 0 6532 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _298_
timestamp 1676037725
transform -1 0 8188 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _299_
timestamp 1676037725
transform 1 0 7544 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _300_
timestamp 1676037725
transform 1 0 2852 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _301_
timestamp 1676037725
transform -1 0 2300 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _302_
timestamp 1676037725
transform -1 0 8556 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_2  _303_
timestamp 1676037725
transform -1 0 6072 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_2  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _305_
timestamp 1676037725
transform -1 0 4416 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _306_
timestamp 1676037725
transform -1 0 4600 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _307_
timestamp 1676037725
transform -1 0 7360 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _308_
timestamp 1676037725
transform -1 0 7176 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _309_
timestamp 1676037725
transform -1 0 8280 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _310_
timestamp 1676037725
transform -1 0 4416 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _311_
timestamp 1676037725
transform 1 0 2392 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_2  _312_
timestamp 1676037725
transform 1 0 3956 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _313_
timestamp 1676037725
transform -1 0 2484 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _314_
timestamp 1676037725
transform -1 0 2392 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6900 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _316_
timestamp 1676037725
transform 1 0 5888 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or3_2  _317_
timestamp 1676037725
transform -1 0 5980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _318_
timestamp 1676037725
transform 1 0 5060 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_2  _319_
timestamp 1676037725
transform 1 0 5060 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _320_
timestamp 1676037725
transform 1 0 4232 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _321_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _322_
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _324_
timestamp 1676037725
transform 1 0 4416 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _325_
timestamp 1676037725
transform 1 0 5152 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _326_
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _327_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _329_
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_2  _331_
timestamp 1676037725
transform 1 0 2024 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _332_
timestamp 1676037725
transform -1 0 2392 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_2  _333_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _334_
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _335_
timestamp 1676037725
transform -1 0 2944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _336_
timestamp 1676037725
transform 1 0 1748 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _337_
timestamp 1676037725
transform -1 0 2668 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_2  _338_
timestamp 1676037725
transform 1 0 1656 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _339_
timestamp 1676037725
transform 1 0 2392 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _340_
timestamp 1676037725
transform -1 0 14536 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _341_
timestamp 1676037725
transform 1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_2  _342_
timestamp 1676037725
transform -1 0 6072 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _343_
timestamp 1676037725
transform 1 0 15548 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _344_
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _345_
timestamp 1676037725
transform -1 0 5060 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _346_
timestamp 1676037725
transform 1 0 5244 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _347_
timestamp 1676037725
transform 1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _348_
timestamp 1676037725
transform 1 0 5060 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_2  _349_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4600 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_2  _350_
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _351_
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _352_
timestamp 1676037725
transform -1 0 17020 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _353_
timestamp 1676037725
transform -1 0 14720 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _354_
timestamp 1676037725
transform -1 0 13708 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _355_
timestamp 1676037725
transform -1 0 15180 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _356_
timestamp 1676037725
transform -1 0 16284 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _357_
timestamp 1676037725
transform 1 0 17848 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _358_
timestamp 1676037725
transform -1 0 16008 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _359_
timestamp 1676037725
transform -1 0 17296 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _360_
timestamp 1676037725
transform -1 0 16744 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _361_
timestamp 1676037725
transform -1 0 17296 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _362_
timestamp 1676037725
transform -1 0 15548 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _363_
timestamp 1676037725
transform -1 0 14996 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _364_
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _365_
timestamp 1676037725
transform -1 0 17664 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _366_
timestamp 1676037725
transform -1 0 17296 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _367_
timestamp 1676037725
transform 1 0 4784 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _368_
timestamp 1676037725
transform -1 0 15824 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _369_
timestamp 1676037725
transform 1 0 16008 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _370_
timestamp 1676037725
transform -1 0 15640 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _371_
timestamp 1676037725
transform -1 0 13616 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _372_
timestamp 1676037725
transform 1 0 10120 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _373_
timestamp 1676037725
transform -1 0 16376 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _374_
timestamp 1676037725
transform -1 0 14996 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _375_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _376_
timestamp 1676037725
transform -1 0 12512 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _377_
timestamp 1676037725
transform -1 0 11684 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _378_
timestamp 1676037725
transform 1 0 7084 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _379_
timestamp 1676037725
transform 1 0 11592 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _380_
timestamp 1676037725
transform -1 0 14076 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _381_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _382_
timestamp 1676037725
transform 1 0 15364 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _383_
timestamp 1676037725
transform -1 0 16376 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _384_
timestamp 1676037725
transform 1 0 15364 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _385_
timestamp 1676037725
transform 1 0 13984 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _386_
timestamp 1676037725
transform -1 0 14168 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1676037725
transform 1 0 15456 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _389_
timestamp 1676037725
transform 1 0 14444 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _390_
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1676037725
transform 1 0 15272 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1676037725
transform 1 0 11684 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1676037725
transform 1 0 11868 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1676037725
transform -1 0 11684 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _396_
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _397_
timestamp 1676037725
transform -1 0 12144 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3312 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1676037725
transform -1 0 3588 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5612 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2208 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1676037725
transform -1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1676037725
transform -1 0 3312 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1676037725
transform -1 0 3588 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1676037725
transform -1 0 5612 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb1
timestamp 1676037725
transform -1 0 2208 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1676037725
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1676037725
transform -1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1676037725
transform -1 0 3312 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1676037725
transform -1 0 3588 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1676037725
transform -1 0 5612 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb1
timestamp 1676037725
transform -1 0 2208 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1676037725
transform 1 0 4048 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1676037725
transform -1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1676037725
transform -1 0 3312 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1676037725
transform -1 0 3588 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1676037725
transform -1 0 5612 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb1
timestamp 1676037725
transform -1 0 2208 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1676037725
transform 1 0 4048 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1676037725
transform -1 0 2576 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1676037725
transform -1 0 3312 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1676037725
transform -1 0 3588 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1676037725
transform -1 0 5612 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb1
timestamp 1676037725
transform -1 0 2208 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1676037725
transform 1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1676037725
transform -1 0 2576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1676037725
transform -1 0 3312 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1676037725
transform -1 0 3588 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1676037725
transform -1 0 5612 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1676037725
transform -1 0 2208 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1676037725
transform 1 0 4048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1676037725
transform -1 0 6716 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1676037725
transform 1 0 7636 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1676037725
transform 1 0 7728 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1676037725
transform 1 0 8924 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1676037725
transform 1 0 6532 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1676037725
transform -1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1676037725
transform -1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1676037725
transform 1 0 7636 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1676037725
transform 1 0 7728 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1676037725
transform 1 0 8924 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb1
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1676037725
transform -1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1676037725
transform -1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1676037725
transform 1 0 7636 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1676037725
transform 1 0 7728 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1676037725
transform 1 0 6532 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1676037725
transform -1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1676037725
transform -1 0 6716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1676037725
transform 1 0 7636 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1676037725
transform 1 0 7728 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1676037725
transform 1 0 8924 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1676037725
transform 1 0 6532 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1676037725
transform -1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1676037725
transform -1 0 6716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1676037725
transform 1 0 7636 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1676037725
transform 1 0 7728 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1676037725
transform 1 0 8924 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb1
timestamp 1676037725
transform 1 0 6532 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1676037725
transform -1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1676037725
transform -1 0 6716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1676037725
transform 1 0 7636 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1676037725
transform 1 0 7728 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1676037725
transform 1 0 8924 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[11\].id.delayenb1
timestamp 1676037725
transform 1 0 6532 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1676037725
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5796 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1676037725
transform 1 0 8280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1676037725
transform -1 0 5796 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1676037725
transform -1 0 3404 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1676037725
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1676037725
transform -1 0 3312 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1676037725
transform -1 0 2944 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1676037725
transform -1 0 5612 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.iss.delayenb1
timestamp 1676037725
transform -1 0 2208 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2024 0 1 2176
box -38 -48 498 592
<< labels >>
flabel metal4 s 5484 2128 6724 17456 0 FreeSans 7680 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 13484 2128 14724 17456 0 FreeSans 7680 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1484 2128 2724 17456 0 FreeSans 7680 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9484 2128 10724 17456 0 FreeSans 7680 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 17484 2128 18724 17456 0 FreeSans 7680 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 416 800 536 0 FreeSans 480 0 0 0 clockp[0]
port 2 nsew signal tristate
flabel metal3 s 0 144 800 264 0 FreeSans 480 0 0 0 clockp[1]
port 3 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 1232 800 1352 0 FreeSans 480 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 960 800 1080 0 FreeSans 480 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 enable
port 10 nsew signal input
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 ext_trim[0]
port 11 nsew signal input
flabel metal2 s 2318 19200 2374 20000 0 FreeSans 224 90 0 0 ext_trim[10]
port 12 nsew signal input
flabel metal2 s 2134 19200 2190 20000 0 FreeSans 224 90 0 0 ext_trim[11]
port 13 nsew signal input
flabel metal2 s 1950 19200 2006 20000 0 FreeSans 224 90 0 0 ext_trim[12]
port 14 nsew signal input
flabel metal2 s 1766 19200 1822 20000 0 FreeSans 224 90 0 0 ext_trim[13]
port 15 nsew signal input
flabel metal2 s 1582 19200 1638 20000 0 FreeSans 224 90 0 0 ext_trim[14]
port 16 nsew signal input
flabel metal2 s 1398 19200 1454 20000 0 FreeSans 224 90 0 0 ext_trim[15]
port 17 nsew signal input
flabel metal2 s 1214 19200 1270 20000 0 FreeSans 224 90 0 0 ext_trim[16]
port 18 nsew signal input
flabel metal2 s 1030 19200 1086 20000 0 FreeSans 224 90 0 0 ext_trim[17]
port 19 nsew signal input
flabel metal2 s 846 19200 902 20000 0 FreeSans 224 90 0 0 ext_trim[18]
port 20 nsew signal input
flabel metal2 s 662 19200 718 20000 0 FreeSans 224 90 0 0 ext_trim[19]
port 21 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 ext_trim[1]
port 22 nsew signal input
flabel metal3 s 19200 1504 20000 1624 0 FreeSans 480 0 0 0 ext_trim[20]
port 23 nsew signal input
flabel metal3 s 19200 1232 20000 1352 0 FreeSans 480 0 0 0 ext_trim[21]
port 24 nsew signal input
flabel metal3 s 19200 960 20000 1080 0 FreeSans 480 0 0 0 ext_trim[22]
port 25 nsew signal input
flabel metal3 s 19200 688 20000 808 0 FreeSans 480 0 0 0 ext_trim[23]
port 26 nsew signal input
flabel metal3 s 19200 416 20000 536 0 FreeSans 480 0 0 0 ext_trim[24]
port 27 nsew signal input
flabel metal3 s 19200 144 20000 264 0 FreeSans 480 0 0 0 ext_trim[25]
port 28 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 ext_trim[2]
port 29 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 ext_trim[3]
port 30 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 ext_trim[4]
port 31 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 ext_trim[5]
port 32 nsew signal input
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 ext_trim[6]
port 33 nsew signal input
flabel metal2 s 110 19200 166 20000 0 FreeSans 224 90 0 0 ext_trim[7]
port 34 nsew signal input
flabel metal2 s 294 19200 350 20000 0 FreeSans 224 90 0 0 ext_trim[8]
port 35 nsew signal input
flabel metal2 s 478 19200 534 20000 0 FreeSans 224 90 0 0 ext_trim[9]
port 36 nsew signal input
flabel metal2 s 294 0 350 800 0 FreeSans 224 90 0 0 osc
port 37 nsew signal input
flabel metal2 s 110 0 166 800 0 FreeSans 224 90 0 0 resetb
port 38 nsew signal input
rlabel metal1 9982 17408 9982 17408 0 VGND
rlabel via1 9982 16864 9982 16864 0 VPWR
rlabel metal2 16698 8670 16698 8670 0 _000_
rlabel metal1 11921 7786 11921 7786 0 _001_
rlabel metal1 11093 6698 11093 6698 0 _002_
rlabel metal1 12328 10778 12328 10778 0 _003_
rlabel metal1 13623 8942 13623 8942 0 _004_
rlabel metal1 14221 7446 14221 7446 0 _005_
rlabel metal2 15686 9724 15686 9724 0 _006_
rlabel metal2 16790 8364 16790 8364 0 _007_
rlabel metal1 15916 13158 15916 13158 0 _008_
rlabel metal1 18262 12682 18262 12682 0 _009_
rlabel metal1 17480 12614 17480 12614 0 _010_
rlabel metal2 15180 8228 15180 8228 0 _011_
rlabel metal1 16836 11050 16836 11050 0 _012_
rlabel metal1 17027 9962 17027 9962 0 _013_
rlabel metal1 16698 11662 16698 11662 0 _014_
rlabel metal1 7643 3434 7643 3434 0 _015_
rlabel metal2 15594 9146 15594 9146 0 _016_
rlabel metal2 16146 8840 16146 8840 0 _017_
rlabel metal2 12282 5576 12282 5576 0 _018_
rlabel metal1 16238 14246 16238 14246 0 _019_
rlabel via2 10718 4539 10718 4539 0 _020_
rlabel metal1 17756 12954 17756 12954 0 _021_
rlabel metal2 14674 5882 14674 5882 0 _022_
rlabel metal1 13570 8568 13570 8568 0 _023_
rlabel metal1 12282 7922 12282 7922 0 _024_
rlabel metal1 11276 6970 11276 6970 0 _025_
rlabel via1 7399 10438 7399 10438 0 _026_
rlabel metal2 11914 9690 11914 9690 0 _027_
rlabel metal1 13524 7310 13524 7310 0 _028_
rlabel metal1 14628 8874 14628 8874 0 _029_
rlabel metal2 15686 5474 15686 5474 0 _030_
rlabel metal1 17673 2618 17673 2618 0 _031_
rlabel metal1 15732 3434 15732 3434 0 _032_
rlabel metal2 14306 4930 14306 4930 0 _033_
rlabel metal2 14398 6086 14398 6086 0 _034_
rlabel metal2 15870 9758 15870 9758 0 _035_
rlabel metal1 17342 9146 17342 9146 0 _036_
rlabel metal1 16054 7310 16054 7310 0 _037_
rlabel metal2 12006 5406 12006 5406 0 _038_
rlabel metal2 12190 3298 12190 3298 0 _039_
rlabel metal1 11730 4658 11730 4658 0 _040_
rlabel metal2 14766 3502 14766 3502 0 _041_
rlabel metal2 11822 6188 11822 6188 0 _042_
rlabel metal1 4370 13396 4370 13396 0 _043_
rlabel metal1 9660 2414 9660 2414 0 _044_
rlabel metal2 9154 2074 9154 2074 0 _045_
rlabel metal1 13846 7854 13846 7854 0 _046_
rlabel metal1 18630 6834 18630 6834 0 _047_
rlabel metal1 18400 8466 18400 8466 0 _048_
rlabel metal1 17434 5066 17434 5066 0 _049_
rlabel metal2 14766 6290 14766 6290 0 _050_
rlabel metal1 14812 4590 14812 4590 0 _051_
rlabel metal1 15318 13226 15318 13226 0 _052_
rlabel metal2 17342 10880 17342 10880 0 _053_
rlabel metal1 18469 10098 18469 10098 0 _054_
rlabel metal1 18538 4114 18538 4114 0 _055_
rlabel metal1 4922 14994 4922 14994 0 _056_
rlabel metal1 9108 12138 9108 12138 0 _057_
rlabel metal1 8004 12206 8004 12206 0 _058_
rlabel metal2 4646 11356 4646 11356 0 _059_
rlabel metal1 16698 14314 16698 14314 0 _060_
rlabel metal2 13340 2414 13340 2414 0 _061_
rlabel metal1 13478 12274 13478 12274 0 _062_
rlabel metal1 18906 2414 18906 2414 0 _063_
rlabel metal1 12374 2346 12374 2346 0 _064_
rlabel metal1 11776 2414 11776 2414 0 _065_
rlabel metal1 13892 14042 13892 14042 0 _066_
rlabel metal1 10836 2414 10836 2414 0 _067_
rlabel metal1 11868 2482 11868 2482 0 _068_
rlabel metal2 12282 2176 12282 2176 0 _069_
rlabel metal1 10764 2482 10764 2482 0 _070_
rlabel metal2 12926 2754 12926 2754 0 _071_
rlabel via2 17986 9435 17986 9435 0 _072_
rlabel metal1 16882 2482 16882 2482 0 _073_
rlabel metal1 10994 14280 10994 14280 0 _074_
rlabel metal1 9706 3026 9706 3026 0 _075_
rlabel metal1 14582 3434 14582 3434 0 _076_
rlabel metal1 17296 3026 17296 3026 0 _077_
rlabel metal1 16974 13838 16974 13838 0 _078_
rlabel metal1 17296 2482 17296 2482 0 _079_
rlabel metal1 9384 2414 9384 2414 0 _080_
rlabel metal1 9430 2516 9430 2516 0 _081_
rlabel metal1 9522 2346 9522 2346 0 _082_
rlabel metal1 7820 2618 7820 2618 0 _083_
rlabel metal1 8326 2482 8326 2482 0 _084_
rlabel metal2 7590 1972 7590 1972 0 _085_
rlabel metal1 8004 3094 8004 3094 0 _086_
rlabel via2 6302 14467 6302 14467 0 _087_
rlabel metal1 5382 4046 5382 4046 0 _088_
rlabel via2 14306 3451 14306 3451 0 _089_
rlabel metal1 6808 14246 6808 14246 0 _090_
rlabel metal1 10534 2312 10534 2312 0 _091_
rlabel metal2 16698 4131 16698 4131 0 _092_
rlabel metal1 7360 3162 7360 3162 0 _093_
rlabel metal1 17848 4590 17848 4590 0 _094_
rlabel metal1 17779 5678 17779 5678 0 _095_
rlabel metal1 10304 12750 10304 12750 0 _096_
rlabel metal2 10810 12988 10810 12988 0 _097_
rlabel metal2 11086 12619 11086 12619 0 _098_
rlabel metal1 10074 12274 10074 12274 0 _099_
rlabel metal1 12052 13294 12052 13294 0 _100_
rlabel metal1 11684 12070 11684 12070 0 _101_
rlabel metal1 12006 13362 12006 13362 0 _102_
rlabel metal1 12696 12886 12696 12886 0 _103_
rlabel metal1 13478 12614 13478 12614 0 _104_
rlabel via1 12719 11730 12719 11730 0 _105_
rlabel metal1 9752 2618 9752 2618 0 _106_
rlabel via1 14674 4811 14674 4811 0 _107_
rlabel metal2 18170 8823 18170 8823 0 _108_
rlabel metal1 12604 13498 12604 13498 0 _109_
rlabel metal1 3450 14858 3450 14858 0 _110_
rlabel metal1 9844 11118 9844 11118 0 _111_
rlabel metal1 5106 12342 5106 12342 0 _112_
rlabel metal1 8142 11628 8142 11628 0 _113_
rlabel metal1 9660 9010 9660 9010 0 _114_
rlabel metal2 9798 7650 9798 7650 0 _115_
rlabel metal2 15410 7259 15410 7259 0 _116_
rlabel metal1 13156 10642 13156 10642 0 _117_
rlabel metal1 10856 8058 10856 8058 0 _118_
rlabel metal1 13570 10982 13570 10982 0 _119_
rlabel metal2 12006 12682 12006 12682 0 _120_
rlabel metal1 13570 11866 13570 11866 0 _121_
rlabel metal1 14306 11152 14306 11152 0 _122_
rlabel metal2 12374 10948 12374 10948 0 _123_
rlabel viali 8970 11728 8970 11728 0 _124_
rlabel metal2 9798 11917 9798 11917 0 _125_
rlabel metal1 8372 11186 8372 11186 0 _126_
rlabel metal1 10534 10166 10534 10166 0 _127_
rlabel metal1 11914 9690 11914 9690 0 _128_
rlabel metal2 3726 15606 3726 15606 0 _129_
rlabel via2 10718 9435 10718 9435 0 _130_
rlabel metal1 15042 9588 15042 9588 0 _131_
rlabel metal1 12374 9418 12374 9418 0 _132_
rlabel via2 1978 13243 1978 13243 0 _133_
rlabel metal1 3174 14382 3174 14382 0 _134_
rlabel metal1 2990 10744 2990 10744 0 _135_
rlabel metal1 5520 2482 5520 2482 0 _136_
rlabel metal2 2714 15521 2714 15521 0 _137_
rlabel metal2 4002 10880 4002 10880 0 _138_
rlabel metal1 6118 11084 6118 11084 0 _139_
rlabel metal1 6716 12818 6716 12818 0 _140_
rlabel metal1 7406 13838 7406 13838 0 _141_
rlabel metal2 7958 13260 7958 13260 0 _142_
rlabel metal1 5014 5338 5014 5338 0 _143_
rlabel metal1 1748 13974 1748 13974 0 _144_
rlabel via2 5566 7293 5566 7293 0 _145_
rlabel metal2 4370 13090 4370 13090 0 _146_
rlabel metal1 6992 15402 6992 15402 0 _147_
rlabel metal1 4370 14994 4370 14994 0 _148_
rlabel metal2 2346 13175 2346 13175 0 _149_
rlabel metal1 3956 10438 3956 10438 0 _150_
rlabel metal2 6486 11424 6486 11424 0 _151_
rlabel metal2 5382 15232 5382 15232 0 _152_
rlabel metal1 4600 15878 4600 15878 0 _153_
rlabel metal1 6808 2618 6808 2618 0 _154_
rlabel metal2 4370 14824 4370 14824 0 _155_
rlabel metal1 2346 13940 2346 13940 0 _156_
rlabel metal1 3864 14042 3864 14042 0 _157_
rlabel metal1 4922 11866 4922 11866 0 _158_
rlabel metal1 4784 15878 4784 15878 0 _159_
rlabel metal1 5980 2278 5980 2278 0 _160_
rlabel metal2 14858 8415 14858 8415 0 _161_
rlabel metal2 9982 8772 9982 8772 0 _162_
rlabel metal1 4219 11730 4219 11730 0 _163_
rlabel metal1 2806 11220 2806 11220 0 _164_
rlabel metal1 2484 11798 2484 11798 0 _165_
rlabel via2 2346 12291 2346 12291 0 _166_
rlabel metal2 1472 12614 1472 12614 0 _167_
rlabel metal2 3266 14892 3266 14892 0 _168_
rlabel metal1 12742 7242 12742 7242 0 _169_
rlabel via1 5566 12189 5566 12189 0 _170_
rlabel metal1 5520 12138 5520 12138 0 _171_
rlabel metal1 6302 5134 6302 5134 0 _172_
rlabel metal1 5382 9554 5382 9554 0 _173_
rlabel metal3 2062 476 2062 476 0 clockp[0]
rlabel metal3 2384 204 2384 204 0 clockp[1]
rlabel metal1 3036 2550 3036 2550 0 dco
rlabel metal3 2062 1836 2062 1836 0 div[0]
rlabel metal3 2108 1564 2108 1564 0 div[1]
rlabel metal3 912 1292 912 1292 0 div[2]
rlabel metal3 2108 1020 2108 1020 0 div[3]
rlabel metal3 2016 748 2016 748 0 div[4]
rlabel metal3 866 2108 866 2108 0 enable
rlabel metal3 820 4284 820 4284 0 ext_trim[0]
rlabel metal1 7636 12886 7636 12886 0 ext_trim[10]
rlabel metal1 552 15266 552 15266 0 ext_trim[11]
rlabel metal1 1564 14382 1564 14382 0 ext_trim[12]
rlabel metal1 1564 15062 1564 15062 0 ext_trim[13]
rlabel metal1 4784 17510 4784 17510 0 ext_trim[14]
rlabel metal2 1380 12716 1380 12716 0 ext_trim[15]
rlabel metal1 1538 13906 1538 13906 0 ext_trim[16]
rlabel via1 2245 12750 2245 12750 0 ext_trim[17]
rlabel metal1 1508 12274 1508 12274 0 ext_trim[18]
rlabel via1 2878 13294 2878 13294 0 ext_trim[19]
rlabel metal3 1050 4012 1050 4012 0 ext_trim[1]
rlabel metal2 15870 1785 15870 1785 0 ext_trim[20]
rlabel via2 15410 1275 15410 1275 0 ext_trim[21]
rlabel metal1 16146 8432 16146 8432 0 ext_trim[22]
rlabel metal3 19144 748 19144 748 0 ext_trim[23]
rlabel metal3 19190 476 19190 476 0 ext_trim[24]
rlabel metal2 19136 204 19136 204 0 ext_trim[25]
rlabel metal1 1288 16082 1288 16082 0 ext_trim[2]
rlabel metal1 1288 16558 1288 16558 0 ext_trim[3]
rlabel metal1 920 13838 920 13838 0 ext_trim[4]
rlabel metal1 966 15402 966 15402 0 ext_trim[5]
rlabel metal3 1027 2652 1027 2652 0 ext_trim[6]
rlabel metal2 138 16058 138 16058 0 ext_trim[7]
rlabel metal2 322 17384 322 17384 0 ext_trim[8]
rlabel metal1 2898 16014 2898 16014 0 ext_trim[9]
rlabel metal2 322 874 322 874 0 osc
rlabel metal1 6026 3468 6026 3468 0 pll_control.clock
rlabel metal1 14582 12784 14582 12784 0 pll_control.count0\[0\]
rlabel metal1 14490 2618 14490 2618 0 pll_control.count0\[1\]
rlabel metal1 17112 3570 17112 3570 0 pll_control.count0\[2\]
rlabel metal1 14674 13974 14674 13974 0 pll_control.count0\[3\]
rlabel metal1 14674 13294 14674 13294 0 pll_control.count0\[4\]
rlabel metal1 13616 12818 13616 12818 0 pll_control.count1\[0\]
rlabel metal1 13478 4114 13478 4114 0 pll_control.count1\[1\]
rlabel metal1 14766 12138 14766 12138 0 pll_control.count1\[2\]
rlabel metal1 17296 13906 17296 13906 0 pll_control.count1\[3\]
rlabel metal1 9338 5882 9338 5882 0 pll_control.count1\[4\]
rlabel metal2 14858 5848 14858 5848 0 pll_control.oscbuf\[0\]
rlabel metal2 16054 6188 16054 6188 0 pll_control.oscbuf\[1\]
rlabel metal2 17802 6528 17802 6528 0 pll_control.oscbuf\[2\]
rlabel metal1 18492 8942 18492 8942 0 pll_control.prep\[0\]
rlabel metal1 17572 8942 17572 8942 0 pll_control.prep\[1\]
rlabel metal1 17802 7242 17802 7242 0 pll_control.prep\[2\]
rlabel metal1 9200 6970 9200 6970 0 pll_control.tint\[0\]
rlabel metal1 4370 11764 4370 11764 0 pll_control.tint\[1\]
rlabel metal2 13202 9248 13202 9248 0 pll_control.tint\[2\]
rlabel metal1 5014 13294 5014 13294 0 pll_control.tint\[3\]
rlabel metal1 12926 11084 12926 11084 0 pll_control.tint\[4\]
rlabel metal1 13110 10064 13110 10064 0 pll_control.tval\[0\]
rlabel metal1 8510 11798 8510 11798 0 pll_control.tval\[1\]
rlabel metal1 276 13022 276 13022 0 resetb
rlabel metal2 5198 7140 5198 7140 0 ringosc.c\[0\]
rlabel metal2 5382 2587 5382 2587 0 ringosc.c\[1\]
rlabel metal1 2645 3978 2645 3978 0 ringosc.dstage\[0\].id.d0
rlabel metal2 3082 4420 3082 4420 0 ringosc.dstage\[0\].id.d1
rlabel metal2 2714 4386 2714 4386 0 ringosc.dstage\[0\].id.d2
rlabel metal1 1518 2618 1518 2618 0 ringosc.dstage\[0\].id.in
rlabel metal1 1702 5168 1702 5168 0 ringosc.dstage\[0\].id.out
rlabel metal1 5566 4624 5566 4624 0 ringosc.dstage\[0\].id.trim\[0\]
rlabel metal1 1656 14790 1656 14790 0 ringosc.dstage\[0\].id.trim\[1\]
rlabel metal2 2346 4284 2346 4284 0 ringosc.dstage\[0\].id.ts
rlabel metal1 8326 5576 8326 5576 0 ringosc.dstage\[10\].id.d0
rlabel metal1 8188 5610 8188 5610 0 ringosc.dstage\[10\].id.d1
rlabel metal1 8694 5270 8694 5270 0 ringosc.dstage\[10\].id.d2
rlabel metal1 9200 6154 9200 6154 0 ringosc.dstage\[10\].id.in
rlabel metal1 9200 5066 9200 5066 0 ringosc.dstage\[10\].id.out
rlabel metal1 7636 5134 7636 5134 0 ringosc.dstage\[10\].id.trim\[0\]
rlabel metal1 13409 7786 13409 7786 0 ringosc.dstage\[10\].id.trim\[1\]
rlabel metal1 7452 5202 7452 5202 0 ringosc.dstage\[10\].id.ts
rlabel metal1 8326 4488 8326 4488 0 ringosc.dstage\[11\].id.d0
rlabel metal1 8188 4522 8188 4522 0 ringosc.dstage\[11\].id.d1
rlabel metal2 8234 4420 8234 4420 0 ringosc.dstage\[11\].id.d2
rlabel metal1 1610 3434 1610 3434 0 ringosc.dstage\[11\].id.out
rlabel via1 1426 3893 1426 3893 0 ringosc.dstage\[11\].id.trim\[0\]
rlabel metal1 6670 4114 6670 4114 0 ringosc.dstage\[11\].id.trim\[1\]
rlabel metal1 7222 4114 7222 4114 0 ringosc.dstage\[11\].id.ts
rlabel metal1 2990 5100 2990 5100 0 ringosc.dstage\[1\].id.d0
rlabel metal1 1702 5576 1702 5576 0 ringosc.dstage\[1\].id.d1
rlabel metal2 4186 5542 4186 5542 0 ringosc.dstage\[1\].id.d2
rlabel metal1 1702 6256 1702 6256 0 ringosc.dstage\[1\].id.out
rlabel metal1 3266 16490 3266 16490 0 ringosc.dstage\[1\].id.trim\[0\]
rlabel metal1 2162 5780 2162 5780 0 ringosc.dstage\[1\].id.trim\[1\]
rlabel metal2 2346 5406 2346 5406 0 ringosc.dstage\[1\].id.ts
rlabel metal1 2990 6188 2990 6188 0 ringosc.dstage\[2\].id.d0
rlabel metal2 2254 6528 2254 6528 0 ringosc.dstage\[2\].id.d1
rlabel metal2 2714 6562 2714 6562 0 ringosc.dstage\[2\].id.d2
rlabel metal1 3404 6698 3404 6698 0 ringosc.dstage\[2\].id.out
rlabel metal2 3174 14246 3174 14246 0 ringosc.dstage\[2\].id.trim\[0\]
rlabel metal1 2668 6766 2668 6766 0 ringosc.dstage\[2\].id.trim\[1\]
rlabel metal1 1610 6800 1610 6800 0 ringosc.dstage\[2\].id.ts
rlabel metal1 2645 7242 2645 7242 0 ringosc.dstage\[3\].id.d0
rlabel metal1 1702 7752 1702 7752 0 ringosc.dstage\[3\].id.d1
rlabel metal2 2714 7650 2714 7650 0 ringosc.dstage\[3\].id.d2
rlabel metal1 1702 8432 1702 8432 0 ringosc.dstage\[3\].id.out
rlabel metal1 3496 7854 3496 7854 0 ringosc.dstage\[3\].id.trim\[0\]
rlabel metal1 1518 13702 1518 13702 0 ringosc.dstage\[3\].id.trim\[1\]
rlabel metal1 1610 7888 1610 7888 0 ringosc.dstage\[3\].id.ts
rlabel metal1 2990 8364 2990 8364 0 ringosc.dstage\[4\].id.d0
rlabel metal2 2254 8704 2254 8704 0 ringosc.dstage\[4\].id.d1
rlabel metal2 2714 8738 2714 8738 0 ringosc.dstage\[4\].id.d2
rlabel metal1 1702 9520 1702 9520 0 ringosc.dstage\[4\].id.out
rlabel metal1 2990 13702 2990 13702 0 ringosc.dstage\[4\].id.trim\[0\]
rlabel metal1 2484 12614 2484 12614 0 ringosc.dstage\[4\].id.trim\[1\]
rlabel metal1 1610 8976 1610 8976 0 ringosc.dstage\[4\].id.ts
rlabel metal1 2990 9452 2990 9452 0 ringosc.dstage\[5\].id.d0
rlabel metal2 2438 9758 2438 9758 0 ringosc.dstage\[5\].id.d1
rlabel metal2 2714 9792 2714 9792 0 ringosc.dstage\[5\].id.d2
rlabel metal1 8556 3502 8556 3502 0 ringosc.dstage\[5\].id.out
rlabel metal1 2162 15368 2162 15368 0 ringosc.dstage\[5\].id.trim\[0\]
rlabel metal2 2530 11985 2530 11985 0 ringosc.dstage\[5\].id.trim\[1\]
rlabel metal2 2346 9826 2346 9826 0 ringosc.dstage\[5\].id.ts
rlabel metal1 8326 9928 8326 9928 0 ringosc.dstage\[6\].id.d0
rlabel metal1 8188 9962 8188 9962 0 ringosc.dstage\[6\].id.d1
rlabel metal1 8694 9622 8694 9622 0 ringosc.dstage\[6\].id.d2
rlabel metal1 9200 9418 9200 9418 0 ringosc.dstage\[6\].id.out
rlabel metal1 7314 9486 7314 9486 0 ringosc.dstage\[6\].id.trim\[0\]
rlabel metal2 6854 11356 6854 11356 0 ringosc.dstage\[6\].id.trim\[1\]
rlabel metal1 7222 9554 7222 9554 0 ringosc.dstage\[6\].id.ts
rlabel metal1 8326 8840 8326 8840 0 ringosc.dstage\[7\].id.d0
rlabel metal1 8188 8874 8188 8874 0 ringosc.dstage\[7\].id.d1
rlabel metal1 8740 8534 8740 8534 0 ringosc.dstage\[7\].id.d2
rlabel metal1 9200 8330 9200 8330 0 ringosc.dstage\[7\].id.out
rlabel metal2 5198 12546 5198 12546 0 ringosc.dstage\[7\].id.trim\[0\]
rlabel metal1 6578 8398 6578 8398 0 ringosc.dstage\[7\].id.trim\[1\]
rlabel metal1 7360 8466 7360 8466 0 ringosc.dstage\[7\].id.ts
rlabel metal1 8326 7752 8326 7752 0 ringosc.dstage\[8\].id.d0
rlabel metal1 8188 7786 8188 7786 0 ringosc.dstage\[8\].id.d1
rlabel metal1 8740 7446 8740 7446 0 ringosc.dstage\[8\].id.d2
rlabel metal1 9200 7242 9200 7242 0 ringosc.dstage\[8\].id.out
rlabel metal1 5796 15538 5796 15538 0 ringosc.dstage\[8\].id.trim\[0\]
rlabel metal1 6716 7378 6716 7378 0 ringosc.dstage\[8\].id.trim\[1\]
rlabel metal1 7222 7378 7222 7378 0 ringosc.dstage\[8\].id.ts
rlabel metal1 8326 6664 8326 6664 0 ringosc.dstage\[9\].id.d0
rlabel metal1 8188 6698 8188 6698 0 ringosc.dstage\[9\].id.d1
rlabel metal1 8740 6358 8740 6358 0 ringosc.dstage\[9\].id.d2
rlabel metal1 7590 6222 7590 6222 0 ringosc.dstage\[9\].id.trim\[0\]
rlabel metal2 13018 7786 13018 7786 0 ringosc.dstage\[9\].id.trim\[1\]
rlabel metal1 7452 6290 7452 6290 0 ringosc.dstage\[9\].id.ts
rlabel metal1 3634 2618 3634 2618 0 ringosc.iss.ctrl0
rlabel metal1 2346 2924 2346 2924 0 ringosc.iss.d0
rlabel metal2 2438 3264 2438 3264 0 ringosc.iss.d1
rlabel metal2 2714 3298 2714 3298 0 ringosc.iss.d2
rlabel metal1 2898 2482 2898 2482 0 ringosc.iss.one
rlabel metal1 2576 2414 2576 2414 0 ringosc.iss.reset
rlabel metal1 1564 14314 1564 14314 0 ringosc.iss.trim\[0\]
rlabel metal1 3174 3468 3174 3468 0 ringosc.iss.trim\[1\]
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
