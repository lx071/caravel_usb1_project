magic
tech sky130A
magscale 1 2
timestamp 1698809212
<< obsli1 >>
rect 1104 2159 88872 77809
<< obsm1 >>
rect 106 76 89134 79756
<< metal2 >>
rect 110 79200 166 80800
rect 294 79200 350 80800
rect 478 79200 534 80800
rect 662 79200 718 80800
rect 846 79200 902 80800
rect 1030 79200 1086 80800
rect 1214 79200 1270 80800
rect 1398 79200 1454 80800
rect 20074 79200 20130 80800
rect 24030 79200 24086 80800
rect 24214 79200 24270 80800
rect 24398 79200 24454 80800
rect 24582 79200 24638 80800
rect 24766 79200 24822 80800
rect 24950 79200 25006 80800
rect 25134 79200 25190 80800
rect 25318 79200 25374 80800
rect 25502 79200 25558 80800
rect 25686 79200 25742 80800
rect 25870 79200 25926 80800
rect 26054 79200 26110 80800
rect 26238 79200 26294 80800
rect 26422 79200 26478 80800
rect 26606 79200 26662 80800
rect 26790 79200 26846 80800
rect 26974 79200 27030 80800
rect 27158 79200 27214 80800
rect 27342 79200 27398 80800
rect 27526 79200 27582 80800
rect 27710 79200 27766 80800
rect 27894 79200 27950 80800
rect 28078 79200 28134 80800
rect 28262 79200 28318 80800
rect 28446 79200 28502 80800
rect 28630 79200 28686 80800
rect 28814 79200 28870 80800
rect 28998 79200 29054 80800
rect 29182 79200 29238 80800
rect 29366 79200 29422 80800
rect 29550 79200 29606 80800
rect 29734 79200 29790 80800
rect 29918 79200 29974 80800
rect 30102 79200 30158 80800
rect 30286 79200 30342 80800
rect 30470 79200 30526 80800
rect 30654 79200 30710 80800
rect 30838 79200 30894 80800
rect 31022 79200 31078 80800
rect 31206 79200 31262 80800
rect 31390 79200 31446 80800
rect 31574 79200 31630 80800
rect 31758 79200 31814 80800
rect 31942 79200 31998 80800
rect 32126 79200 32182 80800
rect 32310 79200 32366 80800
rect 32494 79200 32550 80800
rect 32678 79200 32734 80800
rect 32862 79200 32918 80800
rect 33046 79200 33102 80800
rect 33230 79200 33286 80800
rect 33414 79200 33470 80800
rect 33598 79200 33654 80800
rect 40038 79200 40094 80800
rect 40222 79200 40278 80800
rect 40406 79200 40462 80800
rect 40590 79200 40646 80800
rect 40774 79200 40830 80800
rect 40958 79200 41014 80800
rect 41142 79200 41198 80800
rect 41326 79200 41382 80800
rect 41510 79200 41566 80800
rect 41694 79200 41750 80800
rect 41878 79200 41934 80800
rect 42062 79200 42118 80800
rect 42246 79200 42302 80800
rect 42430 79200 42486 80800
rect 42614 79200 42670 80800
rect 42798 79200 42854 80800
rect 42982 79200 43038 80800
rect 43166 79200 43222 80800
rect 43350 79200 43406 80800
rect 43534 79200 43590 80800
rect 43718 79200 43774 80800
rect 43902 79200 43958 80800
rect 44086 79200 44142 80800
rect 44270 79200 44326 80800
rect 44454 79200 44510 80800
rect 44638 79200 44694 80800
rect 44822 79200 44878 80800
rect 45006 79200 45062 80800
rect 45190 79200 45246 80800
rect 45374 79200 45430 80800
rect 45558 79200 45614 80800
rect 45742 79200 45798 80800
rect 45926 79200 45982 80800
rect 46110 79200 46166 80800
rect 46294 79200 46350 80800
rect 46478 79200 46534 80800
rect 46662 79200 46718 80800
rect 46846 79200 46902 80800
rect 47030 79200 47086 80800
rect 47214 79200 47270 80800
rect 47398 79200 47454 80800
rect 47582 79200 47638 80800
rect 47766 79200 47822 80800
rect 47950 79200 48006 80800
rect 48134 79200 48190 80800
rect 48318 79200 48374 80800
rect 48502 79200 48558 80800
rect 48686 79200 48742 80800
rect 48870 79200 48926 80800
rect 49054 79200 49110 80800
rect 49238 79200 49294 80800
rect 49422 79200 49478 80800
rect 49606 79200 49662 80800
rect 49790 79200 49846 80800
rect 49974 79200 50030 80800
rect 50158 79200 50214 80800
rect 50342 79200 50398 80800
rect 50526 79200 50582 80800
rect 50710 79200 50766 80800
rect 50894 79200 50950 80800
rect 51078 79200 51134 80800
rect 51262 79200 51318 80800
rect 51446 79200 51502 80800
rect 51630 79200 51686 80800
rect 51814 79200 51870 80800
rect 51998 79200 52054 80800
rect 52182 79200 52238 80800
rect 52366 79200 52422 80800
rect 52550 79200 52606 80800
rect 52734 79200 52790 80800
rect 52918 79200 52974 80800
rect 53102 79200 53158 80800
rect 53286 79200 53342 80800
rect 53470 79200 53526 80800
rect 53654 79200 53710 80800
rect 53838 79200 53894 80800
rect 54022 79200 54078 80800
rect 54206 79200 54262 80800
rect 54390 79200 54446 80800
rect 54574 79200 54630 80800
rect 54758 79200 54814 80800
rect 54942 79200 54998 80800
rect 55126 79200 55182 80800
rect 55310 79200 55366 80800
rect 55494 79200 55550 80800
rect 55678 79200 55734 80800
rect 55862 79200 55918 80800
rect 56046 79200 56102 80800
rect 56230 79200 56286 80800
rect 56414 79200 56470 80800
rect 56598 79200 56654 80800
rect 56782 79200 56838 80800
rect 56966 79200 57022 80800
rect 57150 79200 57206 80800
rect 57334 79200 57390 80800
rect 57518 79200 57574 80800
rect 57702 79200 57758 80800
rect 57886 79200 57942 80800
rect 58070 79200 58126 80800
rect 58254 79200 58310 80800
rect 58438 79200 58494 80800
rect 58622 79200 58678 80800
rect 58806 79200 58862 80800
rect 58990 79200 59046 80800
rect 59174 79200 59230 80800
rect 65062 79200 65118 80800
rect 65246 79200 65302 80800
rect 65430 79200 65486 80800
rect 65614 79200 65670 80800
rect 65798 79200 65854 80800
rect 65982 79200 66038 80800
rect 66166 79200 66222 80800
rect 66350 79200 66406 80800
rect 66534 79200 66590 80800
rect 66718 79200 66774 80800
rect 66902 79200 66958 80800
rect 67086 79200 67142 80800
rect 67270 79200 67326 80800
rect 67454 79200 67510 80800
rect 67638 79200 67694 80800
rect 67822 79200 67878 80800
rect 68006 79200 68062 80800
rect 68190 79200 68246 80800
rect 68374 79200 68430 80800
rect 68558 79200 68614 80800
rect 68742 79200 68798 80800
rect 68926 79200 68982 80800
rect 69110 79200 69166 80800
rect 69294 79200 69350 80800
rect 69478 79200 69534 80800
rect 69662 79200 69718 80800
rect 69846 79200 69902 80800
rect 70030 79200 70086 80800
rect 70214 79200 70270 80800
rect 70398 79200 70454 80800
rect 70582 79200 70638 80800
rect 70766 79200 70822 80800
rect 70950 79200 71006 80800
rect 71134 79200 71190 80800
rect 71318 79200 71374 80800
rect 71502 79200 71558 80800
rect 71686 79200 71742 80800
rect 71870 79200 71926 80800
rect 72054 79200 72110 80800
rect 72238 79200 72294 80800
rect 72422 79200 72478 80800
rect 72606 79200 72662 80800
rect 72790 79200 72846 80800
rect 72974 79200 73030 80800
rect 73158 79200 73214 80800
rect 73342 79200 73398 80800
rect 73526 79200 73582 80800
rect 73710 79200 73766 80800
rect 73894 79200 73950 80800
rect 74078 79200 74134 80800
rect 74262 79200 74318 80800
rect 74446 79200 74502 80800
rect 74630 79200 74686 80800
rect 74814 79200 74870 80800
rect 74998 79200 75054 80800
rect 75182 79200 75238 80800
rect 75366 79200 75422 80800
rect 75550 79200 75606 80800
rect 75734 79200 75790 80800
rect 75918 79200 75974 80800
rect 76102 79200 76158 80800
rect 76286 79200 76342 80800
rect 76470 79200 76526 80800
rect 76654 79200 76710 80800
rect 76838 79200 76894 80800
rect 77022 79200 77078 80800
rect 77206 79200 77262 80800
rect 77390 79200 77446 80800
rect 77574 79200 77630 80800
rect 77758 79200 77814 80800
rect 77942 79200 77998 80800
rect 78126 79200 78182 80800
rect 78310 79200 78366 80800
rect 78494 79200 78550 80800
rect 78678 79200 78734 80800
rect 78862 79200 78918 80800
rect 79046 79200 79102 80800
rect 79230 79200 79286 80800
rect 79414 79200 79470 80800
rect 79598 79200 79654 80800
rect 79782 79200 79838 80800
rect 79966 79200 80022 80800
rect 80150 79200 80206 80800
rect 80334 79200 80390 80800
rect 110 -800 166 800
rect 294 -800 350 800
rect 478 -800 534 800
rect 662 -800 718 800
rect 846 -800 902 800
rect 1030 -800 1086 800
rect 1214 -800 1270 800
rect 1398 -800 1454 800
rect 1582 -800 1638 800
rect 1766 -800 1822 800
rect 1950 -800 2006 800
rect 2134 -800 2190 800
rect 2318 -800 2374 800
rect 2502 -800 2558 800
rect 2686 -800 2742 800
rect 2870 -800 2926 800
rect 3054 -800 3110 800
rect 3238 -800 3294 800
rect 3422 -800 3478 800
rect 3606 -800 3662 800
rect 3790 -800 3846 800
rect 3974 -800 4030 800
rect 4158 -800 4214 800
rect 4342 -800 4398 800
rect 4526 -800 4582 800
rect 4710 -800 4766 800
rect 4894 -800 4950 800
rect 5078 -800 5134 800
rect 5262 -800 5318 800
rect 5446 -800 5502 800
rect 5630 -800 5686 800
rect 5814 -800 5870 800
rect 5998 -800 6054 800
rect 6182 -800 6238 800
rect 6366 -800 6422 800
rect 6550 -800 6606 800
rect 6734 -800 6790 800
rect 6918 -800 6974 800
rect 7102 -800 7158 800
rect 7286 -800 7342 800
rect 7470 -800 7526 800
rect 7654 -800 7710 800
rect 7838 -800 7894 800
rect 8022 -800 8078 800
rect 8206 -800 8262 800
rect 8390 -800 8446 800
rect 8574 -800 8630 800
rect 8758 -800 8814 800
rect 8942 -800 8998 800
rect 9126 -800 9182 800
rect 9310 -800 9366 800
rect 9494 -800 9550 800
rect 9678 -800 9734 800
rect 9862 -800 9918 800
rect 10046 -800 10102 800
rect 10230 -800 10286 800
rect 10414 -800 10470 800
rect 10598 -800 10654 800
rect 10782 -800 10838 800
rect 10966 -800 11022 800
rect 11150 -800 11206 800
rect 11334 -800 11390 800
rect 11518 -800 11574 800
rect 11702 -800 11758 800
rect 11886 -800 11942 800
rect 12070 -800 12126 800
rect 12254 -800 12310 800
rect 12438 -800 12494 800
rect 12622 -800 12678 800
rect 12806 -800 12862 800
rect 12990 -800 13046 800
rect 13174 -800 13230 800
rect 13358 -800 13414 800
rect 13542 -800 13598 800
rect 13726 -800 13782 800
rect 13910 -800 13966 800
rect 14094 -800 14150 800
rect 14278 -800 14334 800
rect 14462 -800 14518 800
rect 14646 -800 14702 800
rect 14830 -800 14886 800
rect 15014 -800 15070 800
rect 15198 -800 15254 800
rect 15382 -800 15438 800
rect 15566 -800 15622 800
rect 15750 -800 15806 800
rect 15934 -800 15990 800
rect 16118 -800 16174 800
rect 16302 -800 16358 800
rect 16486 -800 16542 800
rect 16670 -800 16726 800
rect 16854 -800 16910 800
rect 17038 -800 17094 800
rect 17222 -800 17278 800
rect 17406 -800 17462 800
rect 17590 -800 17646 800
rect 17774 -800 17830 800
rect 17958 -800 18014 800
rect 18142 -800 18198 800
rect 18326 -800 18382 800
rect 18510 -800 18566 800
rect 18694 -800 18750 800
rect 18878 -800 18934 800
rect 19062 -800 19118 800
rect 19246 -800 19302 800
rect 19430 -800 19486 800
rect 19614 -800 19670 800
rect 19798 -800 19854 800
rect 19982 -800 20038 800
rect 50066 -800 50122 800
rect 50250 -800 50306 800
rect 50434 -800 50490 800
rect 50618 -800 50674 800
rect 50802 -800 50858 800
rect 50986 -800 51042 800
rect 51170 -800 51226 800
rect 51354 -800 51410 800
rect 51538 -800 51594 800
rect 51722 -800 51778 800
rect 51906 -800 51962 800
rect 52090 -800 52146 800
rect 52274 -800 52330 800
rect 52458 -800 52514 800
rect 52642 -800 52698 800
rect 52826 -800 52882 800
rect 53010 -800 53066 800
rect 53194 -800 53250 800
<< obsm2 >>
rect 222 79144 238 79762
rect 406 79144 422 79762
rect 590 79144 606 79762
rect 774 79144 790 79762
rect 958 79144 974 79762
rect 1142 79144 1158 79762
rect 1326 79144 1342 79762
rect 1510 79144 20018 79762
rect 20186 79144 23974 79762
rect 24142 79144 24158 79762
rect 24326 79144 24342 79762
rect 24510 79144 24526 79762
rect 24694 79144 24710 79762
rect 24878 79144 24894 79762
rect 25062 79144 25078 79762
rect 25246 79144 25262 79762
rect 25430 79144 25446 79762
rect 25614 79144 25630 79762
rect 25798 79144 25814 79762
rect 25982 79144 25998 79762
rect 26166 79144 26182 79762
rect 26350 79144 26366 79762
rect 26534 79144 26550 79762
rect 26718 79144 26734 79762
rect 26902 79144 26918 79762
rect 27086 79144 27102 79762
rect 27270 79144 27286 79762
rect 27454 79144 27470 79762
rect 27638 79144 27654 79762
rect 27822 79144 27838 79762
rect 28006 79144 28022 79762
rect 28190 79144 28206 79762
rect 28374 79144 28390 79762
rect 28558 79144 28574 79762
rect 28742 79144 28758 79762
rect 28926 79144 28942 79762
rect 29110 79144 29126 79762
rect 29294 79144 29310 79762
rect 29478 79144 29494 79762
rect 29662 79144 29678 79762
rect 29846 79144 29862 79762
rect 30030 79144 30046 79762
rect 30214 79144 30230 79762
rect 30398 79144 30414 79762
rect 30582 79144 30598 79762
rect 30766 79144 30782 79762
rect 30950 79144 30966 79762
rect 31134 79144 31150 79762
rect 31318 79144 31334 79762
rect 31502 79144 31518 79762
rect 31686 79144 31702 79762
rect 31870 79144 31886 79762
rect 32054 79144 32070 79762
rect 32238 79144 32254 79762
rect 32422 79144 32438 79762
rect 32606 79144 32622 79762
rect 32790 79144 32806 79762
rect 32974 79144 32990 79762
rect 33158 79144 33174 79762
rect 33342 79144 33358 79762
rect 33526 79144 33542 79762
rect 33710 79144 39982 79762
rect 40150 79144 40166 79762
rect 40334 79144 40350 79762
rect 40518 79144 40534 79762
rect 40702 79144 40718 79762
rect 40886 79144 40902 79762
rect 41070 79144 41086 79762
rect 41254 79144 41270 79762
rect 41438 79144 41454 79762
rect 41622 79144 41638 79762
rect 41806 79144 41822 79762
rect 41990 79144 42006 79762
rect 42174 79144 42190 79762
rect 42358 79144 42374 79762
rect 42542 79144 42558 79762
rect 42726 79144 42742 79762
rect 42910 79144 42926 79762
rect 43094 79144 43110 79762
rect 43278 79144 43294 79762
rect 43462 79144 43478 79762
rect 43646 79144 43662 79762
rect 43830 79144 43846 79762
rect 44014 79144 44030 79762
rect 44198 79144 44214 79762
rect 44382 79144 44398 79762
rect 44566 79144 44582 79762
rect 44750 79144 44766 79762
rect 44934 79144 44950 79762
rect 45118 79144 45134 79762
rect 45302 79144 45318 79762
rect 45486 79144 45502 79762
rect 45670 79144 45686 79762
rect 45854 79144 45870 79762
rect 46038 79144 46054 79762
rect 46222 79144 46238 79762
rect 46406 79144 46422 79762
rect 46590 79144 46606 79762
rect 46774 79144 46790 79762
rect 46958 79144 46974 79762
rect 47142 79144 47158 79762
rect 47326 79144 47342 79762
rect 47510 79144 47526 79762
rect 47694 79144 47710 79762
rect 47878 79144 47894 79762
rect 48062 79144 48078 79762
rect 48246 79144 48262 79762
rect 48430 79144 48446 79762
rect 48614 79144 48630 79762
rect 48798 79144 48814 79762
rect 48982 79144 48998 79762
rect 49166 79144 49182 79762
rect 49350 79144 49366 79762
rect 49534 79144 49550 79762
rect 49718 79144 49734 79762
rect 49902 79144 49918 79762
rect 50086 79144 50102 79762
rect 50270 79144 50286 79762
rect 50454 79144 50470 79762
rect 50638 79144 50654 79762
rect 50822 79144 50838 79762
rect 51006 79144 51022 79762
rect 51190 79144 51206 79762
rect 51374 79144 51390 79762
rect 51558 79144 51574 79762
rect 51742 79144 51758 79762
rect 51926 79144 51942 79762
rect 52110 79144 52126 79762
rect 52294 79144 52310 79762
rect 52478 79144 52494 79762
rect 52662 79144 52678 79762
rect 52846 79144 52862 79762
rect 53030 79144 53046 79762
rect 53214 79144 53230 79762
rect 53398 79144 53414 79762
rect 53582 79144 53598 79762
rect 53766 79144 53782 79762
rect 53950 79144 53966 79762
rect 54134 79144 54150 79762
rect 54318 79144 54334 79762
rect 54502 79144 54518 79762
rect 54686 79144 54702 79762
rect 54870 79144 54886 79762
rect 55054 79144 55070 79762
rect 55238 79144 55254 79762
rect 55422 79144 55438 79762
rect 55606 79144 55622 79762
rect 55790 79144 55806 79762
rect 55974 79144 55990 79762
rect 56158 79144 56174 79762
rect 56342 79144 56358 79762
rect 56526 79144 56542 79762
rect 56710 79144 56726 79762
rect 56894 79144 56910 79762
rect 57078 79144 57094 79762
rect 57262 79144 57278 79762
rect 57446 79144 57462 79762
rect 57630 79144 57646 79762
rect 57814 79144 57830 79762
rect 57998 79144 58014 79762
rect 58182 79144 58198 79762
rect 58366 79144 58382 79762
rect 58550 79144 58566 79762
rect 58734 79144 58750 79762
rect 58918 79144 58934 79762
rect 59102 79144 59118 79762
rect 59286 79144 65006 79762
rect 65174 79144 65190 79762
rect 65358 79144 65374 79762
rect 65542 79144 65558 79762
rect 65726 79144 65742 79762
rect 65910 79144 65926 79762
rect 66094 79144 66110 79762
rect 66278 79144 66294 79762
rect 66462 79144 66478 79762
rect 66646 79144 66662 79762
rect 66830 79144 66846 79762
rect 67014 79144 67030 79762
rect 67198 79144 67214 79762
rect 67382 79144 67398 79762
rect 67566 79144 67582 79762
rect 67750 79144 67766 79762
rect 67934 79144 67950 79762
rect 68118 79144 68134 79762
rect 68302 79144 68318 79762
rect 68486 79144 68502 79762
rect 68670 79144 68686 79762
rect 68854 79144 68870 79762
rect 69038 79144 69054 79762
rect 69222 79144 69238 79762
rect 69406 79144 69422 79762
rect 69590 79144 69606 79762
rect 69774 79144 69790 79762
rect 69958 79144 69974 79762
rect 70142 79144 70158 79762
rect 70326 79144 70342 79762
rect 70510 79144 70526 79762
rect 70694 79144 70710 79762
rect 70878 79144 70894 79762
rect 71062 79144 71078 79762
rect 71246 79144 71262 79762
rect 71430 79144 71446 79762
rect 71614 79144 71630 79762
rect 71798 79144 71814 79762
rect 71982 79144 71998 79762
rect 72166 79144 72182 79762
rect 72350 79144 72366 79762
rect 72534 79144 72550 79762
rect 72718 79144 72734 79762
rect 72902 79144 72918 79762
rect 73086 79144 73102 79762
rect 73270 79144 73286 79762
rect 73454 79144 73470 79762
rect 73638 79144 73654 79762
rect 73822 79144 73838 79762
rect 74006 79144 74022 79762
rect 74190 79144 74206 79762
rect 74374 79144 74390 79762
rect 74558 79144 74574 79762
rect 74742 79144 74758 79762
rect 74926 79144 74942 79762
rect 75110 79144 75126 79762
rect 75294 79144 75310 79762
rect 75478 79144 75494 79762
rect 75662 79144 75678 79762
rect 75846 79144 75862 79762
rect 76030 79144 76046 79762
rect 76214 79144 76230 79762
rect 76398 79144 76414 79762
rect 76582 79144 76598 79762
rect 76766 79144 76782 79762
rect 76950 79144 76966 79762
rect 77134 79144 77150 79762
rect 77318 79144 77334 79762
rect 77502 79144 77518 79762
rect 77686 79144 77702 79762
rect 77870 79144 77886 79762
rect 78054 79144 78070 79762
rect 78238 79144 78254 79762
rect 78422 79144 78438 79762
rect 78606 79144 78622 79762
rect 78790 79144 78806 79762
rect 78974 79144 78990 79762
rect 79158 79144 79174 79762
rect 79342 79144 79358 79762
rect 79526 79144 79542 79762
rect 79710 79144 79726 79762
rect 79894 79144 79910 79762
rect 80078 79144 80094 79762
rect 80262 79144 80278 79762
rect 80446 79144 89130 79762
rect 112 856 89130 79144
rect 222 70 238 856
rect 406 70 422 856
rect 590 70 606 856
rect 774 70 790 856
rect 958 70 974 856
rect 1142 70 1158 856
rect 1326 70 1342 856
rect 1510 70 1526 856
rect 1694 70 1710 856
rect 1878 70 1894 856
rect 2062 70 2078 856
rect 2246 70 2262 856
rect 2430 70 2446 856
rect 2614 70 2630 856
rect 2798 70 2814 856
rect 2982 70 2998 856
rect 3166 70 3182 856
rect 3350 70 3366 856
rect 3534 70 3550 856
rect 3718 70 3734 856
rect 3902 70 3918 856
rect 4086 70 4102 856
rect 4270 70 4286 856
rect 4454 70 4470 856
rect 4638 70 4654 856
rect 4822 70 4838 856
rect 5006 70 5022 856
rect 5190 70 5206 856
rect 5374 70 5390 856
rect 5558 70 5574 856
rect 5742 70 5758 856
rect 5926 70 5942 856
rect 6110 70 6126 856
rect 6294 70 6310 856
rect 6478 70 6494 856
rect 6662 70 6678 856
rect 6846 70 6862 856
rect 7030 70 7046 856
rect 7214 70 7230 856
rect 7398 70 7414 856
rect 7582 70 7598 856
rect 7766 70 7782 856
rect 7950 70 7966 856
rect 8134 70 8150 856
rect 8318 70 8334 856
rect 8502 70 8518 856
rect 8686 70 8702 856
rect 8870 70 8886 856
rect 9054 70 9070 856
rect 9238 70 9254 856
rect 9422 70 9438 856
rect 9606 70 9622 856
rect 9790 70 9806 856
rect 9974 70 9990 856
rect 10158 70 10174 856
rect 10342 70 10358 856
rect 10526 70 10542 856
rect 10710 70 10726 856
rect 10894 70 10910 856
rect 11078 70 11094 856
rect 11262 70 11278 856
rect 11446 70 11462 856
rect 11630 70 11646 856
rect 11814 70 11830 856
rect 11998 70 12014 856
rect 12182 70 12198 856
rect 12366 70 12382 856
rect 12550 70 12566 856
rect 12734 70 12750 856
rect 12918 70 12934 856
rect 13102 70 13118 856
rect 13286 70 13302 856
rect 13470 70 13486 856
rect 13654 70 13670 856
rect 13838 70 13854 856
rect 14022 70 14038 856
rect 14206 70 14222 856
rect 14390 70 14406 856
rect 14574 70 14590 856
rect 14758 70 14774 856
rect 14942 70 14958 856
rect 15126 70 15142 856
rect 15310 70 15326 856
rect 15494 70 15510 856
rect 15678 70 15694 856
rect 15862 70 15878 856
rect 16046 70 16062 856
rect 16230 70 16246 856
rect 16414 70 16430 856
rect 16598 70 16614 856
rect 16782 70 16798 856
rect 16966 70 16982 856
rect 17150 70 17166 856
rect 17334 70 17350 856
rect 17518 70 17534 856
rect 17702 70 17718 856
rect 17886 70 17902 856
rect 18070 70 18086 856
rect 18254 70 18270 856
rect 18438 70 18454 856
rect 18622 70 18638 856
rect 18806 70 18822 856
rect 18990 70 19006 856
rect 19174 70 19190 856
rect 19358 70 19374 856
rect 19542 70 19558 856
rect 19726 70 19742 856
rect 19910 70 19926 856
rect 20094 70 50010 856
rect 50178 70 50194 856
rect 50362 70 50378 856
rect 50546 70 50562 856
rect 50730 70 50746 856
rect 50914 70 50930 856
rect 51098 70 51114 856
rect 51282 70 51298 856
rect 51466 70 51482 856
rect 51650 70 51666 856
rect 51834 70 51850 856
rect 52018 70 52034 856
rect 52202 70 52218 856
rect 52386 70 52402 856
rect 52570 70 52586 856
rect 52754 70 52770 856
rect 52938 70 52954 856
rect 53122 70 53138 856
rect 53306 70 89130 856
<< metal3 >>
rect 89200 61752 90800 61872
rect 89200 61480 90800 61600
rect 89200 61208 90800 61328
rect 89200 60936 90800 61056
rect 89200 60664 90800 60784
rect 89200 60392 90800 60512
rect 89200 60120 90800 60240
rect 89200 416 90800 536
rect 89200 144 90800 264
<< obsm3 >>
rect 289 61952 89200 78845
rect 289 60040 89120 61952
rect 289 616 89200 60040
rect 289 171 89120 616
<< metal4 >>
rect 3748 2128 4988 77840
rect 13748 2128 14988 77840
rect 23748 2128 24988 77840
rect 33748 2128 34988 77840
rect 43748 2128 44988 77840
rect 53748 2128 54988 77840
rect 63748 2128 64988 77840
rect 73748 2128 74988 77840
rect 83748 2128 84988 77840
<< obsm4 >>
rect 5211 77920 85317 78845
rect 5211 2483 13668 77920
rect 15068 2483 23668 77920
rect 25068 2483 33668 77920
rect 35068 2483 43668 77920
rect 45068 2483 53668 77920
rect 55068 2483 63668 77920
rect 65068 2483 73668 77920
rect 75068 2483 83668 77920
rect 85068 2483 85317 77920
<< labels >>
rlabel metal2 s 32862 79200 32918 80800 6 cfg_clk_skew_ctrl1[0]
port 1 nsew signal output
rlabel metal2 s 31758 79200 31814 80800 6 cfg_clk_skew_ctrl1[10]
port 2 nsew signal output
rlabel metal2 s 31574 79200 31630 80800 6 cfg_clk_skew_ctrl1[11]
port 3 nsew signal output
rlabel metal2 s 31390 79200 31446 80800 6 cfg_clk_skew_ctrl1[12]
port 4 nsew signal output
rlabel metal2 s 31206 79200 31262 80800 6 cfg_clk_skew_ctrl1[13]
port 5 nsew signal output
rlabel metal2 s 31022 79200 31078 80800 6 cfg_clk_skew_ctrl1[14]
port 6 nsew signal output
rlabel metal2 s 30838 79200 30894 80800 6 cfg_clk_skew_ctrl1[15]
port 7 nsew signal output
rlabel metal2 s 30654 79200 30710 80800 6 cfg_clk_skew_ctrl1[16]
port 8 nsew signal output
rlabel metal2 s 30470 79200 30526 80800 6 cfg_clk_skew_ctrl1[17]
port 9 nsew signal output
rlabel metal2 s 30286 79200 30342 80800 6 cfg_clk_skew_ctrl1[18]
port 10 nsew signal output
rlabel metal2 s 30102 79200 30158 80800 6 cfg_clk_skew_ctrl1[19]
port 11 nsew signal output
rlabel metal2 s 32678 79200 32734 80800 6 cfg_clk_skew_ctrl1[1]
port 12 nsew signal output
rlabel metal2 s 29918 79200 29974 80800 6 cfg_clk_skew_ctrl1[20]
port 13 nsew signal output
rlabel metal2 s 29734 79200 29790 80800 6 cfg_clk_skew_ctrl1[21]
port 14 nsew signal output
rlabel metal2 s 29550 79200 29606 80800 6 cfg_clk_skew_ctrl1[22]
port 15 nsew signal output
rlabel metal2 s 29366 79200 29422 80800 6 cfg_clk_skew_ctrl1[23]
port 16 nsew signal output
rlabel metal2 s 29182 79200 29238 80800 6 cfg_clk_skew_ctrl1[24]
port 17 nsew signal output
rlabel metal2 s 28998 79200 29054 80800 6 cfg_clk_skew_ctrl1[25]
port 18 nsew signal output
rlabel metal2 s 28814 79200 28870 80800 6 cfg_clk_skew_ctrl1[26]
port 19 nsew signal output
rlabel metal2 s 28630 79200 28686 80800 6 cfg_clk_skew_ctrl1[27]
port 20 nsew signal output
rlabel metal2 s 65614 79200 65670 80800 6 cfg_clk_skew_ctrl1[28]
port 21 nsew signal output
rlabel metal2 s 65430 79200 65486 80800 6 cfg_clk_skew_ctrl1[29]
port 22 nsew signal output
rlabel metal2 s 32494 79200 32550 80800 6 cfg_clk_skew_ctrl1[2]
port 23 nsew signal output
rlabel metal2 s 65246 79200 65302 80800 6 cfg_clk_skew_ctrl1[30]
port 24 nsew signal output
rlabel metal2 s 65062 79200 65118 80800 6 cfg_clk_skew_ctrl1[31]
port 25 nsew signal output
rlabel metal2 s 32310 79200 32366 80800 6 cfg_clk_skew_ctrl1[3]
port 26 nsew signal output
rlabel metal2 s 1214 79200 1270 80800 6 cfg_clk_skew_ctrl1[4]
port 27 nsew signal output
rlabel metal2 s 846 79200 902 80800 6 cfg_clk_skew_ctrl1[5]
port 28 nsew signal output
rlabel metal2 s 478 79200 534 80800 6 cfg_clk_skew_ctrl1[6]
port 29 nsew signal output
rlabel metal2 s 110 79200 166 80800 6 cfg_clk_skew_ctrl1[7]
port 30 nsew signal output
rlabel metal2 s 32126 79200 32182 80800 6 cfg_clk_skew_ctrl1[8]
port 31 nsew signal output
rlabel metal2 s 31942 79200 31998 80800 6 cfg_clk_skew_ctrl1[9]
port 32 nsew signal output
rlabel metal2 s 28446 79200 28502 80800 6 cfg_clk_skew_ctrl2[0]
port 33 nsew signal output
rlabel metal2 s 26606 79200 26662 80800 6 cfg_clk_skew_ctrl2[10]
port 34 nsew signal output
rlabel metal2 s 26422 79200 26478 80800 6 cfg_clk_skew_ctrl2[11]
port 35 nsew signal output
rlabel metal2 s 26238 79200 26294 80800 6 cfg_clk_skew_ctrl2[12]
port 36 nsew signal output
rlabel metal2 s 26054 79200 26110 80800 6 cfg_clk_skew_ctrl2[13]
port 37 nsew signal output
rlabel metal2 s 25870 79200 25926 80800 6 cfg_clk_skew_ctrl2[14]
port 38 nsew signal output
rlabel metal2 s 25686 79200 25742 80800 6 cfg_clk_skew_ctrl2[15]
port 39 nsew signal output
rlabel metal2 s 25502 79200 25558 80800 6 cfg_clk_skew_ctrl2[16]
port 40 nsew signal output
rlabel metal2 s 25318 79200 25374 80800 6 cfg_clk_skew_ctrl2[17]
port 41 nsew signal output
rlabel metal2 s 25134 79200 25190 80800 6 cfg_clk_skew_ctrl2[18]
port 42 nsew signal output
rlabel metal2 s 24950 79200 25006 80800 6 cfg_clk_skew_ctrl2[19]
port 43 nsew signal output
rlabel metal2 s 28262 79200 28318 80800 6 cfg_clk_skew_ctrl2[1]
port 44 nsew signal output
rlabel metal2 s 24766 79200 24822 80800 6 cfg_clk_skew_ctrl2[20]
port 45 nsew signal output
rlabel metal2 s 24582 79200 24638 80800 6 cfg_clk_skew_ctrl2[21]
port 46 nsew signal output
rlabel metal2 s 24398 79200 24454 80800 6 cfg_clk_skew_ctrl2[22]
port 47 nsew signal output
rlabel metal2 s 24214 79200 24270 80800 6 cfg_clk_skew_ctrl2[23]
port 48 nsew signal output
rlabel metal2 s 67086 79200 67142 80800 6 cfg_clk_skew_ctrl2[24]
port 49 nsew signal output
rlabel metal2 s 66902 79200 66958 80800 6 cfg_clk_skew_ctrl2[25]
port 50 nsew signal output
rlabel metal2 s 66718 79200 66774 80800 6 cfg_clk_skew_ctrl2[26]
port 51 nsew signal output
rlabel metal2 s 66534 79200 66590 80800 6 cfg_clk_skew_ctrl2[27]
port 52 nsew signal output
rlabel metal2 s 66350 79200 66406 80800 6 cfg_clk_skew_ctrl2[28]
port 53 nsew signal output
rlabel metal2 s 66166 79200 66222 80800 6 cfg_clk_skew_ctrl2[29]
port 54 nsew signal output
rlabel metal2 s 28078 79200 28134 80800 6 cfg_clk_skew_ctrl2[2]
port 55 nsew signal output
rlabel metal2 s 65982 79200 66038 80800 6 cfg_clk_skew_ctrl2[30]
port 56 nsew signal output
rlabel metal2 s 65798 79200 65854 80800 6 cfg_clk_skew_ctrl2[31]
port 57 nsew signal output
rlabel metal2 s 27894 79200 27950 80800 6 cfg_clk_skew_ctrl2[3]
port 58 nsew signal output
rlabel metal2 s 27710 79200 27766 80800 6 cfg_clk_skew_ctrl2[4]
port 59 nsew signal output
rlabel metal2 s 27526 79200 27582 80800 6 cfg_clk_skew_ctrl2[5]
port 60 nsew signal output
rlabel metal2 s 27342 79200 27398 80800 6 cfg_clk_skew_ctrl2[6]
port 61 nsew signal output
rlabel metal2 s 27158 79200 27214 80800 6 cfg_clk_skew_ctrl2[7]
port 62 nsew signal output
rlabel metal2 s 26974 79200 27030 80800 6 cfg_clk_skew_ctrl2[8]
port 63 nsew signal output
rlabel metal2 s 26790 79200 26846 80800 6 cfg_clk_skew_ctrl2[9]
port 64 nsew signal output
rlabel metal2 s 1398 79200 1454 80800 6 cfg_cska_wh[0]
port 65 nsew signal input
rlabel metal2 s 1030 79200 1086 80800 6 cfg_cska_wh[1]
port 66 nsew signal input
rlabel metal2 s 662 79200 718 80800 6 cfg_cska_wh[2]
port 67 nsew signal input
rlabel metal2 s 294 79200 350 80800 6 cfg_cska_wh[3]
port 68 nsew signal input
rlabel metal3 s 89200 416 90800 536 6 cfg_fast_sim
port 69 nsew signal output
rlabel metal2 s 79414 79200 79470 80800 6 cfg_strap_pad_ctrl
port 70 nsew signal output
rlabel metal2 s 20074 79200 20130 80800 6 cpu_clk
port 71 nsew signal output
rlabel metal2 s 79598 79200 79654 80800 6 e_reset_n
port 72 nsew signal output
rlabel metal2 s 79966 79200 80022 80800 6 int_pll_clock
port 73 nsew signal input
rlabel metal2 s 50066 -800 50122 800 8 la_data_in[0]
port 74 nsew signal input
rlabel metal2 s 51906 -800 51962 800 8 la_data_in[10]
port 75 nsew signal input
rlabel metal2 s 52090 -800 52146 800 8 la_data_in[11]
port 76 nsew signal input
rlabel metal2 s 52274 -800 52330 800 8 la_data_in[12]
port 77 nsew signal input
rlabel metal2 s 52458 -800 52514 800 8 la_data_in[13]
port 78 nsew signal input
rlabel metal2 s 52642 -800 52698 800 8 la_data_in[14]
port 79 nsew signal input
rlabel metal2 s 52826 -800 52882 800 8 la_data_in[15]
port 80 nsew signal input
rlabel metal2 s 53010 -800 53066 800 8 la_data_in[16]
port 81 nsew signal input
rlabel metal2 s 53194 -800 53250 800 8 la_data_in[17]
port 82 nsew signal input
rlabel metal2 s 50250 -800 50306 800 8 la_data_in[1]
port 83 nsew signal input
rlabel metal2 s 50434 -800 50490 800 8 la_data_in[2]
port 84 nsew signal input
rlabel metal2 s 50618 -800 50674 800 8 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 50802 -800 50858 800 8 la_data_in[4]
port 86 nsew signal input
rlabel metal2 s 50986 -800 51042 800 8 la_data_in[5]
port 87 nsew signal input
rlabel metal2 s 51170 -800 51226 800 8 la_data_in[6]
port 88 nsew signal input
rlabel metal2 s 51354 -800 51410 800 8 la_data_in[7]
port 89 nsew signal input
rlabel metal2 s 51538 -800 51594 800 8 la_data_in[8]
port 90 nsew signal input
rlabel metal2 s 51722 -800 51778 800 8 la_data_in[9]
port 91 nsew signal input
rlabel metal2 s 79782 79200 79838 80800 6 p_reset_n
port 92 nsew signal output
rlabel metal2 s 80334 79200 80390 80800 6 s_reset_n
port 93 nsew signal output
rlabel metal3 s 89200 60664 90800 60784 6 sclk
port 94 nsew signal input
rlabel metal3 s 89200 61208 90800 61328 6 sdin
port 95 nsew signal input
rlabel metal3 s 89200 61480 90800 61600 6 sdout
port 96 nsew signal output
rlabel metal3 s 89200 61752 90800 61872 6 sdout_oen
port 97 nsew signal output
rlabel metal3 s 89200 60936 90800 61056 6 ssn
port 98 nsew signal input
rlabel metal2 s 72974 79200 73030 80800 6 strap_sticky[0]
port 99 nsew signal input
rlabel metal2 s 71134 79200 71190 80800 6 strap_sticky[10]
port 100 nsew signal input
rlabel metal2 s 70950 79200 71006 80800 6 strap_sticky[11]
port 101 nsew signal input
rlabel metal2 s 70766 79200 70822 80800 6 strap_sticky[12]
port 102 nsew signal input
rlabel metal2 s 70582 79200 70638 80800 6 strap_sticky[13]
port 103 nsew signal input
rlabel metal2 s 70398 79200 70454 80800 6 strap_sticky[14]
port 104 nsew signal input
rlabel metal2 s 70214 79200 70270 80800 6 strap_sticky[15]
port 105 nsew signal input
rlabel metal2 s 70030 79200 70086 80800 6 strap_sticky[16]
port 106 nsew signal input
rlabel metal2 s 69846 79200 69902 80800 6 strap_sticky[17]
port 107 nsew signal input
rlabel metal2 s 69662 79200 69718 80800 6 strap_sticky[18]
port 108 nsew signal input
rlabel metal2 s 69478 79200 69534 80800 6 strap_sticky[19]
port 109 nsew signal input
rlabel metal2 s 72790 79200 72846 80800 6 strap_sticky[1]
port 110 nsew signal input
rlabel metal2 s 69294 79200 69350 80800 6 strap_sticky[20]
port 111 nsew signal input
rlabel metal2 s 69110 79200 69166 80800 6 strap_sticky[21]
port 112 nsew signal input
rlabel metal2 s 68926 79200 68982 80800 6 strap_sticky[22]
port 113 nsew signal input
rlabel metal2 s 68742 79200 68798 80800 6 strap_sticky[23]
port 114 nsew signal input
rlabel metal2 s 68558 79200 68614 80800 6 strap_sticky[24]
port 115 nsew signal input
rlabel metal2 s 68374 79200 68430 80800 6 strap_sticky[25]
port 116 nsew signal input
rlabel metal2 s 68190 79200 68246 80800 6 strap_sticky[26]
port 117 nsew signal input
rlabel metal2 s 68006 79200 68062 80800 6 strap_sticky[27]
port 118 nsew signal input
rlabel metal2 s 67822 79200 67878 80800 6 strap_sticky[28]
port 119 nsew signal input
rlabel metal2 s 67638 79200 67694 80800 6 strap_sticky[29]
port 120 nsew signal input
rlabel metal2 s 72606 79200 72662 80800 6 strap_sticky[2]
port 121 nsew signal input
rlabel metal2 s 67454 79200 67510 80800 6 strap_sticky[30]
port 122 nsew signal input
rlabel metal2 s 67270 79200 67326 80800 6 strap_sticky[31]
port 123 nsew signal input
rlabel metal2 s 72422 79200 72478 80800 6 strap_sticky[3]
port 124 nsew signal input
rlabel metal2 s 72238 79200 72294 80800 6 strap_sticky[4]
port 125 nsew signal input
rlabel metal2 s 72054 79200 72110 80800 6 strap_sticky[5]
port 126 nsew signal input
rlabel metal2 s 71870 79200 71926 80800 6 strap_sticky[6]
port 127 nsew signal input
rlabel metal2 s 71686 79200 71742 80800 6 strap_sticky[7]
port 128 nsew signal input
rlabel metal2 s 71502 79200 71558 80800 6 strap_sticky[8]
port 129 nsew signal input
rlabel metal2 s 71318 79200 71374 80800 6 strap_sticky[9]
port 130 nsew signal input
rlabel metal2 s 73342 79200 73398 80800 6 strap_uartm[0]
port 131 nsew signal input
rlabel metal2 s 73158 79200 73214 80800 6 strap_uartm[1]
port 132 nsew signal input
rlabel metal2 s 79230 79200 79286 80800 6 system_strap[0]
port 133 nsew signal output
rlabel metal2 s 77390 79200 77446 80800 6 system_strap[10]
port 134 nsew signal output
rlabel metal2 s 77206 79200 77262 80800 6 system_strap[11]
port 135 nsew signal output
rlabel metal2 s 77022 79200 77078 80800 6 system_strap[12]
port 136 nsew signal output
rlabel metal2 s 76838 79200 76894 80800 6 system_strap[13]
port 137 nsew signal output
rlabel metal2 s 76654 79200 76710 80800 6 system_strap[14]
port 138 nsew signal output
rlabel metal2 s 76470 79200 76526 80800 6 system_strap[15]
port 139 nsew signal output
rlabel metal2 s 76286 79200 76342 80800 6 system_strap[16]
port 140 nsew signal output
rlabel metal2 s 76102 79200 76158 80800 6 system_strap[17]
port 141 nsew signal output
rlabel metal2 s 75918 79200 75974 80800 6 system_strap[18]
port 142 nsew signal output
rlabel metal2 s 75734 79200 75790 80800 6 system_strap[19]
port 143 nsew signal output
rlabel metal2 s 79046 79200 79102 80800 6 system_strap[1]
port 144 nsew signal output
rlabel metal2 s 75550 79200 75606 80800 6 system_strap[20]
port 145 nsew signal output
rlabel metal2 s 75366 79200 75422 80800 6 system_strap[21]
port 146 nsew signal output
rlabel metal2 s 75182 79200 75238 80800 6 system_strap[22]
port 147 nsew signal output
rlabel metal2 s 74998 79200 75054 80800 6 system_strap[23]
port 148 nsew signal output
rlabel metal2 s 74814 79200 74870 80800 6 system_strap[24]
port 149 nsew signal output
rlabel metal2 s 74630 79200 74686 80800 6 system_strap[25]
port 150 nsew signal output
rlabel metal2 s 74446 79200 74502 80800 6 system_strap[26]
port 151 nsew signal output
rlabel metal2 s 74262 79200 74318 80800 6 system_strap[27]
port 152 nsew signal output
rlabel metal2 s 74078 79200 74134 80800 6 system_strap[28]
port 153 nsew signal output
rlabel metal2 s 73894 79200 73950 80800 6 system_strap[29]
port 154 nsew signal output
rlabel metal2 s 78862 79200 78918 80800 6 system_strap[2]
port 155 nsew signal output
rlabel metal2 s 73710 79200 73766 80800 6 system_strap[30]
port 156 nsew signal output
rlabel metal2 s 73526 79200 73582 80800 6 system_strap[31]
port 157 nsew signal output
rlabel metal2 s 78678 79200 78734 80800 6 system_strap[3]
port 158 nsew signal output
rlabel metal2 s 78494 79200 78550 80800 6 system_strap[4]
port 159 nsew signal output
rlabel metal2 s 78310 79200 78366 80800 6 system_strap[5]
port 160 nsew signal output
rlabel metal2 s 78126 79200 78182 80800 6 system_strap[6]
port 161 nsew signal output
rlabel metal2 s 77942 79200 77998 80800 6 system_strap[7]
port 162 nsew signal output
rlabel metal2 s 77758 79200 77814 80800 6 system_strap[8]
port 163 nsew signal output
rlabel metal2 s 77574 79200 77630 80800 6 system_strap[9]
port 164 nsew signal output
rlabel metal3 s 89200 60120 90800 60240 6 uartm_rxd
port 165 nsew signal input
rlabel metal3 s 89200 60392 90800 60512 6 uartm_txd
port 166 nsew signal output
rlabel metal2 s 294 -800 350 800 8 user_clock1
port 167 nsew signal input
rlabel metal2 s 110 -800 166 800 8 user_clock2
port 168 nsew signal input
rlabel metal4 s 3748 2128 4988 77840 6 vccd1
port 169 nsew power bidirectional
rlabel metal4 s 23748 2128 24988 77840 6 vccd1
port 169 nsew power bidirectional
rlabel metal4 s 43748 2128 44988 77840 6 vccd1
port 169 nsew power bidirectional
rlabel metal4 s 63748 2128 64988 77840 6 vccd1
port 169 nsew power bidirectional
rlabel metal4 s 83748 2128 84988 77840 6 vccd1
port 169 nsew power bidirectional
rlabel metal4 s 13748 2128 14988 77840 6 vssd1
port 170 nsew ground bidirectional
rlabel metal4 s 33748 2128 34988 77840 6 vssd1
port 170 nsew ground bidirectional
rlabel metal4 s 53748 2128 54988 77840 6 vssd1
port 170 nsew ground bidirectional
rlabel metal4 s 73748 2128 74988 77840 6 vssd1
port 170 nsew ground bidirectional
rlabel metal2 s 33046 79200 33102 80800 6 wbd_clk_int
port 171 nsew signal input
rlabel metal2 s 33598 79200 33654 80800 6 wbd_clk_wh
port 172 nsew signal output
rlabel metal2 s 24030 79200 24086 80800 6 wbd_int_rst_n
port 173 nsew signal output
rlabel metal3 s 89200 144 90800 264 6 wbd_pll_rst_n
port 174 nsew signal output
rlabel metal2 s 846 -800 902 800 8 wbm_ack_o
port 175 nsew signal output
rlabel metal2 s 1582 -800 1638 800 8 wbm_adr_i[0]
port 176 nsew signal input
rlabel metal2 s 7838 -800 7894 800 8 wbm_adr_i[10]
port 177 nsew signal input
rlabel metal2 s 8390 -800 8446 800 8 wbm_adr_i[11]
port 178 nsew signal input
rlabel metal2 s 8942 -800 8998 800 8 wbm_adr_i[12]
port 179 nsew signal input
rlabel metal2 s 9494 -800 9550 800 8 wbm_adr_i[13]
port 180 nsew signal input
rlabel metal2 s 10046 -800 10102 800 8 wbm_adr_i[14]
port 181 nsew signal input
rlabel metal2 s 10598 -800 10654 800 8 wbm_adr_i[15]
port 182 nsew signal input
rlabel metal2 s 11150 -800 11206 800 8 wbm_adr_i[16]
port 183 nsew signal input
rlabel metal2 s 11702 -800 11758 800 8 wbm_adr_i[17]
port 184 nsew signal input
rlabel metal2 s 12254 -800 12310 800 8 wbm_adr_i[18]
port 185 nsew signal input
rlabel metal2 s 12806 -800 12862 800 8 wbm_adr_i[19]
port 186 nsew signal input
rlabel metal2 s 2318 -800 2374 800 8 wbm_adr_i[1]
port 187 nsew signal input
rlabel metal2 s 13358 -800 13414 800 8 wbm_adr_i[20]
port 188 nsew signal input
rlabel metal2 s 13910 -800 13966 800 8 wbm_adr_i[21]
port 189 nsew signal input
rlabel metal2 s 14462 -800 14518 800 8 wbm_adr_i[22]
port 190 nsew signal input
rlabel metal2 s 15014 -800 15070 800 8 wbm_adr_i[23]
port 191 nsew signal input
rlabel metal2 s 15566 -800 15622 800 8 wbm_adr_i[24]
port 192 nsew signal input
rlabel metal2 s 16118 -800 16174 800 8 wbm_adr_i[25]
port 193 nsew signal input
rlabel metal2 s 16670 -800 16726 800 8 wbm_adr_i[26]
port 194 nsew signal input
rlabel metal2 s 17222 -800 17278 800 8 wbm_adr_i[27]
port 195 nsew signal input
rlabel metal2 s 17774 -800 17830 800 8 wbm_adr_i[28]
port 196 nsew signal input
rlabel metal2 s 18326 -800 18382 800 8 wbm_adr_i[29]
port 197 nsew signal input
rlabel metal2 s 3054 -800 3110 800 8 wbm_adr_i[2]
port 198 nsew signal input
rlabel metal2 s 18878 -800 18934 800 8 wbm_adr_i[30]
port 199 nsew signal input
rlabel metal2 s 19430 -800 19486 800 8 wbm_adr_i[31]
port 200 nsew signal input
rlabel metal2 s 3790 -800 3846 800 8 wbm_adr_i[3]
port 201 nsew signal input
rlabel metal2 s 4526 -800 4582 800 8 wbm_adr_i[4]
port 202 nsew signal input
rlabel metal2 s 5078 -800 5134 800 8 wbm_adr_i[5]
port 203 nsew signal input
rlabel metal2 s 5630 -800 5686 800 8 wbm_adr_i[6]
port 204 nsew signal input
rlabel metal2 s 6182 -800 6238 800 8 wbm_adr_i[7]
port 205 nsew signal input
rlabel metal2 s 6734 -800 6790 800 8 wbm_adr_i[8]
port 206 nsew signal input
rlabel metal2 s 7286 -800 7342 800 8 wbm_adr_i[9]
port 207 nsew signal input
rlabel metal2 s 478 -800 534 800 8 wbm_clk_i
port 208 nsew signal input
rlabel metal2 s 1030 -800 1086 800 8 wbm_cyc_i
port 209 nsew signal input
rlabel metal2 s 1766 -800 1822 800 8 wbm_dat_i[0]
port 210 nsew signal input
rlabel metal2 s 8022 -800 8078 800 8 wbm_dat_i[10]
port 211 nsew signal input
rlabel metal2 s 8574 -800 8630 800 8 wbm_dat_i[11]
port 212 nsew signal input
rlabel metal2 s 9126 -800 9182 800 8 wbm_dat_i[12]
port 213 nsew signal input
rlabel metal2 s 9678 -800 9734 800 8 wbm_dat_i[13]
port 214 nsew signal input
rlabel metal2 s 10230 -800 10286 800 8 wbm_dat_i[14]
port 215 nsew signal input
rlabel metal2 s 10782 -800 10838 800 8 wbm_dat_i[15]
port 216 nsew signal input
rlabel metal2 s 11334 -800 11390 800 8 wbm_dat_i[16]
port 217 nsew signal input
rlabel metal2 s 11886 -800 11942 800 8 wbm_dat_i[17]
port 218 nsew signal input
rlabel metal2 s 12438 -800 12494 800 8 wbm_dat_i[18]
port 219 nsew signal input
rlabel metal2 s 12990 -800 13046 800 8 wbm_dat_i[19]
port 220 nsew signal input
rlabel metal2 s 2502 -800 2558 800 8 wbm_dat_i[1]
port 221 nsew signal input
rlabel metal2 s 13542 -800 13598 800 8 wbm_dat_i[20]
port 222 nsew signal input
rlabel metal2 s 14094 -800 14150 800 8 wbm_dat_i[21]
port 223 nsew signal input
rlabel metal2 s 14646 -800 14702 800 8 wbm_dat_i[22]
port 224 nsew signal input
rlabel metal2 s 15198 -800 15254 800 8 wbm_dat_i[23]
port 225 nsew signal input
rlabel metal2 s 15750 -800 15806 800 8 wbm_dat_i[24]
port 226 nsew signal input
rlabel metal2 s 16302 -800 16358 800 8 wbm_dat_i[25]
port 227 nsew signal input
rlabel metal2 s 16854 -800 16910 800 8 wbm_dat_i[26]
port 228 nsew signal input
rlabel metal2 s 17406 -800 17462 800 8 wbm_dat_i[27]
port 229 nsew signal input
rlabel metal2 s 17958 -800 18014 800 8 wbm_dat_i[28]
port 230 nsew signal input
rlabel metal2 s 18510 -800 18566 800 8 wbm_dat_i[29]
port 231 nsew signal input
rlabel metal2 s 3238 -800 3294 800 8 wbm_dat_i[2]
port 232 nsew signal input
rlabel metal2 s 19062 -800 19118 800 8 wbm_dat_i[30]
port 233 nsew signal input
rlabel metal2 s 19614 -800 19670 800 8 wbm_dat_i[31]
port 234 nsew signal input
rlabel metal2 s 3974 -800 4030 800 8 wbm_dat_i[3]
port 235 nsew signal input
rlabel metal2 s 4710 -800 4766 800 8 wbm_dat_i[4]
port 236 nsew signal input
rlabel metal2 s 5262 -800 5318 800 8 wbm_dat_i[5]
port 237 nsew signal input
rlabel metal2 s 5814 -800 5870 800 8 wbm_dat_i[6]
port 238 nsew signal input
rlabel metal2 s 6366 -800 6422 800 8 wbm_dat_i[7]
port 239 nsew signal input
rlabel metal2 s 6918 -800 6974 800 8 wbm_dat_i[8]
port 240 nsew signal input
rlabel metal2 s 7470 -800 7526 800 8 wbm_dat_i[9]
port 241 nsew signal input
rlabel metal2 s 1950 -800 2006 800 8 wbm_dat_o[0]
port 242 nsew signal output
rlabel metal2 s 8206 -800 8262 800 8 wbm_dat_o[10]
port 243 nsew signal output
rlabel metal2 s 8758 -800 8814 800 8 wbm_dat_o[11]
port 244 nsew signal output
rlabel metal2 s 9310 -800 9366 800 8 wbm_dat_o[12]
port 245 nsew signal output
rlabel metal2 s 9862 -800 9918 800 8 wbm_dat_o[13]
port 246 nsew signal output
rlabel metal2 s 10414 -800 10470 800 8 wbm_dat_o[14]
port 247 nsew signal output
rlabel metal2 s 10966 -800 11022 800 8 wbm_dat_o[15]
port 248 nsew signal output
rlabel metal2 s 11518 -800 11574 800 8 wbm_dat_o[16]
port 249 nsew signal output
rlabel metal2 s 12070 -800 12126 800 8 wbm_dat_o[17]
port 250 nsew signal output
rlabel metal2 s 12622 -800 12678 800 8 wbm_dat_o[18]
port 251 nsew signal output
rlabel metal2 s 13174 -800 13230 800 8 wbm_dat_o[19]
port 252 nsew signal output
rlabel metal2 s 2686 -800 2742 800 8 wbm_dat_o[1]
port 253 nsew signal output
rlabel metal2 s 13726 -800 13782 800 8 wbm_dat_o[20]
port 254 nsew signal output
rlabel metal2 s 14278 -800 14334 800 8 wbm_dat_o[21]
port 255 nsew signal output
rlabel metal2 s 14830 -800 14886 800 8 wbm_dat_o[22]
port 256 nsew signal output
rlabel metal2 s 15382 -800 15438 800 8 wbm_dat_o[23]
port 257 nsew signal output
rlabel metal2 s 15934 -800 15990 800 8 wbm_dat_o[24]
port 258 nsew signal output
rlabel metal2 s 16486 -800 16542 800 8 wbm_dat_o[25]
port 259 nsew signal output
rlabel metal2 s 17038 -800 17094 800 8 wbm_dat_o[26]
port 260 nsew signal output
rlabel metal2 s 17590 -800 17646 800 8 wbm_dat_o[27]
port 261 nsew signal output
rlabel metal2 s 18142 -800 18198 800 8 wbm_dat_o[28]
port 262 nsew signal output
rlabel metal2 s 18694 -800 18750 800 8 wbm_dat_o[29]
port 263 nsew signal output
rlabel metal2 s 3422 -800 3478 800 8 wbm_dat_o[2]
port 264 nsew signal output
rlabel metal2 s 19246 -800 19302 800 8 wbm_dat_o[30]
port 265 nsew signal output
rlabel metal2 s 19798 -800 19854 800 8 wbm_dat_o[31]
port 266 nsew signal output
rlabel metal2 s 4158 -800 4214 800 8 wbm_dat_o[3]
port 267 nsew signal output
rlabel metal2 s 4894 -800 4950 800 8 wbm_dat_o[4]
port 268 nsew signal output
rlabel metal2 s 5446 -800 5502 800 8 wbm_dat_o[5]
port 269 nsew signal output
rlabel metal2 s 5998 -800 6054 800 8 wbm_dat_o[6]
port 270 nsew signal output
rlabel metal2 s 6550 -800 6606 800 8 wbm_dat_o[7]
port 271 nsew signal output
rlabel metal2 s 7102 -800 7158 800 8 wbm_dat_o[8]
port 272 nsew signal output
rlabel metal2 s 7654 -800 7710 800 8 wbm_dat_o[9]
port 273 nsew signal output
rlabel metal2 s 19982 -800 20038 800 8 wbm_err_o
port 274 nsew signal output
rlabel metal2 s 662 -800 718 800 8 wbm_rst_i
port 275 nsew signal input
rlabel metal2 s 2134 -800 2190 800 8 wbm_sel_i[0]
port 276 nsew signal input
rlabel metal2 s 2870 -800 2926 800 8 wbm_sel_i[1]
port 277 nsew signal input
rlabel metal2 s 3606 -800 3662 800 8 wbm_sel_i[2]
port 278 nsew signal input
rlabel metal2 s 4342 -800 4398 800 8 wbm_sel_i[3]
port 279 nsew signal input
rlabel metal2 s 1214 -800 1270 800 8 wbm_stb_i
port 280 nsew signal input
rlabel metal2 s 1398 -800 1454 800 8 wbm_we_i
port 281 nsew signal input
rlabel metal2 s 58806 79200 58862 80800 6 wbs_ack_i
port 282 nsew signal input
rlabel metal2 s 46110 79200 46166 80800 6 wbs_adr_o[0]
port 283 nsew signal output
rlabel metal2 s 44270 79200 44326 80800 6 wbs_adr_o[10]
port 284 nsew signal output
rlabel metal2 s 44086 79200 44142 80800 6 wbs_adr_o[11]
port 285 nsew signal output
rlabel metal2 s 43902 79200 43958 80800 6 wbs_adr_o[12]
port 286 nsew signal output
rlabel metal2 s 43718 79200 43774 80800 6 wbs_adr_o[13]
port 287 nsew signal output
rlabel metal2 s 43534 79200 43590 80800 6 wbs_adr_o[14]
port 288 nsew signal output
rlabel metal2 s 43350 79200 43406 80800 6 wbs_adr_o[15]
port 289 nsew signal output
rlabel metal2 s 43166 79200 43222 80800 6 wbs_adr_o[16]
port 290 nsew signal output
rlabel metal2 s 42982 79200 43038 80800 6 wbs_adr_o[17]
port 291 nsew signal output
rlabel metal2 s 42798 79200 42854 80800 6 wbs_adr_o[18]
port 292 nsew signal output
rlabel metal2 s 42614 79200 42670 80800 6 wbs_adr_o[19]
port 293 nsew signal output
rlabel metal2 s 45926 79200 45982 80800 6 wbs_adr_o[1]
port 294 nsew signal output
rlabel metal2 s 42430 79200 42486 80800 6 wbs_adr_o[20]
port 295 nsew signal output
rlabel metal2 s 42246 79200 42302 80800 6 wbs_adr_o[21]
port 296 nsew signal output
rlabel metal2 s 42062 79200 42118 80800 6 wbs_adr_o[22]
port 297 nsew signal output
rlabel metal2 s 41878 79200 41934 80800 6 wbs_adr_o[23]
port 298 nsew signal output
rlabel metal2 s 41694 79200 41750 80800 6 wbs_adr_o[24]
port 299 nsew signal output
rlabel metal2 s 41510 79200 41566 80800 6 wbs_adr_o[25]
port 300 nsew signal output
rlabel metal2 s 41326 79200 41382 80800 6 wbs_adr_o[26]
port 301 nsew signal output
rlabel metal2 s 41142 79200 41198 80800 6 wbs_adr_o[27]
port 302 nsew signal output
rlabel metal2 s 40958 79200 41014 80800 6 wbs_adr_o[28]
port 303 nsew signal output
rlabel metal2 s 40774 79200 40830 80800 6 wbs_adr_o[29]
port 304 nsew signal output
rlabel metal2 s 45742 79200 45798 80800 6 wbs_adr_o[2]
port 305 nsew signal output
rlabel metal2 s 40590 79200 40646 80800 6 wbs_adr_o[30]
port 306 nsew signal output
rlabel metal2 s 40406 79200 40462 80800 6 wbs_adr_o[31]
port 307 nsew signal output
rlabel metal2 s 45558 79200 45614 80800 6 wbs_adr_o[3]
port 308 nsew signal output
rlabel metal2 s 45374 79200 45430 80800 6 wbs_adr_o[4]
port 309 nsew signal output
rlabel metal2 s 45190 79200 45246 80800 6 wbs_adr_o[5]
port 310 nsew signal output
rlabel metal2 s 45006 79200 45062 80800 6 wbs_adr_o[6]
port 311 nsew signal output
rlabel metal2 s 44822 79200 44878 80800 6 wbs_adr_o[7]
port 312 nsew signal output
rlabel metal2 s 44638 79200 44694 80800 6 wbs_adr_o[8]
port 313 nsew signal output
rlabel metal2 s 44454 79200 44510 80800 6 wbs_adr_o[9]
port 314 nsew signal output
rlabel metal2 s 33414 79200 33470 80800 6 wbs_clk_i
port 315 nsew signal input
rlabel metal2 s 33230 79200 33286 80800 6 wbs_clk_out
port 316 nsew signal output
rlabel metal2 s 59174 79200 59230 80800 6 wbs_cyc_o
port 317 nsew signal output
rlabel metal2 s 58622 79200 58678 80800 6 wbs_dat_i[0]
port 318 nsew signal input
rlabel metal2 s 56782 79200 56838 80800 6 wbs_dat_i[10]
port 319 nsew signal input
rlabel metal2 s 56598 79200 56654 80800 6 wbs_dat_i[11]
port 320 nsew signal input
rlabel metal2 s 56414 79200 56470 80800 6 wbs_dat_i[12]
port 321 nsew signal input
rlabel metal2 s 56230 79200 56286 80800 6 wbs_dat_i[13]
port 322 nsew signal input
rlabel metal2 s 56046 79200 56102 80800 6 wbs_dat_i[14]
port 323 nsew signal input
rlabel metal2 s 55862 79200 55918 80800 6 wbs_dat_i[15]
port 324 nsew signal input
rlabel metal2 s 55678 79200 55734 80800 6 wbs_dat_i[16]
port 325 nsew signal input
rlabel metal2 s 55494 79200 55550 80800 6 wbs_dat_i[17]
port 326 nsew signal input
rlabel metal2 s 55310 79200 55366 80800 6 wbs_dat_i[18]
port 327 nsew signal input
rlabel metal2 s 55126 79200 55182 80800 6 wbs_dat_i[19]
port 328 nsew signal input
rlabel metal2 s 58438 79200 58494 80800 6 wbs_dat_i[1]
port 329 nsew signal input
rlabel metal2 s 54942 79200 54998 80800 6 wbs_dat_i[20]
port 330 nsew signal input
rlabel metal2 s 54758 79200 54814 80800 6 wbs_dat_i[21]
port 331 nsew signal input
rlabel metal2 s 54574 79200 54630 80800 6 wbs_dat_i[22]
port 332 nsew signal input
rlabel metal2 s 54390 79200 54446 80800 6 wbs_dat_i[23]
port 333 nsew signal input
rlabel metal2 s 54206 79200 54262 80800 6 wbs_dat_i[24]
port 334 nsew signal input
rlabel metal2 s 54022 79200 54078 80800 6 wbs_dat_i[25]
port 335 nsew signal input
rlabel metal2 s 53838 79200 53894 80800 6 wbs_dat_i[26]
port 336 nsew signal input
rlabel metal2 s 53654 79200 53710 80800 6 wbs_dat_i[27]
port 337 nsew signal input
rlabel metal2 s 53470 79200 53526 80800 6 wbs_dat_i[28]
port 338 nsew signal input
rlabel metal2 s 53286 79200 53342 80800 6 wbs_dat_i[29]
port 339 nsew signal input
rlabel metal2 s 58254 79200 58310 80800 6 wbs_dat_i[2]
port 340 nsew signal input
rlabel metal2 s 53102 79200 53158 80800 6 wbs_dat_i[30]
port 341 nsew signal input
rlabel metal2 s 52918 79200 52974 80800 6 wbs_dat_i[31]
port 342 nsew signal input
rlabel metal2 s 58070 79200 58126 80800 6 wbs_dat_i[3]
port 343 nsew signal input
rlabel metal2 s 57886 79200 57942 80800 6 wbs_dat_i[4]
port 344 nsew signal input
rlabel metal2 s 57702 79200 57758 80800 6 wbs_dat_i[5]
port 345 nsew signal input
rlabel metal2 s 57518 79200 57574 80800 6 wbs_dat_i[6]
port 346 nsew signal input
rlabel metal2 s 57334 79200 57390 80800 6 wbs_dat_i[7]
port 347 nsew signal input
rlabel metal2 s 57150 79200 57206 80800 6 wbs_dat_i[8]
port 348 nsew signal input
rlabel metal2 s 56966 79200 57022 80800 6 wbs_dat_i[9]
port 349 nsew signal input
rlabel metal2 s 52734 79200 52790 80800 6 wbs_dat_o[0]
port 350 nsew signal output
rlabel metal2 s 50894 79200 50950 80800 6 wbs_dat_o[10]
port 351 nsew signal output
rlabel metal2 s 50710 79200 50766 80800 6 wbs_dat_o[11]
port 352 nsew signal output
rlabel metal2 s 50526 79200 50582 80800 6 wbs_dat_o[12]
port 353 nsew signal output
rlabel metal2 s 50342 79200 50398 80800 6 wbs_dat_o[13]
port 354 nsew signal output
rlabel metal2 s 50158 79200 50214 80800 6 wbs_dat_o[14]
port 355 nsew signal output
rlabel metal2 s 49974 79200 50030 80800 6 wbs_dat_o[15]
port 356 nsew signal output
rlabel metal2 s 49790 79200 49846 80800 6 wbs_dat_o[16]
port 357 nsew signal output
rlabel metal2 s 49606 79200 49662 80800 6 wbs_dat_o[17]
port 358 nsew signal output
rlabel metal2 s 49422 79200 49478 80800 6 wbs_dat_o[18]
port 359 nsew signal output
rlabel metal2 s 49238 79200 49294 80800 6 wbs_dat_o[19]
port 360 nsew signal output
rlabel metal2 s 52550 79200 52606 80800 6 wbs_dat_o[1]
port 361 nsew signal output
rlabel metal2 s 49054 79200 49110 80800 6 wbs_dat_o[20]
port 362 nsew signal output
rlabel metal2 s 48870 79200 48926 80800 6 wbs_dat_o[21]
port 363 nsew signal output
rlabel metal2 s 48686 79200 48742 80800 6 wbs_dat_o[22]
port 364 nsew signal output
rlabel metal2 s 48502 79200 48558 80800 6 wbs_dat_o[23]
port 365 nsew signal output
rlabel metal2 s 48318 79200 48374 80800 6 wbs_dat_o[24]
port 366 nsew signal output
rlabel metal2 s 48134 79200 48190 80800 6 wbs_dat_o[25]
port 367 nsew signal output
rlabel metal2 s 47950 79200 48006 80800 6 wbs_dat_o[26]
port 368 nsew signal output
rlabel metal2 s 47766 79200 47822 80800 6 wbs_dat_o[27]
port 369 nsew signal output
rlabel metal2 s 47582 79200 47638 80800 6 wbs_dat_o[28]
port 370 nsew signal output
rlabel metal2 s 47398 79200 47454 80800 6 wbs_dat_o[29]
port 371 nsew signal output
rlabel metal2 s 52366 79200 52422 80800 6 wbs_dat_o[2]
port 372 nsew signal output
rlabel metal2 s 47214 79200 47270 80800 6 wbs_dat_o[30]
port 373 nsew signal output
rlabel metal2 s 47030 79200 47086 80800 6 wbs_dat_o[31]
port 374 nsew signal output
rlabel metal2 s 52182 79200 52238 80800 6 wbs_dat_o[3]
port 375 nsew signal output
rlabel metal2 s 51998 79200 52054 80800 6 wbs_dat_o[4]
port 376 nsew signal output
rlabel metal2 s 51814 79200 51870 80800 6 wbs_dat_o[5]
port 377 nsew signal output
rlabel metal2 s 51630 79200 51686 80800 6 wbs_dat_o[6]
port 378 nsew signal output
rlabel metal2 s 51446 79200 51502 80800 6 wbs_dat_o[7]
port 379 nsew signal output
rlabel metal2 s 51262 79200 51318 80800 6 wbs_dat_o[8]
port 380 nsew signal output
rlabel metal2 s 51078 79200 51134 80800 6 wbs_dat_o[9]
port 381 nsew signal output
rlabel metal2 s 58990 79200 59046 80800 6 wbs_err_i
port 382 nsew signal input
rlabel metal2 s 46846 79200 46902 80800 6 wbs_sel_o[0]
port 383 nsew signal output
rlabel metal2 s 46662 79200 46718 80800 6 wbs_sel_o[1]
port 384 nsew signal output
rlabel metal2 s 46478 79200 46534 80800 6 wbs_sel_o[2]
port 385 nsew signal output
rlabel metal2 s 46294 79200 46350 80800 6 wbs_sel_o[3]
port 386 nsew signal output
rlabel metal2 s 40038 79200 40094 80800 6 wbs_stb_o
port 387 nsew signal output
rlabel metal2 s 40222 79200 40278 80800 6 wbs_we_o
port 388 nsew signal output
rlabel metal2 s 80150 79200 80206 80800 6 xtal_clk
port 389 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 90000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 20737318
string GDS_FILE /home/lx/projects/caravel_env/caravel_usb_test/openlane/wb_host/runs/wb_host/results/signoff/wb_host.magic.gds
string GDS_START 959072
<< end >>

