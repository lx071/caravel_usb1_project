// This is the unpowered netlist.
module wb_host (cfg_fast_sim,
    cfg_strap_pad_ctrl,
    cpu_clk,
    e_reset_n,
    int_pll_clock,
    p_reset_n,
    s_reset_n,
    sclk,
    sdin,
    sdout,
    sdout_oen,
    ssn,
    uartm_rxd,
    uartm_txd,
    user_clock1,
    user_clock2,
    wbd_clk_int,
    wbd_clk_wh,
    wbd_int_rst_n,
    wbd_pll_rst_n,
    wbm_ack_o,
    wbm_clk_i,
    wbm_cyc_i,
    wbm_err_o,
    wbm_rst_i,
    wbm_stb_i,
    wbm_we_i,
    wbs_ack_i,
    wbs_clk_i,
    wbs_clk_out,
    wbs_cyc_o,
    wbs_err_i,
    wbs_stb_o,
    wbs_we_o,
    xtal_clk,
    cfg_clk_skew_ctrl1,
    cfg_clk_skew_ctrl2,
    cfg_cska_wh,
    la_data_in,
    strap_sticky,
    strap_uartm,
    system_strap,
    wbm_adr_i,
    wbm_dat_i,
    wbm_dat_o,
    wbm_sel_i,
    wbs_adr_o,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_o);
 output cfg_fast_sim;
 output cfg_strap_pad_ctrl;
 output cpu_clk;
 output e_reset_n;
 input int_pll_clock;
 output p_reset_n;
 output s_reset_n;
 input sclk;
 input sdin;
 output sdout;
 output sdout_oen;
 input ssn;
 input uartm_rxd;
 output uartm_txd;
 input user_clock1;
 input user_clock2;
 input wbd_clk_int;
 output wbd_clk_wh;
 output wbd_int_rst_n;
 output wbd_pll_rst_n;
 output wbm_ack_o;
 input wbm_clk_i;
 input wbm_cyc_i;
 output wbm_err_o;
 input wbm_rst_i;
 input wbm_stb_i;
 input wbm_we_i;
 input wbs_ack_i;
 input wbs_clk_i;
 output wbs_clk_out;
 output wbs_cyc_o;
 input wbs_err_i;
 output wbs_stb_o;
 output wbs_we_o;
 input xtal_clk;
 output [31:0] cfg_clk_skew_ctrl1;
 output [31:0] cfg_clk_skew_ctrl2;
 input [3:0] cfg_cska_wh;
 input [17:0] la_data_in;
 input [31:0] strap_sticky;
 input [1:0] strap_uartm;
 output [31:0] system_strap;
 input [31:0] wbm_adr_i;
 input [31:0] wbm_dat_i;
 output [31:0] wbm_dat_o;
 input [3:0] wbm_sel_i;
 output [31:0] wbs_adr_o;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 output [3:0] wbs_sel_o;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire \clknet_0_u_async_wb.u_cmd_if.rd_clk ;
 wire \clknet_0_u_uart2wb.baud_clk_16x ;
 wire clknet_0_wbm_clk_i;
 wire \clknet_1_0__leaf_u_uart2wb.baud_clk_16x ;
 wire \clknet_1_1__leaf_u_uart2wb.baud_clk_16x ;
 wire \clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ;
 wire clknet_3_0__leaf_wbm_clk_i;
 wire \clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ;
 wire clknet_3_1__leaf_wbm_clk_i;
 wire \clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ;
 wire clknet_3_2__leaf_wbm_clk_i;
 wire \clknet_3_3__leaf_u_async_wb.u_cmd_if.rd_clk ;
 wire clknet_3_3__leaf_wbm_clk_i;
 wire \clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ;
 wire clknet_3_4__leaf_wbm_clk_i;
 wire \clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ;
 wire clknet_3_5__leaf_wbm_clk_i;
 wire \clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ;
 wire clknet_3_6__leaf_wbm_clk_i;
 wire \clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ;
 wire clknet_3_7__leaf_wbm_clk_i;
 wire \clknet_leaf_0_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_0_wbm_clk_i;
 wire \clknet_leaf_10_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_10_wbm_clk_i;
 wire \clknet_leaf_11_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_11_wbm_clk_i;
 wire \clknet_leaf_12_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_12_wbm_clk_i;
 wire \clknet_leaf_13_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_13_wbm_clk_i;
 wire \clknet_leaf_14_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_14_wbm_clk_i;
 wire \clknet_leaf_15_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_15_wbm_clk_i;
 wire \clknet_leaf_16_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_16_wbm_clk_i;
 wire \clknet_leaf_17_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_17_wbm_clk_i;
 wire \clknet_leaf_18_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_18_wbm_clk_i;
 wire \clknet_leaf_19_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_19_wbm_clk_i;
 wire \clknet_leaf_1_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_1_wbm_clk_i;
 wire \clknet_leaf_20_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_20_wbm_clk_i;
 wire \clknet_leaf_21_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_21_wbm_clk_i;
 wire \clknet_leaf_22_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_22_wbm_clk_i;
 wire \clknet_leaf_23_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_23_wbm_clk_i;
 wire \clknet_leaf_24_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_24_wbm_clk_i;
 wire \clknet_leaf_25_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_25_wbm_clk_i;
 wire \clknet_leaf_26_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_26_wbm_clk_i;
 wire \clknet_leaf_27_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_27_wbm_clk_i;
 wire clknet_leaf_28_wbm_clk_i;
 wire clknet_leaf_29_wbm_clk_i;
 wire \clknet_leaf_2_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_2_wbm_clk_i;
 wire clknet_leaf_30_wbm_clk_i;
 wire clknet_leaf_31_wbm_clk_i;
 wire clknet_leaf_32_wbm_clk_i;
 wire clknet_leaf_33_wbm_clk_i;
 wire clknet_leaf_34_wbm_clk_i;
 wire clknet_leaf_35_wbm_clk_i;
 wire clknet_leaf_36_wbm_clk_i;
 wire clknet_leaf_37_wbm_clk_i;
 wire clknet_leaf_38_wbm_clk_i;
 wire clknet_leaf_39_wbm_clk_i;
 wire \clknet_leaf_3_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_3_wbm_clk_i;
 wire clknet_leaf_40_wbm_clk_i;
 wire clknet_leaf_41_wbm_clk_i;
 wire clknet_leaf_42_wbm_clk_i;
 wire clknet_leaf_43_wbm_clk_i;
 wire clknet_leaf_44_wbm_clk_i;
 wire clknet_leaf_45_wbm_clk_i;
 wire clknet_leaf_46_wbm_clk_i;
 wire clknet_leaf_47_wbm_clk_i;
 wire clknet_leaf_48_wbm_clk_i;
 wire clknet_leaf_49_wbm_clk_i;
 wire \clknet_leaf_4_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_4_wbm_clk_i;
 wire clknet_leaf_50_wbm_clk_i;
 wire clknet_leaf_51_wbm_clk_i;
 wire clknet_leaf_52_wbm_clk_i;
 wire clknet_leaf_53_wbm_clk_i;
 wire clknet_leaf_54_wbm_clk_i;
 wire clknet_leaf_55_wbm_clk_i;
 wire clknet_leaf_56_wbm_clk_i;
 wire clknet_leaf_57_wbm_clk_i;
 wire clknet_leaf_58_wbm_clk_i;
 wire clknet_leaf_59_wbm_clk_i;
 wire \clknet_leaf_5_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_5_wbm_clk_i;
 wire clknet_leaf_60_wbm_clk_i;
 wire clknet_leaf_61_wbm_clk_i;
 wire clknet_leaf_62_wbm_clk_i;
 wire clknet_leaf_63_wbm_clk_i;
 wire clknet_leaf_64_wbm_clk_i;
 wire clknet_leaf_65_wbm_clk_i;
 wire clknet_leaf_66_wbm_clk_i;
 wire clknet_leaf_67_wbm_clk_i;
 wire clknet_leaf_68_wbm_clk_i;
 wire clknet_leaf_69_wbm_clk_i;
 wire \clknet_leaf_6_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_6_wbm_clk_i;
 wire clknet_leaf_70_wbm_clk_i;
 wire clknet_leaf_71_wbm_clk_i;
 wire clknet_leaf_72_wbm_clk_i;
 wire clknet_leaf_73_wbm_clk_i;
 wire clknet_leaf_74_wbm_clk_i;
 wire clknet_leaf_75_wbm_clk_i;
 wire clknet_leaf_76_wbm_clk_i;
 wire clknet_leaf_77_wbm_clk_i;
 wire clknet_leaf_78_wbm_clk_i;
 wire clknet_leaf_79_wbm_clk_i;
 wire \clknet_leaf_7_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_7_wbm_clk_i;
 wire clknet_leaf_80_wbm_clk_i;
 wire clknet_leaf_81_wbm_clk_i;
 wire clknet_leaf_82_wbm_clk_i;
 wire clknet_leaf_83_wbm_clk_i;
 wire clknet_leaf_84_wbm_clk_i;
 wire clknet_leaf_85_wbm_clk_i;
 wire clknet_leaf_86_wbm_clk_i;
 wire clknet_leaf_87_wbm_clk_i;
 wire clknet_leaf_88_wbm_clk_i;
 wire clknet_leaf_89_wbm_clk_i;
 wire \clknet_leaf_8_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_8_wbm_clk_i;
 wire clknet_leaf_90_wbm_clk_i;
 wire clknet_leaf_91_wbm_clk_i;
 wire clknet_leaf_92_wbm_clk_i;
 wire clknet_leaf_93_wbm_clk_i;
 wire clknet_leaf_94_wbm_clk_i;
 wire \clknet_leaf_9_u_uart2wb.baud_clk_16x ;
 wire clknet_leaf_9_wbm_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \u_arb.gnt[0] ;
 wire \u_arb.gnt[1] ;
 wire \u_async_wb.PendingRd ;
 wire \u_async_wb.m_cmd_wr_data[56] ;
 wire \u_async_wb.m_cmd_wr_data[57] ;
 wire \u_async_wb.m_cmd_wr_data[58] ;
 wire \u_async_wb.m_cmd_wr_data[59] ;
 wire \u_async_wb.m_cmd_wr_data[60] ;
 wire \u_async_wb.m_cmd_wr_data[61] ;
 wire \u_async_wb.m_cmd_wr_data[62] ;
 wire \u_async_wb.m_cmd_wr_data[63] ;
 wire \u_async_wb.m_cmd_wr_data[64] ;
 wire \u_async_wb.m_cmd_wr_data[65] ;
 wire \u_async_wb.m_cmd_wr_data[66] ;
 wire \u_async_wb.m_cmd_wr_data[67] ;
 wire \u_async_wb.m_cmd_wr_data[68] ;
 wire \u_async_wb.u_cmd_if.grey_rd_ptr[0] ;
 wire \u_async_wb.u_cmd_if.grey_rd_ptr[1] ;
 wire \u_async_wb.u_cmd_if.grey_rd_ptr[2] ;
 wire \u_async_wb.u_cmd_if.grey_wr_ptr[0] ;
 wire \u_async_wb.u_cmd_if.grey_wr_ptr[1] ;
 wire \u_async_wb.u_cmd_if.grey_wr_ptr[2] ;
 wire \u_async_wb.u_cmd_if.mem[0][0] ;
 wire \u_async_wb.u_cmd_if.mem[0][10] ;
 wire \u_async_wb.u_cmd_if.mem[0][11] ;
 wire \u_async_wb.u_cmd_if.mem[0][12] ;
 wire \u_async_wb.u_cmd_if.mem[0][13] ;
 wire \u_async_wb.u_cmd_if.mem[0][14] ;
 wire \u_async_wb.u_cmd_if.mem[0][15] ;
 wire \u_async_wb.u_cmd_if.mem[0][16] ;
 wire \u_async_wb.u_cmd_if.mem[0][17] ;
 wire \u_async_wb.u_cmd_if.mem[0][18] ;
 wire \u_async_wb.u_cmd_if.mem[0][19] ;
 wire \u_async_wb.u_cmd_if.mem[0][1] ;
 wire \u_async_wb.u_cmd_if.mem[0][20] ;
 wire \u_async_wb.u_cmd_if.mem[0][21] ;
 wire \u_async_wb.u_cmd_if.mem[0][22] ;
 wire \u_async_wb.u_cmd_if.mem[0][23] ;
 wire \u_async_wb.u_cmd_if.mem[0][24] ;
 wire \u_async_wb.u_cmd_if.mem[0][25] ;
 wire \u_async_wb.u_cmd_if.mem[0][26] ;
 wire \u_async_wb.u_cmd_if.mem[0][27] ;
 wire \u_async_wb.u_cmd_if.mem[0][28] ;
 wire \u_async_wb.u_cmd_if.mem[0][29] ;
 wire \u_async_wb.u_cmd_if.mem[0][2] ;
 wire \u_async_wb.u_cmd_if.mem[0][30] ;
 wire \u_async_wb.u_cmd_if.mem[0][31] ;
 wire \u_async_wb.u_cmd_if.mem[0][32] ;
 wire \u_async_wb.u_cmd_if.mem[0][33] ;
 wire \u_async_wb.u_cmd_if.mem[0][34] ;
 wire \u_async_wb.u_cmd_if.mem[0][35] ;
 wire \u_async_wb.u_cmd_if.mem[0][36] ;
 wire \u_async_wb.u_cmd_if.mem[0][37] ;
 wire \u_async_wb.u_cmd_if.mem[0][38] ;
 wire \u_async_wb.u_cmd_if.mem[0][39] ;
 wire \u_async_wb.u_cmd_if.mem[0][3] ;
 wire \u_async_wb.u_cmd_if.mem[0][40] ;
 wire \u_async_wb.u_cmd_if.mem[0][41] ;
 wire \u_async_wb.u_cmd_if.mem[0][42] ;
 wire \u_async_wb.u_cmd_if.mem[0][43] ;
 wire \u_async_wb.u_cmd_if.mem[0][44] ;
 wire \u_async_wb.u_cmd_if.mem[0][45] ;
 wire \u_async_wb.u_cmd_if.mem[0][46] ;
 wire \u_async_wb.u_cmd_if.mem[0][47] ;
 wire \u_async_wb.u_cmd_if.mem[0][48] ;
 wire \u_async_wb.u_cmd_if.mem[0][49] ;
 wire \u_async_wb.u_cmd_if.mem[0][4] ;
 wire \u_async_wb.u_cmd_if.mem[0][50] ;
 wire \u_async_wb.u_cmd_if.mem[0][51] ;
 wire \u_async_wb.u_cmd_if.mem[0][52] ;
 wire \u_async_wb.u_cmd_if.mem[0][53] ;
 wire \u_async_wb.u_cmd_if.mem[0][54] ;
 wire \u_async_wb.u_cmd_if.mem[0][55] ;
 wire \u_async_wb.u_cmd_if.mem[0][56] ;
 wire \u_async_wb.u_cmd_if.mem[0][57] ;
 wire \u_async_wb.u_cmd_if.mem[0][58] ;
 wire \u_async_wb.u_cmd_if.mem[0][59] ;
 wire \u_async_wb.u_cmd_if.mem[0][5] ;
 wire \u_async_wb.u_cmd_if.mem[0][60] ;
 wire \u_async_wb.u_cmd_if.mem[0][61] ;
 wire \u_async_wb.u_cmd_if.mem[0][62] ;
 wire \u_async_wb.u_cmd_if.mem[0][63] ;
 wire \u_async_wb.u_cmd_if.mem[0][64] ;
 wire \u_async_wb.u_cmd_if.mem[0][65] ;
 wire \u_async_wb.u_cmd_if.mem[0][66] ;
 wire \u_async_wb.u_cmd_if.mem[0][67] ;
 wire \u_async_wb.u_cmd_if.mem[0][68] ;
 wire \u_async_wb.u_cmd_if.mem[0][6] ;
 wire \u_async_wb.u_cmd_if.mem[0][7] ;
 wire \u_async_wb.u_cmd_if.mem[0][8] ;
 wire \u_async_wb.u_cmd_if.mem[0][9] ;
 wire \u_async_wb.u_cmd_if.mem[1][0] ;
 wire \u_async_wb.u_cmd_if.mem[1][10] ;
 wire \u_async_wb.u_cmd_if.mem[1][11] ;
 wire \u_async_wb.u_cmd_if.mem[1][12] ;
 wire \u_async_wb.u_cmd_if.mem[1][13] ;
 wire \u_async_wb.u_cmd_if.mem[1][14] ;
 wire \u_async_wb.u_cmd_if.mem[1][15] ;
 wire \u_async_wb.u_cmd_if.mem[1][16] ;
 wire \u_async_wb.u_cmd_if.mem[1][17] ;
 wire \u_async_wb.u_cmd_if.mem[1][18] ;
 wire \u_async_wb.u_cmd_if.mem[1][19] ;
 wire \u_async_wb.u_cmd_if.mem[1][1] ;
 wire \u_async_wb.u_cmd_if.mem[1][20] ;
 wire \u_async_wb.u_cmd_if.mem[1][21] ;
 wire \u_async_wb.u_cmd_if.mem[1][22] ;
 wire \u_async_wb.u_cmd_if.mem[1][23] ;
 wire \u_async_wb.u_cmd_if.mem[1][24] ;
 wire \u_async_wb.u_cmd_if.mem[1][25] ;
 wire \u_async_wb.u_cmd_if.mem[1][26] ;
 wire \u_async_wb.u_cmd_if.mem[1][27] ;
 wire \u_async_wb.u_cmd_if.mem[1][28] ;
 wire \u_async_wb.u_cmd_if.mem[1][29] ;
 wire \u_async_wb.u_cmd_if.mem[1][2] ;
 wire \u_async_wb.u_cmd_if.mem[1][30] ;
 wire \u_async_wb.u_cmd_if.mem[1][31] ;
 wire \u_async_wb.u_cmd_if.mem[1][32] ;
 wire \u_async_wb.u_cmd_if.mem[1][33] ;
 wire \u_async_wb.u_cmd_if.mem[1][34] ;
 wire \u_async_wb.u_cmd_if.mem[1][35] ;
 wire \u_async_wb.u_cmd_if.mem[1][36] ;
 wire \u_async_wb.u_cmd_if.mem[1][37] ;
 wire \u_async_wb.u_cmd_if.mem[1][38] ;
 wire \u_async_wb.u_cmd_if.mem[1][39] ;
 wire \u_async_wb.u_cmd_if.mem[1][3] ;
 wire \u_async_wb.u_cmd_if.mem[1][40] ;
 wire \u_async_wb.u_cmd_if.mem[1][41] ;
 wire \u_async_wb.u_cmd_if.mem[1][42] ;
 wire \u_async_wb.u_cmd_if.mem[1][43] ;
 wire \u_async_wb.u_cmd_if.mem[1][44] ;
 wire \u_async_wb.u_cmd_if.mem[1][45] ;
 wire \u_async_wb.u_cmd_if.mem[1][46] ;
 wire \u_async_wb.u_cmd_if.mem[1][47] ;
 wire \u_async_wb.u_cmd_if.mem[1][48] ;
 wire \u_async_wb.u_cmd_if.mem[1][49] ;
 wire \u_async_wb.u_cmd_if.mem[1][4] ;
 wire \u_async_wb.u_cmd_if.mem[1][50] ;
 wire \u_async_wb.u_cmd_if.mem[1][51] ;
 wire \u_async_wb.u_cmd_if.mem[1][52] ;
 wire \u_async_wb.u_cmd_if.mem[1][53] ;
 wire \u_async_wb.u_cmd_if.mem[1][54] ;
 wire \u_async_wb.u_cmd_if.mem[1][55] ;
 wire \u_async_wb.u_cmd_if.mem[1][56] ;
 wire \u_async_wb.u_cmd_if.mem[1][57] ;
 wire \u_async_wb.u_cmd_if.mem[1][58] ;
 wire \u_async_wb.u_cmd_if.mem[1][59] ;
 wire \u_async_wb.u_cmd_if.mem[1][5] ;
 wire \u_async_wb.u_cmd_if.mem[1][60] ;
 wire \u_async_wb.u_cmd_if.mem[1][61] ;
 wire \u_async_wb.u_cmd_if.mem[1][62] ;
 wire \u_async_wb.u_cmd_if.mem[1][63] ;
 wire \u_async_wb.u_cmd_if.mem[1][64] ;
 wire \u_async_wb.u_cmd_if.mem[1][65] ;
 wire \u_async_wb.u_cmd_if.mem[1][66] ;
 wire \u_async_wb.u_cmd_if.mem[1][67] ;
 wire \u_async_wb.u_cmd_if.mem[1][68] ;
 wire \u_async_wb.u_cmd_if.mem[1][6] ;
 wire \u_async_wb.u_cmd_if.mem[1][7] ;
 wire \u_async_wb.u_cmd_if.mem[1][8] ;
 wire \u_async_wb.u_cmd_if.mem[1][9] ;
 wire \u_async_wb.u_cmd_if.mem[2][0] ;
 wire \u_async_wb.u_cmd_if.mem[2][10] ;
 wire \u_async_wb.u_cmd_if.mem[2][11] ;
 wire \u_async_wb.u_cmd_if.mem[2][12] ;
 wire \u_async_wb.u_cmd_if.mem[2][13] ;
 wire \u_async_wb.u_cmd_if.mem[2][14] ;
 wire \u_async_wb.u_cmd_if.mem[2][15] ;
 wire \u_async_wb.u_cmd_if.mem[2][16] ;
 wire \u_async_wb.u_cmd_if.mem[2][17] ;
 wire \u_async_wb.u_cmd_if.mem[2][18] ;
 wire \u_async_wb.u_cmd_if.mem[2][19] ;
 wire \u_async_wb.u_cmd_if.mem[2][1] ;
 wire \u_async_wb.u_cmd_if.mem[2][20] ;
 wire \u_async_wb.u_cmd_if.mem[2][21] ;
 wire \u_async_wb.u_cmd_if.mem[2][22] ;
 wire \u_async_wb.u_cmd_if.mem[2][23] ;
 wire \u_async_wb.u_cmd_if.mem[2][24] ;
 wire \u_async_wb.u_cmd_if.mem[2][25] ;
 wire \u_async_wb.u_cmd_if.mem[2][26] ;
 wire \u_async_wb.u_cmd_if.mem[2][27] ;
 wire \u_async_wb.u_cmd_if.mem[2][28] ;
 wire \u_async_wb.u_cmd_if.mem[2][29] ;
 wire \u_async_wb.u_cmd_if.mem[2][2] ;
 wire \u_async_wb.u_cmd_if.mem[2][30] ;
 wire \u_async_wb.u_cmd_if.mem[2][31] ;
 wire \u_async_wb.u_cmd_if.mem[2][32] ;
 wire \u_async_wb.u_cmd_if.mem[2][33] ;
 wire \u_async_wb.u_cmd_if.mem[2][34] ;
 wire \u_async_wb.u_cmd_if.mem[2][35] ;
 wire \u_async_wb.u_cmd_if.mem[2][36] ;
 wire \u_async_wb.u_cmd_if.mem[2][37] ;
 wire \u_async_wb.u_cmd_if.mem[2][38] ;
 wire \u_async_wb.u_cmd_if.mem[2][39] ;
 wire \u_async_wb.u_cmd_if.mem[2][3] ;
 wire \u_async_wb.u_cmd_if.mem[2][40] ;
 wire \u_async_wb.u_cmd_if.mem[2][41] ;
 wire \u_async_wb.u_cmd_if.mem[2][42] ;
 wire \u_async_wb.u_cmd_if.mem[2][43] ;
 wire \u_async_wb.u_cmd_if.mem[2][44] ;
 wire \u_async_wb.u_cmd_if.mem[2][45] ;
 wire \u_async_wb.u_cmd_if.mem[2][46] ;
 wire \u_async_wb.u_cmd_if.mem[2][47] ;
 wire \u_async_wb.u_cmd_if.mem[2][48] ;
 wire \u_async_wb.u_cmd_if.mem[2][49] ;
 wire \u_async_wb.u_cmd_if.mem[2][4] ;
 wire \u_async_wb.u_cmd_if.mem[2][50] ;
 wire \u_async_wb.u_cmd_if.mem[2][51] ;
 wire \u_async_wb.u_cmd_if.mem[2][52] ;
 wire \u_async_wb.u_cmd_if.mem[2][53] ;
 wire \u_async_wb.u_cmd_if.mem[2][54] ;
 wire \u_async_wb.u_cmd_if.mem[2][55] ;
 wire \u_async_wb.u_cmd_if.mem[2][56] ;
 wire \u_async_wb.u_cmd_if.mem[2][57] ;
 wire \u_async_wb.u_cmd_if.mem[2][58] ;
 wire \u_async_wb.u_cmd_if.mem[2][59] ;
 wire \u_async_wb.u_cmd_if.mem[2][5] ;
 wire \u_async_wb.u_cmd_if.mem[2][60] ;
 wire \u_async_wb.u_cmd_if.mem[2][61] ;
 wire \u_async_wb.u_cmd_if.mem[2][62] ;
 wire \u_async_wb.u_cmd_if.mem[2][63] ;
 wire \u_async_wb.u_cmd_if.mem[2][64] ;
 wire \u_async_wb.u_cmd_if.mem[2][65] ;
 wire \u_async_wb.u_cmd_if.mem[2][66] ;
 wire \u_async_wb.u_cmd_if.mem[2][67] ;
 wire \u_async_wb.u_cmd_if.mem[2][68] ;
 wire \u_async_wb.u_cmd_if.mem[2][6] ;
 wire \u_async_wb.u_cmd_if.mem[2][7] ;
 wire \u_async_wb.u_cmd_if.mem[2][8] ;
 wire \u_async_wb.u_cmd_if.mem[2][9] ;
 wire \u_async_wb.u_cmd_if.mem[3][0] ;
 wire \u_async_wb.u_cmd_if.mem[3][10] ;
 wire \u_async_wb.u_cmd_if.mem[3][11] ;
 wire \u_async_wb.u_cmd_if.mem[3][12] ;
 wire \u_async_wb.u_cmd_if.mem[3][13] ;
 wire \u_async_wb.u_cmd_if.mem[3][14] ;
 wire \u_async_wb.u_cmd_if.mem[3][15] ;
 wire \u_async_wb.u_cmd_if.mem[3][16] ;
 wire \u_async_wb.u_cmd_if.mem[3][17] ;
 wire \u_async_wb.u_cmd_if.mem[3][18] ;
 wire \u_async_wb.u_cmd_if.mem[3][19] ;
 wire \u_async_wb.u_cmd_if.mem[3][1] ;
 wire \u_async_wb.u_cmd_if.mem[3][20] ;
 wire \u_async_wb.u_cmd_if.mem[3][21] ;
 wire \u_async_wb.u_cmd_if.mem[3][22] ;
 wire \u_async_wb.u_cmd_if.mem[3][23] ;
 wire \u_async_wb.u_cmd_if.mem[3][24] ;
 wire \u_async_wb.u_cmd_if.mem[3][25] ;
 wire \u_async_wb.u_cmd_if.mem[3][26] ;
 wire \u_async_wb.u_cmd_if.mem[3][27] ;
 wire \u_async_wb.u_cmd_if.mem[3][28] ;
 wire \u_async_wb.u_cmd_if.mem[3][29] ;
 wire \u_async_wb.u_cmd_if.mem[3][2] ;
 wire \u_async_wb.u_cmd_if.mem[3][30] ;
 wire \u_async_wb.u_cmd_if.mem[3][31] ;
 wire \u_async_wb.u_cmd_if.mem[3][32] ;
 wire \u_async_wb.u_cmd_if.mem[3][33] ;
 wire \u_async_wb.u_cmd_if.mem[3][34] ;
 wire \u_async_wb.u_cmd_if.mem[3][35] ;
 wire \u_async_wb.u_cmd_if.mem[3][36] ;
 wire \u_async_wb.u_cmd_if.mem[3][37] ;
 wire \u_async_wb.u_cmd_if.mem[3][38] ;
 wire \u_async_wb.u_cmd_if.mem[3][39] ;
 wire \u_async_wb.u_cmd_if.mem[3][3] ;
 wire \u_async_wb.u_cmd_if.mem[3][40] ;
 wire \u_async_wb.u_cmd_if.mem[3][41] ;
 wire \u_async_wb.u_cmd_if.mem[3][42] ;
 wire \u_async_wb.u_cmd_if.mem[3][43] ;
 wire \u_async_wb.u_cmd_if.mem[3][44] ;
 wire \u_async_wb.u_cmd_if.mem[3][45] ;
 wire \u_async_wb.u_cmd_if.mem[3][46] ;
 wire \u_async_wb.u_cmd_if.mem[3][47] ;
 wire \u_async_wb.u_cmd_if.mem[3][48] ;
 wire \u_async_wb.u_cmd_if.mem[3][49] ;
 wire \u_async_wb.u_cmd_if.mem[3][4] ;
 wire \u_async_wb.u_cmd_if.mem[3][50] ;
 wire \u_async_wb.u_cmd_if.mem[3][51] ;
 wire \u_async_wb.u_cmd_if.mem[3][52] ;
 wire \u_async_wb.u_cmd_if.mem[3][53] ;
 wire \u_async_wb.u_cmd_if.mem[3][54] ;
 wire \u_async_wb.u_cmd_if.mem[3][55] ;
 wire \u_async_wb.u_cmd_if.mem[3][56] ;
 wire \u_async_wb.u_cmd_if.mem[3][57] ;
 wire \u_async_wb.u_cmd_if.mem[3][58] ;
 wire \u_async_wb.u_cmd_if.mem[3][59] ;
 wire \u_async_wb.u_cmd_if.mem[3][5] ;
 wire \u_async_wb.u_cmd_if.mem[3][60] ;
 wire \u_async_wb.u_cmd_if.mem[3][61] ;
 wire \u_async_wb.u_cmd_if.mem[3][62] ;
 wire \u_async_wb.u_cmd_if.mem[3][63] ;
 wire \u_async_wb.u_cmd_if.mem[3][64] ;
 wire \u_async_wb.u_cmd_if.mem[3][65] ;
 wire \u_async_wb.u_cmd_if.mem[3][66] ;
 wire \u_async_wb.u_cmd_if.mem[3][67] ;
 wire \u_async_wb.u_cmd_if.mem[3][68] ;
 wire \u_async_wb.u_cmd_if.mem[3][6] ;
 wire \u_async_wb.u_cmd_if.mem[3][7] ;
 wire \u_async_wb.u_cmd_if.mem[3][8] ;
 wire \u_async_wb.u_cmd_if.mem[3][9] ;
 wire \u_async_wb.u_cmd_if.rd_clk ;
 wire \u_async_wb.u_cmd_if.rd_ptr[0] ;
 wire \u_async_wb.u_cmd_if.rd_ptr[1] ;
 wire \u_async_wb.u_cmd_if.rd_reset_n ;
 wire \u_async_wb.u_cmd_if.sync_rd_ptr[2] ;
 wire \u_async_wb.u_cmd_if.sync_rd_ptr_0[0] ;
 wire \u_async_wb.u_cmd_if.sync_rd_ptr_0[1] ;
 wire \u_async_wb.u_cmd_if.sync_rd_ptr_0[2] ;
 wire \u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ;
 wire \u_async_wb.u_cmd_if.sync_rd_ptr_1[1] ;
 wire \u_async_wb.u_cmd_if.sync_wr_ptr[2] ;
 wire \u_async_wb.u_cmd_if.sync_wr_ptr_0[0] ;
 wire \u_async_wb.u_cmd_if.sync_wr_ptr_0[1] ;
 wire \u_async_wb.u_cmd_if.sync_wr_ptr_0[2] ;
 wire \u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ;
 wire \u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ;
 wire \u_async_wb.u_cmd_if.wr_ptr[0] ;
 wire \u_async_wb.u_cmd_if.wr_ptr[1] ;
 wire \u_async_wb.u_resp_if.grey_rd_ptr[0] ;
 wire \u_async_wb.u_resp_if.grey_rd_ptr[1] ;
 wire \u_async_wb.u_resp_if.grey_wr_ptr[0] ;
 wire \u_async_wb.u_resp_if.grey_wr_ptr[1] ;
 wire \u_async_wb.u_resp_if.mem[0][0] ;
 wire \u_async_wb.u_resp_if.mem[0][10] ;
 wire \u_async_wb.u_resp_if.mem[0][11] ;
 wire \u_async_wb.u_resp_if.mem[0][12] ;
 wire \u_async_wb.u_resp_if.mem[0][13] ;
 wire \u_async_wb.u_resp_if.mem[0][14] ;
 wire \u_async_wb.u_resp_if.mem[0][15] ;
 wire \u_async_wb.u_resp_if.mem[0][16] ;
 wire \u_async_wb.u_resp_if.mem[0][17] ;
 wire \u_async_wb.u_resp_if.mem[0][18] ;
 wire \u_async_wb.u_resp_if.mem[0][19] ;
 wire \u_async_wb.u_resp_if.mem[0][1] ;
 wire \u_async_wb.u_resp_if.mem[0][20] ;
 wire \u_async_wb.u_resp_if.mem[0][21] ;
 wire \u_async_wb.u_resp_if.mem[0][22] ;
 wire \u_async_wb.u_resp_if.mem[0][23] ;
 wire \u_async_wb.u_resp_if.mem[0][24] ;
 wire \u_async_wb.u_resp_if.mem[0][25] ;
 wire \u_async_wb.u_resp_if.mem[0][26] ;
 wire \u_async_wb.u_resp_if.mem[0][27] ;
 wire \u_async_wb.u_resp_if.mem[0][28] ;
 wire \u_async_wb.u_resp_if.mem[0][29] ;
 wire \u_async_wb.u_resp_if.mem[0][2] ;
 wire \u_async_wb.u_resp_if.mem[0][30] ;
 wire \u_async_wb.u_resp_if.mem[0][31] ;
 wire \u_async_wb.u_resp_if.mem[0][32] ;
 wire \u_async_wb.u_resp_if.mem[0][3] ;
 wire \u_async_wb.u_resp_if.mem[0][4] ;
 wire \u_async_wb.u_resp_if.mem[0][5] ;
 wire \u_async_wb.u_resp_if.mem[0][6] ;
 wire \u_async_wb.u_resp_if.mem[0][7] ;
 wire \u_async_wb.u_resp_if.mem[0][8] ;
 wire \u_async_wb.u_resp_if.mem[0][9] ;
 wire \u_async_wb.u_resp_if.mem[1][0] ;
 wire \u_async_wb.u_resp_if.mem[1][10] ;
 wire \u_async_wb.u_resp_if.mem[1][11] ;
 wire \u_async_wb.u_resp_if.mem[1][12] ;
 wire \u_async_wb.u_resp_if.mem[1][13] ;
 wire \u_async_wb.u_resp_if.mem[1][14] ;
 wire \u_async_wb.u_resp_if.mem[1][15] ;
 wire \u_async_wb.u_resp_if.mem[1][16] ;
 wire \u_async_wb.u_resp_if.mem[1][17] ;
 wire \u_async_wb.u_resp_if.mem[1][18] ;
 wire \u_async_wb.u_resp_if.mem[1][19] ;
 wire \u_async_wb.u_resp_if.mem[1][1] ;
 wire \u_async_wb.u_resp_if.mem[1][20] ;
 wire \u_async_wb.u_resp_if.mem[1][21] ;
 wire \u_async_wb.u_resp_if.mem[1][22] ;
 wire \u_async_wb.u_resp_if.mem[1][23] ;
 wire \u_async_wb.u_resp_if.mem[1][24] ;
 wire \u_async_wb.u_resp_if.mem[1][25] ;
 wire \u_async_wb.u_resp_if.mem[1][26] ;
 wire \u_async_wb.u_resp_if.mem[1][27] ;
 wire \u_async_wb.u_resp_if.mem[1][28] ;
 wire \u_async_wb.u_resp_if.mem[1][29] ;
 wire \u_async_wb.u_resp_if.mem[1][2] ;
 wire \u_async_wb.u_resp_if.mem[1][30] ;
 wire \u_async_wb.u_resp_if.mem[1][31] ;
 wire \u_async_wb.u_resp_if.mem[1][32] ;
 wire \u_async_wb.u_resp_if.mem[1][3] ;
 wire \u_async_wb.u_resp_if.mem[1][4] ;
 wire \u_async_wb.u_resp_if.mem[1][5] ;
 wire \u_async_wb.u_resp_if.mem[1][6] ;
 wire \u_async_wb.u_resp_if.mem[1][7] ;
 wire \u_async_wb.u_resp_if.mem[1][8] ;
 wire \u_async_wb.u_resp_if.mem[1][9] ;
 wire \u_async_wb.u_resp_if.rd_ptr[0] ;
 wire \u_async_wb.u_resp_if.rd_ptr[1] ;
 wire \u_async_wb.u_resp_if.sync_rd_ptr_0[0] ;
 wire \u_async_wb.u_resp_if.sync_rd_ptr_0[1] ;
 wire \u_async_wb.u_resp_if.sync_rd_ptr_1[0] ;
 wire \u_async_wb.u_resp_if.sync_rd_ptr_1[1] ;
 wire \u_async_wb.u_resp_if.sync_wr_ptr_0[0] ;
 wire \u_async_wb.u_resp_if.sync_wr_ptr_0[1] ;
 wire \u_async_wb.u_resp_if.sync_wr_ptr_1[0] ;
 wire \u_async_wb.u_resp_if.sync_wr_ptr_1[1] ;
 wire \u_async_wb.u_resp_if.wr_ptr[0] ;
 wire \u_async_wb.u_resp_if.wr_ptr[1] ;
 wire \u_async_wb.wbs_ack_f ;
 wire \u_delay1_stb0.A ;
 wire \u_delay1_stb0.X ;
 wire \u_delay2_stb1.X ;
 wire \u_delay2_stb2.X ;
 wire \u_reg.cfg_clk_ctrl[0] ;
 wire \u_reg.cfg_clk_ctrl[1] ;
 wire \u_reg.cfg_clk_ctrl[2] ;
 wire \u_reg.cfg_clk_ctrl[3] ;
 wire \u_reg.cfg_clk_ctrl[4] ;
 wire \u_reg.cfg_clk_ctrl[5] ;
 wire \u_reg.cfg_clk_ctrl[6] ;
 wire \u_reg.cfg_clk_ctrl[7] ;
 wire \u_reg.cfg_glb_ctrl[0] ;
 wire \u_reg.cfg_glb_ctrl[10] ;
 wire \u_reg.cfg_glb_ctrl[11] ;
 wire \u_reg.cfg_glb_ctrl[12] ;
 wire \u_reg.cfg_glb_ctrl[13] ;
 wire \u_reg.cfg_glb_ctrl[14] ;
 wire \u_reg.cfg_glb_ctrl[15] ;
 wire \u_reg.cfg_glb_ctrl[1] ;
 wire \u_reg.cfg_glb_ctrl[2] ;
 wire \u_reg.cfg_glb_ctrl[3] ;
 wire \u_reg.cfg_glb_ctrl[4] ;
 wire \u_reg.cfg_glb_ctrl[5] ;
 wire \u_reg.cfg_glb_ctrl[6] ;
 wire \u_reg.cfg_glb_ctrl[7] ;
 wire \u_reg.cfg_glb_ctrl[8] ;
 wire \u_reg.cfg_glb_ctrl[9] ;
 wire \u_reg.clk_enb ;
 wire \u_reg.cpu_clk_div ;
 wire \u_reg.cpu_ref_clk ;
 wire \u_reg.cpu_ref_clk_div_2 ;
 wire \u_reg.cpu_ref_clk_div_4 ;
 wire \u_reg.cpu_ref_clk_div_8 ;
 wire \u_reg.cpu_ref_clk_int ;
 wire \u_reg.force_refclk ;
 wire \u_reg.reg_ack ;
 wire \u_reg.reg_rdata[0] ;
 wire \u_reg.reg_rdata[10] ;
 wire \u_reg.reg_rdata[11] ;
 wire \u_reg.reg_rdata[12] ;
 wire \u_reg.reg_rdata[13] ;
 wire \u_reg.reg_rdata[14] ;
 wire \u_reg.reg_rdata[15] ;
 wire \u_reg.reg_rdata[16] ;
 wire \u_reg.reg_rdata[17] ;
 wire \u_reg.reg_rdata[18] ;
 wire \u_reg.reg_rdata[19] ;
 wire \u_reg.reg_rdata[1] ;
 wire \u_reg.reg_rdata[20] ;
 wire \u_reg.reg_rdata[21] ;
 wire \u_reg.reg_rdata[22] ;
 wire \u_reg.reg_rdata[23] ;
 wire \u_reg.reg_rdata[24] ;
 wire \u_reg.reg_rdata[25] ;
 wire \u_reg.reg_rdata[26] ;
 wire \u_reg.reg_rdata[27] ;
 wire \u_reg.reg_rdata[28] ;
 wire \u_reg.reg_rdata[29] ;
 wire \u_reg.reg_rdata[2] ;
 wire \u_reg.reg_rdata[30] ;
 wire \u_reg.reg_rdata[31] ;
 wire \u_reg.reg_rdata[3] ;
 wire \u_reg.reg_rdata[4] ;
 wire \u_reg.reg_rdata[5] ;
 wire \u_reg.reg_rdata[6] ;
 wire \u_reg.reg_rdata[7] ;
 wire \u_reg.reg_rdata[8] ;
 wire \u_reg.reg_rdata[9] ;
 wire \u_reg.soft_reboot ;
 wire \u_reg.u_bank_sel.gen_bit_reg[0].u_bit_reg.data_out ;
 wire \u_reg.u_bank_sel.gen_bit_reg[1].u_bit_reg.data_out ;
 wire \u_reg.u_bank_sel.gen_bit_reg[2].u_bit_reg.data_out ;
 wire \u_reg.u_buf_pll_rst.A ;
 wire \u_reg.u_buf_wb_rst.A ;
 wire \u_reg.u_clkgate_wbs.CLK ;
 wire \u_reg.u_wbclk.clk_div_2 ;
 wire \u_reg.u_wbclk.clk_div_4 ;
 wire \u_reg.u_wbclk.clk_div_8 ;
 wire \u_reg.u_wbclk.mclk ;
 wire \u_reg.u_wbs_ref_clkbuf.A ;
 wire \u_reset_fsm.boot_req_s ;
 wire \u_reset_fsm.boot_req_ss ;
 wire \u_reset_fsm.clk_cnt[0] ;
 wire \u_reset_fsm.clk_cnt[10] ;
 wire \u_reset_fsm.clk_cnt[11] ;
 wire \u_reset_fsm.clk_cnt[12] ;
 wire \u_reset_fsm.clk_cnt[13] ;
 wire \u_reset_fsm.clk_cnt[14] ;
 wire \u_reset_fsm.clk_cnt[15] ;
 wire \u_reset_fsm.clk_cnt[1] ;
 wire \u_reset_fsm.clk_cnt[2] ;
 wire \u_reset_fsm.clk_cnt[3] ;
 wire \u_reset_fsm.clk_cnt[4] ;
 wire \u_reset_fsm.clk_cnt[5] ;
 wire \u_reset_fsm.clk_cnt[6] ;
 wire \u_reset_fsm.clk_cnt[7] ;
 wire \u_reset_fsm.clk_cnt[8] ;
 wire \u_reset_fsm.clk_cnt[9] ;
 wire \u_reset_fsm.state[0] ;
 wire \u_reset_fsm.state[1] ;
 wire \u_reset_fsm.state[2] ;
 wire \u_skew_wh.clk_d1 ;
 wire \u_skew_wh.clk_d10 ;
 wire \u_skew_wh.clk_d11 ;
 wire \u_skew_wh.clk_d12 ;
 wire \u_skew_wh.clk_d13 ;
 wire \u_skew_wh.clk_d14 ;
 wire \u_skew_wh.clk_d15 ;
 wire \u_skew_wh.clk_d2 ;
 wire \u_skew_wh.clk_d3 ;
 wire \u_skew_wh.clk_d4 ;
 wire \u_skew_wh.clk_d5 ;
 wire \u_skew_wh.clk_d6 ;
 wire \u_skew_wh.clk_d7 ;
 wire \u_skew_wh.clk_d8 ;
 wire \u_skew_wh.clk_d9 ;
 wire \u_skew_wh.clk_inbuf ;
 wire \u_skew_wh.clkbuf_1.X1 ;
 wire \u_skew_wh.clkbuf_1.X2 ;
 wire \u_skew_wh.clkbuf_1.X3 ;
 wire \u_skew_wh.clkbuf_10.X1 ;
 wire \u_skew_wh.clkbuf_10.X2 ;
 wire \u_skew_wh.clkbuf_10.X3 ;
 wire \u_skew_wh.clkbuf_11.X1 ;
 wire \u_skew_wh.clkbuf_11.X2 ;
 wire \u_skew_wh.clkbuf_11.X3 ;
 wire \u_skew_wh.clkbuf_12.X1 ;
 wire \u_skew_wh.clkbuf_12.X2 ;
 wire \u_skew_wh.clkbuf_12.X3 ;
 wire \u_skew_wh.clkbuf_13.X1 ;
 wire \u_skew_wh.clkbuf_13.X2 ;
 wire \u_skew_wh.clkbuf_13.X3 ;
 wire \u_skew_wh.clkbuf_14.X1 ;
 wire \u_skew_wh.clkbuf_14.X2 ;
 wire \u_skew_wh.clkbuf_14.X3 ;
 wire \u_skew_wh.clkbuf_15.X1 ;
 wire \u_skew_wh.clkbuf_15.X2 ;
 wire \u_skew_wh.clkbuf_15.X3 ;
 wire \u_skew_wh.clkbuf_2.X1 ;
 wire \u_skew_wh.clkbuf_2.X2 ;
 wire \u_skew_wh.clkbuf_2.X3 ;
 wire \u_skew_wh.clkbuf_3.X1 ;
 wire \u_skew_wh.clkbuf_3.X2 ;
 wire \u_skew_wh.clkbuf_3.X3 ;
 wire \u_skew_wh.clkbuf_4.X1 ;
 wire \u_skew_wh.clkbuf_4.X2 ;
 wire \u_skew_wh.clkbuf_4.X3 ;
 wire \u_skew_wh.clkbuf_5.X1 ;
 wire \u_skew_wh.clkbuf_5.X2 ;
 wire \u_skew_wh.clkbuf_5.X3 ;
 wire \u_skew_wh.clkbuf_6.X1 ;
 wire \u_skew_wh.clkbuf_6.X2 ;
 wire \u_skew_wh.clkbuf_6.X3 ;
 wire \u_skew_wh.clkbuf_7.X1 ;
 wire \u_skew_wh.clkbuf_7.X2 ;
 wire \u_skew_wh.clkbuf_7.X3 ;
 wire \u_skew_wh.clkbuf_8.X1 ;
 wire \u_skew_wh.clkbuf_8.X2 ;
 wire \u_skew_wh.clkbuf_8.X3 ;
 wire \u_skew_wh.clkbuf_9.X1 ;
 wire \u_skew_wh.clkbuf_9.X2 ;
 wire \u_skew_wh.clkbuf_9.X3 ;
 wire \u_skew_wh.d00 ;
 wire \u_skew_wh.d01 ;
 wire \u_skew_wh.d02 ;
 wire \u_skew_wh.d03 ;
 wire \u_skew_wh.d04 ;
 wire \u_skew_wh.d05 ;
 wire \u_skew_wh.d06 ;
 wire \u_skew_wh.d07 ;
 wire \u_skew_wh.d10 ;
 wire \u_skew_wh.d11 ;
 wire \u_skew_wh.d12 ;
 wire \u_skew_wh.d13 ;
 wire \u_skew_wh.d20 ;
 wire \u_skew_wh.d21 ;
 wire \u_skew_wh.d30 ;
 wire \u_skew_wh.in0 ;
 wire \u_skew_wh.in1 ;
 wire \u_skew_wh.in10 ;
 wire \u_skew_wh.in11 ;
 wire \u_skew_wh.in12 ;
 wire \u_skew_wh.in13 ;
 wire \u_skew_wh.in14 ;
 wire \u_skew_wh.in15 ;
 wire \u_skew_wh.in2 ;
 wire \u_skew_wh.in3 ;
 wire \u_skew_wh.in4 ;
 wire \u_skew_wh.in5 ;
 wire \u_skew_wh.in6 ;
 wire \u_skew_wh.in7 ;
 wire \u_skew_wh.in8 ;
 wire \u_skew_wh.in9 ;
 wire \u_spi2wb.reg_addr[0] ;
 wire \u_spi2wb.reg_addr[10] ;
 wire \u_spi2wb.reg_addr[11] ;
 wire \u_spi2wb.reg_addr[12] ;
 wire \u_spi2wb.reg_addr[13] ;
 wire \u_spi2wb.reg_addr[14] ;
 wire \u_spi2wb.reg_addr[15] ;
 wire \u_spi2wb.reg_addr[16] ;
 wire \u_spi2wb.reg_addr[17] ;
 wire \u_spi2wb.reg_addr[18] ;
 wire \u_spi2wb.reg_addr[19] ;
 wire \u_spi2wb.reg_addr[1] ;
 wire \u_spi2wb.reg_addr[2] ;
 wire \u_spi2wb.reg_addr[3] ;
 wire \u_spi2wb.reg_addr[4] ;
 wire \u_spi2wb.reg_addr[5] ;
 wire \u_spi2wb.reg_addr[6] ;
 wire \u_spi2wb.reg_addr[7] ;
 wire \u_spi2wb.reg_addr[8] ;
 wire \u_spi2wb.reg_addr[9] ;
 wire \u_spi2wb.reg_be[0] ;
 wire \u_spi2wb.reg_be[1] ;
 wire \u_spi2wb.reg_be[2] ;
 wire \u_spi2wb.reg_be[3] ;
 wire \u_spi2wb.reg_rd ;
 wire \u_spi2wb.reg_wdata[0] ;
 wire \u_spi2wb.reg_wdata[10] ;
 wire \u_spi2wb.reg_wdata[11] ;
 wire \u_spi2wb.reg_wdata[12] ;
 wire \u_spi2wb.reg_wdata[13] ;
 wire \u_spi2wb.reg_wdata[14] ;
 wire \u_spi2wb.reg_wdata[15] ;
 wire \u_spi2wb.reg_wdata[16] ;
 wire \u_spi2wb.reg_wdata[17] ;
 wire \u_spi2wb.reg_wdata[18] ;
 wire \u_spi2wb.reg_wdata[19] ;
 wire \u_spi2wb.reg_wdata[1] ;
 wire \u_spi2wb.reg_wdata[20] ;
 wire \u_spi2wb.reg_wdata[21] ;
 wire \u_spi2wb.reg_wdata[22] ;
 wire \u_spi2wb.reg_wdata[23] ;
 wire \u_spi2wb.reg_wdata[24] ;
 wire \u_spi2wb.reg_wdata[25] ;
 wire \u_spi2wb.reg_wdata[26] ;
 wire \u_spi2wb.reg_wdata[27] ;
 wire \u_spi2wb.reg_wdata[28] ;
 wire \u_spi2wb.reg_wdata[29] ;
 wire \u_spi2wb.reg_wdata[2] ;
 wire \u_spi2wb.reg_wdata[30] ;
 wire \u_spi2wb.reg_wdata[31] ;
 wire \u_spi2wb.reg_wdata[3] ;
 wire \u_spi2wb.reg_wdata[4] ;
 wire \u_spi2wb.reg_wdata[5] ;
 wire \u_spi2wb.reg_wdata[6] ;
 wire \u_spi2wb.reg_wdata[7] ;
 wire \u_spi2wb.reg_wdata[8] ;
 wire \u_spi2wb.reg_wdata[9] ;
 wire \u_spi2wb.reg_wr ;
 wire \u_spi2wb.u_if.RegSdOut[0] ;
 wire \u_spi2wb.u_if.RegSdOut[10] ;
 wire \u_spi2wb.u_if.RegSdOut[11] ;
 wire \u_spi2wb.u_if.RegSdOut[12] ;
 wire \u_spi2wb.u_if.RegSdOut[13] ;
 wire \u_spi2wb.u_if.RegSdOut[14] ;
 wire \u_spi2wb.u_if.RegSdOut[15] ;
 wire \u_spi2wb.u_if.RegSdOut[16] ;
 wire \u_spi2wb.u_if.RegSdOut[17] ;
 wire \u_spi2wb.u_if.RegSdOut[18] ;
 wire \u_spi2wb.u_if.RegSdOut[19] ;
 wire \u_spi2wb.u_if.RegSdOut[1] ;
 wire \u_spi2wb.u_if.RegSdOut[20] ;
 wire \u_spi2wb.u_if.RegSdOut[21] ;
 wire \u_spi2wb.u_if.RegSdOut[22] ;
 wire \u_spi2wb.u_if.RegSdOut[23] ;
 wire \u_spi2wb.u_if.RegSdOut[24] ;
 wire \u_spi2wb.u_if.RegSdOut[25] ;
 wire \u_spi2wb.u_if.RegSdOut[26] ;
 wire \u_spi2wb.u_if.RegSdOut[27] ;
 wire \u_spi2wb.u_if.RegSdOut[28] ;
 wire \u_spi2wb.u_if.RegSdOut[29] ;
 wire \u_spi2wb.u_if.RegSdOut[2] ;
 wire \u_spi2wb.u_if.RegSdOut[30] ;
 wire \u_spi2wb.u_if.RegSdOut[31] ;
 wire \u_spi2wb.u_if.RegSdOut[3] ;
 wire \u_spi2wb.u_if.RegSdOut[4] ;
 wire \u_spi2wb.u_if.RegSdOut[5] ;
 wire \u_spi2wb.u_if.RegSdOut[6] ;
 wire \u_spi2wb.u_if.RegSdOut[7] ;
 wire \u_spi2wb.u_if.RegSdOut[8] ;
 wire \u_spi2wb.u_if.RegSdOut[9] ;
 wire \u_spi2wb.u_if.adr_phase ;
 wire \u_spi2wb.u_if.bitcnt[0] ;
 wire \u_spi2wb.u_if.bitcnt[1] ;
 wire \u_spi2wb.u_if.bitcnt[2] ;
 wire \u_spi2wb.u_if.bitcnt[3] ;
 wire \u_spi2wb.u_if.bitcnt[4] ;
 wire \u_spi2wb.u_if.bitcnt[5] ;
 wire \u_spi2wb.u_if.cmd_phase ;
 wire \u_spi2wb.u_if.cmd_reg[4] ;
 wire \u_spi2wb.u_if.cmd_reg[5] ;
 wire \u_spi2wb.u_if.cmd_reg[6] ;
 wire \u_spi2wb.u_if.cmd_reg[7] ;
 wire \u_spi2wb.u_if.rd_phase ;
 wire \u_spi2wb.u_if.sck_l0 ;
 wire \u_spi2wb.u_if.sck_l1 ;
 wire \u_spi2wb.u_if.sck_l2 ;
 wire \u_spi2wb.u_if.spi_if_st[0] ;
 wire \u_spi2wb.u_if.spi_if_st[1] ;
 wire \u_spi2wb.u_if.spi_if_st[5] ;
 wire \u_spi2wb.u_if.ssn_l0 ;
 wire \u_spi2wb.u_if.ssn_l1 ;
 wire \u_spi2wb.u_if.wr_phase ;
 wire \u_uart2wb.arst_ssn ;
 wire \u_uart2wb.auto_baud_16x[0] ;
 wire \u_uart2wb.auto_baud_16x[10] ;
 wire \u_uart2wb.auto_baud_16x[11] ;
 wire \u_uart2wb.auto_baud_16x[1] ;
 wire \u_uart2wb.auto_baud_16x[2] ;
 wire \u_uart2wb.auto_baud_16x[3] ;
 wire \u_uart2wb.auto_baud_16x[4] ;
 wire \u_uart2wb.auto_baud_16x[5] ;
 wire \u_uart2wb.auto_baud_16x[6] ;
 wire \u_uart2wb.auto_baud_16x[7] ;
 wire \u_uart2wb.auto_baud_16x[8] ;
 wire \u_uart2wb.auto_baud_16x[9] ;
 wire \u_uart2wb.auto_rx_enb ;
 wire \u_uart2wb.baud_clk_16x ;
 wire \u_uart2wb.line_reset_n ;
 wire \u_uart2wb.reg_ack ;
 wire \u_uart2wb.reg_addr[0] ;
 wire \u_uart2wb.reg_addr[10] ;
 wire \u_uart2wb.reg_addr[11] ;
 wire \u_uart2wb.reg_addr[12] ;
 wire \u_uart2wb.reg_addr[13] ;
 wire \u_uart2wb.reg_addr[14] ;
 wire \u_uart2wb.reg_addr[15] ;
 wire \u_uart2wb.reg_addr[16] ;
 wire \u_uart2wb.reg_addr[17] ;
 wire \u_uart2wb.reg_addr[18] ;
 wire \u_uart2wb.reg_addr[19] ;
 wire \u_uart2wb.reg_addr[1] ;
 wire \u_uart2wb.reg_addr[2] ;
 wire \u_uart2wb.reg_addr[3] ;
 wire \u_uart2wb.reg_addr[4] ;
 wire \u_uart2wb.reg_addr[5] ;
 wire \u_uart2wb.reg_addr[6] ;
 wire \u_uart2wb.reg_addr[7] ;
 wire \u_uart2wb.reg_addr[8] ;
 wire \u_uart2wb.reg_addr[9] ;
 wire \u_uart2wb.reg_rdata[0] ;
 wire \u_uart2wb.reg_rdata[10] ;
 wire \u_uart2wb.reg_rdata[11] ;
 wire \u_uart2wb.reg_rdata[12] ;
 wire \u_uart2wb.reg_rdata[13] ;
 wire \u_uart2wb.reg_rdata[14] ;
 wire \u_uart2wb.reg_rdata[15] ;
 wire \u_uart2wb.reg_rdata[16] ;
 wire \u_uart2wb.reg_rdata[17] ;
 wire \u_uart2wb.reg_rdata[18] ;
 wire \u_uart2wb.reg_rdata[19] ;
 wire \u_uart2wb.reg_rdata[1] ;
 wire \u_uart2wb.reg_rdata[20] ;
 wire \u_uart2wb.reg_rdata[21] ;
 wire \u_uart2wb.reg_rdata[22] ;
 wire \u_uart2wb.reg_rdata[23] ;
 wire \u_uart2wb.reg_rdata[24] ;
 wire \u_uart2wb.reg_rdata[25] ;
 wire \u_uart2wb.reg_rdata[26] ;
 wire \u_uart2wb.reg_rdata[27] ;
 wire \u_uart2wb.reg_rdata[28] ;
 wire \u_uart2wb.reg_rdata[29] ;
 wire \u_uart2wb.reg_rdata[2] ;
 wire \u_uart2wb.reg_rdata[30] ;
 wire \u_uart2wb.reg_rdata[31] ;
 wire \u_uart2wb.reg_rdata[3] ;
 wire \u_uart2wb.reg_rdata[4] ;
 wire \u_uart2wb.reg_rdata[5] ;
 wire \u_uart2wb.reg_rdata[6] ;
 wire \u_uart2wb.reg_rdata[7] ;
 wire \u_uart2wb.reg_rdata[8] ;
 wire \u_uart2wb.reg_rdata[9] ;
 wire \u_uart2wb.reg_req ;
 wire \u_uart2wb.reg_wdata[0] ;
 wire \u_uart2wb.reg_wdata[10] ;
 wire \u_uart2wb.reg_wdata[11] ;
 wire \u_uart2wb.reg_wdata[12] ;
 wire \u_uart2wb.reg_wdata[13] ;
 wire \u_uart2wb.reg_wdata[14] ;
 wire \u_uart2wb.reg_wdata[15] ;
 wire \u_uart2wb.reg_wdata[16] ;
 wire \u_uart2wb.reg_wdata[17] ;
 wire \u_uart2wb.reg_wdata[18] ;
 wire \u_uart2wb.reg_wdata[19] ;
 wire \u_uart2wb.reg_wdata[1] ;
 wire \u_uart2wb.reg_wdata[20] ;
 wire \u_uart2wb.reg_wdata[21] ;
 wire \u_uart2wb.reg_wdata[22] ;
 wire \u_uart2wb.reg_wdata[23] ;
 wire \u_uart2wb.reg_wdata[24] ;
 wire \u_uart2wb.reg_wdata[25] ;
 wire \u_uart2wb.reg_wdata[26] ;
 wire \u_uart2wb.reg_wdata[27] ;
 wire \u_uart2wb.reg_wdata[28] ;
 wire \u_uart2wb.reg_wdata[29] ;
 wire \u_uart2wb.reg_wdata[2] ;
 wire \u_uart2wb.reg_wdata[30] ;
 wire \u_uart2wb.reg_wdata[31] ;
 wire \u_uart2wb.reg_wdata[3] ;
 wire \u_uart2wb.reg_wdata[4] ;
 wire \u_uart2wb.reg_wdata[5] ;
 wire \u_uart2wb.reg_wdata[6] ;
 wire \u_uart2wb.reg_wdata[7] ;
 wire \u_uart2wb.reg_wdata[8] ;
 wire \u_uart2wb.reg_wdata[9] ;
 wire \u_uart2wb.reg_wr ;
 wire \u_uart2wb.rx_data[0] ;
 wire \u_uart2wb.rx_data[1] ;
 wire \u_uart2wb.rx_data[2] ;
 wire \u_uart2wb.rx_data[3] ;
 wire \u_uart2wb.rx_data[4] ;
 wire \u_uart2wb.rx_data[5] ;
 wire \u_uart2wb.rx_data[6] ;
 wire \u_uart2wb.rx_data[7] ;
 wire \u_uart2wb.rx_wr ;
 wire \u_uart2wb.tx_data[0] ;
 wire \u_uart2wb.tx_data[1] ;
 wire \u_uart2wb.tx_data[2] ;
 wire \u_uart2wb.tx_data[3] ;
 wire \u_uart2wb.tx_data[4] ;
 wire \u_uart2wb.tx_data[5] ;
 wire \u_uart2wb.tx_data[6] ;
 wire \u_uart2wb.tx_data_avail ;
 wire \u_uart2wb.tx_rd ;
 wire \u_uart2wb.u_arst_sync.in_data_2s ;
 wire \u_uart2wb.u_arst_sync.in_data_s ;
 wire \u_uart2wb.u_async_reg_bus.in_flag ;
 wire \u_uart2wb.u_async_reg_bus.in_flag_s ;
 wire \u_uart2wb.u_async_reg_bus.in_flag_ss ;
 wire \u_uart2wb.u_async_reg_bus.in_state[0] ;
 wire \u_uart2wb.u_async_reg_bus.in_state[1] ;
 wire \u_uart2wb.u_async_reg_bus.in_timer[0] ;
 wire \u_uart2wb.u_async_reg_bus.in_timer[1] ;
 wire \u_uart2wb.u_async_reg_bus.in_timer[2] ;
 wire \u_uart2wb.u_async_reg_bus.in_timer[3] ;
 wire \u_uart2wb.u_async_reg_bus.in_timer[4] ;
 wire \u_uart2wb.u_async_reg_bus.in_timer[5] ;
 wire \u_uart2wb.u_async_reg_bus.in_timer[6] ;
 wire \u_uart2wb.u_async_reg_bus.in_timer[7] ;
 wire \u_uart2wb.u_async_reg_bus.in_timer[8] ;
 wire \u_uart2wb.u_async_reg_bus.out_flag ;
 wire \u_uart2wb.u_async_reg_bus.out_flag_s ;
 wire \u_uart2wb.u_async_reg_bus.out_flag_ss ;
 wire \u_uart2wb.u_async_reg_bus.out_reg_cs ;
 wire \u_uart2wb.u_async_reg_bus.out_state[0] ;
 wire \u_uart2wb.u_async_reg_bus.out_state[1] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[0] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[10] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[11] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[12] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[13] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[14] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[15] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[16] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[17] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[18] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[19] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[1] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[2] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[3] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[4] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[5] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[6] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[7] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[8] ;
 wire \u_uart2wb.u_aut_det.clk_cnt[9] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[0] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[10] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[11] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[12] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[13] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[14] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[15] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[16] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[17] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[18] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[19] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[1] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[2] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[3] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[4] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[5] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[6] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[7] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[8] ;
 wire \u_uart2wb.u_aut_det.ref1_cnt[9] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[0] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[10] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[11] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[12] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[13] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[14] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[15] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[16] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[17] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[18] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[19] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[1] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[2] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[3] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[4] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[5] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[6] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[7] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[8] ;
 wire \u_uart2wb.u_aut_det.ref2_cnt[9] ;
 wire \u_uart2wb.u_aut_det.rxd_sync[0] ;
 wire \u_uart2wb.u_aut_det.rxd_sync[1] ;
 wire \u_uart2wb.u_aut_det.rxd_sync[2] ;
 wire \u_uart2wb.u_aut_det.state[0] ;
 wire \u_uart2wb.u_aut_det.state[1] ;
 wire \u_uart2wb.u_aut_det.state[2] ;
 wire \u_uart2wb.u_aut_det.state[3] ;
 wire \u_uart2wb.u_aut_det.state[4] ;
 wire \u_uart2wb.u_aut_det.state[5] ;
 wire \u_uart2wb.u_aut_det.state[6] ;
 wire \u_uart2wb.u_aut_det.state[7] ;
 wire \u_uart2wb.u_core.line_clk_16x ;
 wire \u_uart2wb.u_core.si_ss ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[0] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[10] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[11] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[1] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[2] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[3] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[4] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[5] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[6] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[7] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[8] ;
 wire \u_uart2wb.u_core.u_clk_ctl.high_count[9] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[0] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[10] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[11] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[1] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[2] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[3] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[4] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[5] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[6] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[7] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[8] ;
 wire \u_uart2wb.u_core.u_clk_ctl.low_count[9] ;
 wire \u_uart2wb.u_core.u_line_rst.in_data_2s ;
 wire \u_uart2wb.u_core.u_line_rst.in_data_s ;
 wire \u_uart2wb.u_core.u_rxd_sync.in_data_2s ;
 wire \u_uart2wb.u_core.u_rxd_sync.in_data_s ;
 wire \u_uart2wb.u_core.u_rxfsm.cnt[0] ;
 wire \u_uart2wb.u_core.u_rxfsm.cnt[1] ;
 wire \u_uart2wb.u_core.u_rxfsm.cnt[2] ;
 wire \u_uart2wb.u_core.u_rxfsm.offset[0] ;
 wire \u_uart2wb.u_core.u_rxfsm.offset[1] ;
 wire \u_uart2wb.u_core.u_rxfsm.offset[2] ;
 wire \u_uart2wb.u_core.u_rxfsm.offset[3] ;
 wire \u_uart2wb.u_core.u_rxfsm.rxpos[0] ;
 wire \u_uart2wb.u_core.u_rxfsm.rxpos[1] ;
 wire \u_uart2wb.u_core.u_rxfsm.rxpos[2] ;
 wire \u_uart2wb.u_core.u_rxfsm.rxpos[3] ;
 wire \u_uart2wb.u_core.u_rxfsm.rxstate[0] ;
 wire \u_uart2wb.u_core.u_rxfsm.rxstate[1] ;
 wire \u_uart2wb.u_core.u_rxfsm.rxstate[2] ;
 wire \u_uart2wb.u_core.u_txfsm.cnt[0] ;
 wire \u_uart2wb.u_core.u_txfsm.cnt[1] ;
 wire \u_uart2wb.u_core.u_txfsm.cnt[2] ;
 wire \u_uart2wb.u_core.u_txfsm.divcnt[0] ;
 wire \u_uart2wb.u_core.u_txfsm.divcnt[1] ;
 wire \u_uart2wb.u_core.u_txfsm.divcnt[2] ;
 wire \u_uart2wb.u_core.u_txfsm.divcnt[3] ;
 wire \u_uart2wb.u_core.u_txfsm.txdata[0] ;
 wire \u_uart2wb.u_core.u_txfsm.txdata[1] ;
 wire \u_uart2wb.u_core.u_txfsm.txdata[2] ;
 wire \u_uart2wb.u_core.u_txfsm.txdata[3] ;
 wire \u_uart2wb.u_core.u_txfsm.txdata[4] ;
 wire \u_uart2wb.u_core.u_txfsm.txdata[5] ;
 wire \u_uart2wb.u_core.u_txfsm.txdata[6] ;
 wire \u_uart2wb.u_core.u_txfsm.txstate[0] ;
 wire \u_uart2wb.u_core.u_txfsm.txstate[1] ;
 wire \u_uart2wb.u_core.u_txfsm.txstate[2] ;
 wire \u_uart2wb.u_core.u_txfsm.txstate[3] ;
 wire \u_uart2wb.u_core.u_txfsm.txstate[4] ;
 wire \u_uart2wb.u_msg.NextState[0] ;
 wire \u_uart2wb.u_msg.NextState[1] ;
 wire \u_uart2wb.u_msg.NextState[2] ;
 wire \u_uart2wb.u_msg.NextState[3] ;
 wire \u_uart2wb.u_msg.RxMsgCnt[0] ;
 wire \u_uart2wb.u_msg.RxMsgCnt[1] ;
 wire \u_uart2wb.u_msg.RxMsgCnt[2] ;
 wire \u_uart2wb.u_msg.RxMsgCnt[3] ;
 wire \u_uart2wb.u_msg.RxMsgCnt[4] ;
 wire \u_uart2wb.u_msg.State[0] ;
 wire \u_uart2wb.u_msg.State[1] ;
 wire \u_uart2wb.u_msg.State[2] ;
 wire \u_uart2wb.u_msg.State[3] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[100] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[101] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[102] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[104] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[105] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[106] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[107] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[108] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[109] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[110] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[112] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[113] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[114] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[115] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[116] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[117] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[118] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[11] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[120] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[121] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[122] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[123] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[124] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[125] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[126] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[12] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[13] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[17] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[18] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[20] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[21] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[24] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[25] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[26] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[28] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[29] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[32] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[33] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[34] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[35] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[36] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[37] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[38] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[40] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[41] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[42] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[43] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[44] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[45] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[46] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[48] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[49] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[50] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[51] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[52] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[53] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[54] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[56] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[57] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[58] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[59] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[5] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[60] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[61] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[62] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[64] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[65] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[66] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[67] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[68] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[69] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[70] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[72] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[73] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[74] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[75] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[76] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[77] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[78] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[80] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[81] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[82] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[83] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[84] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[85] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[86] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[88] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[89] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[90] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[91] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[92] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[93] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[94] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[96] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[97] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[98] ;
 wire \u_uart2wb.u_msg.TxMsgBuf[99] ;
 wire \u_uart2wb.u_msg.TxMsgSize[0] ;
 wire \u_uart2wb.u_msg.TxMsgSize[1] ;
 wire \u_uart2wb.u_msg.TxMsgSize[2] ;
 wire \u_uart2wb.u_msg.TxMsgSize[3] ;
 wire \u_uart2wb.u_msg.TxMsgSize[4] ;
 wire \u_uart2wb.u_msg.cmd[0] ;
 wire \u_uart2wb.u_msg.cmd[10] ;
 wire \u_uart2wb.u_msg.cmd[11] ;
 wire \u_uart2wb.u_msg.cmd[12] ;
 wire \u_uart2wb.u_msg.cmd[13] ;
 wire \u_uart2wb.u_msg.cmd[14] ;
 wire \u_uart2wb.u_msg.cmd[15] ;
 wire \u_uart2wb.u_msg.cmd[1] ;
 wire \u_uart2wb.u_msg.cmd[2] ;
 wire \u_uart2wb.u_msg.cmd[3] ;
 wire \u_uart2wb.u_msg.cmd[4] ;
 wire \u_uart2wb.u_msg.cmd[5] ;
 wire \u_uart2wb.u_msg.cmd[6] ;
 wire \u_uart2wb.u_msg.cmd[7] ;
 wire \u_uart2wb.u_msg.cmd[8] ;
 wire \u_uart2wb.u_msg.cmd[9] ;
 wire \u_uart2wb.u_msg.wait_cnt[0] ;
 wire \u_uart2wb.u_msg.wait_cnt[1] ;
 wire \u_uart2wb.u_msg.wait_cnt[2] ;
 wire \u_uart2wb.u_msg.wait_cnt[3] ;
 wire \u_uart2wb.u_msg.wait_cnt[4] ;
 wire \u_uart2wb.u_msg.wait_cnt[5] ;
 wire \u_uart2wb.u_msg.wait_cnt[6] ;
 wire \u_uart2wb.u_msg.wait_cnt[7] ;
 wire \u_wbm_rst.arst_n ;
 wire \u_wbm_rst.in_data_2s ;
 wire \u_wbm_rst.in_data_s ;
 wire \u_wbs_rst.in_data_2s ;
 wire \u_wbs_rst.in_data_s ;
 wire wb_ack_o;
 wire wb_ack_o1;
 wire \wb_dat_o[0] ;
 wire \wb_dat_o[10] ;
 wire \wb_dat_o[11] ;
 wire \wb_dat_o[12] ;
 wire \wb_dat_o[13] ;
 wire \wb_dat_o[14] ;
 wire \wb_dat_o[15] ;
 wire \wb_dat_o[16] ;
 wire \wb_dat_o[17] ;
 wire \wb_dat_o[18] ;
 wire \wb_dat_o[19] ;
 wire \wb_dat_o[1] ;
 wire \wb_dat_o[20] ;
 wire \wb_dat_o[21] ;
 wire \wb_dat_o[22] ;
 wire \wb_dat_o[23] ;
 wire \wb_dat_o[24] ;
 wire \wb_dat_o[25] ;
 wire \wb_dat_o[26] ;
 wire \wb_dat_o[27] ;
 wire \wb_dat_o[28] ;
 wire \wb_dat_o[29] ;
 wire \wb_dat_o[2] ;
 wire \wb_dat_o[30] ;
 wire \wb_dat_o[31] ;
 wire \wb_dat_o[3] ;
 wire \wb_dat_o[4] ;
 wire \wb_dat_o[5] ;
 wire \wb_dat_o[6] ;
 wire \wb_dat_o[7] ;
 wire \wb_dat_o[8] ;
 wire \wb_dat_o[9] ;
 wire wb_err_o;
 wire wb_err_o1;
 wire wb_req;

 sky130_fd_sc_hd__diode_2 ANTENNA__04633__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__04635__A (.DIODE(_01107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04638__A (.DIODE(\u_spi2wb.u_if.ssn_l1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04642__B_N (.DIODE(\u_spi2wb.u_if.sck_l1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04658__B (.DIODE(\u_spi2wb.u_if.sck_l1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04674__A (.DIODE(strap_uartm[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__04675__A (.DIODE(strap_uartm[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__04678__A (.DIODE(la_data_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__04678__B (.DIODE(la_data_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__04681__B2 (.DIODE(_01149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04684__A (.DIODE(strap_uartm[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__04689__A1 (.DIODE(la_data_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__04689__A2 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04689__B1 (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04689__B2 (.DIODE(\u_uart2wb.auto_rx_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04691__A (.DIODE(\u_uart2wb.tx_data_avail ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04696__A (.DIODE(la_data_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__04696__B (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04697__B (.DIODE(_01163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04715__B1 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04718__B (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04721__A1 (.DIODE(\u_uart2wb.tx_data_avail ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04723__A2 (.DIODE(_01163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04975__B (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04988__A1 (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04994__A (.DIODE(\u_spi2wb.u_if.ssn_l1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05004__A (.DIODE(\u_spi2wb.u_if.ssn_l1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05017__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05019__A (.DIODE(wbm_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__05024__A (.DIODE(wbm_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05026__A (.DIODE(wb_req));
 sky130_fd_sc_hd__diode_2 ANTENNA__05026__B (.DIODE(_01476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05032__A2 (.DIODE(\u_spi2wb.reg_wr ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05032__B1 (.DIODE(wbm_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__05034__A (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05035__A (.DIODE(wb_req));
 sky130_fd_sc_hd__diode_2 ANTENNA__05036__B (.DIODE(_01476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05042__B (.DIODE(\u_async_wb.u_cmd_if.grey_wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05051__A (.DIODE(_01485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05057__A (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05057__C (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05059__A1 (.DIODE(_01479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05063__A (.DIODE(_01511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05063__B (.DIODE(wb_ack_o1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05064__A0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__05064__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__05064__A2 (.DIODE(int_pll_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__05064__A3 (.DIODE(xtal_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__05064__S0 (.DIODE(\u_reg.cfg_clk_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05064__S1 (.DIODE(\u_reg.cfg_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05066__A (.DIODE(\u_reg.cfg_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05067__S (.DIODE(\u_reg.cfg_clk_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05069__A (.DIODE(\u_reg.cfg_clk_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05074__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__05075__A0 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__05075__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__05075__A2 (.DIODE(int_pll_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA__05075__A3 (.DIODE(xtal_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__05075__S0 (.DIODE(\u_reg.cfg_clk_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05075__S1 (.DIODE(\u_reg.cfg_clk_ctrl[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05079__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05081__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05083__A (.DIODE(_01526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05086__A (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05087__A (.DIODE(_01530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05088__S0 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05088__S1 (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05091__S0 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05091__S1 (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05095__S1 (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05098__A (.DIODE(_01530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05102__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05108__A (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05109__A (.DIODE(_01526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05110__A (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05115__A (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05116__A (.DIODE(_01552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05117__A (.DIODE(_01553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05121__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05123__B (.DIODE(_01558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05126__B (.DIODE(_01560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05129__S0 (.DIODE(_01562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05130__B (.DIODE(_01563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05132__A (.DIODE(_01553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05133__S0 (.DIODE(_01562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05136__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05137__S0 (.DIODE(_01562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05138__B (.DIODE(_01569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05139__A (.DIODE(_01570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05140__S0 (.DIODE(_01562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05141__B (.DIODE(_01571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05142__A (.DIODE(_01572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05145__B (.DIODE(_01574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05146__A (.DIODE(_01575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05147__A (.DIODE(_01553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05149__B (.DIODE(_01577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05150__A (.DIODE(_01578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05152__A (.DIODE(_01579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05154__B (.DIODE(_01581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05157__B (.DIODE(_01583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05160__S0 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05161__B (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05163__A (.DIODE(_01553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05164__S0 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05165__B (.DIODE(_01589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05167__A (.DIODE(_01579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05168__S0 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05171__S0 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05174__A (.DIODE(_01526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05179__A (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05184__A (.DIODE(_01579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05199__A (.DIODE(_01579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05237__A (.DIODE(_01526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05242__A (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05245__B (.DIODE(_01649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05252__B (.DIODE(_01654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05256__B (.DIODE(_01657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05260__B (.DIODE(_01660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05264__B (.DIODE(_01663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05267__B (.DIODE(_01665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05271__B (.DIODE(_01668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05275__B (.DIODE(_01671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05277__A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05296__A (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05299__A (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05300__A (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05303__A (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05304__A (.DIODE(_01552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05307__A (.DIODE(_01695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05311__A (.DIODE(_01698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05314__A (.DIODE(_01700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05315__A (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05318__A (.DIODE(_01703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05319__A (.DIODE(_01552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05326__A (.DIODE(_01709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05330__A (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05333__A (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05334__A (.DIODE(_01552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05337__A (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05340__B (.DIODE(_01719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05343__B (.DIODE(_01721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05346__B (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05348__S1 (.DIODE(_01530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05349__B (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05357__A (.DIODE(\u_spi2wb.reg_wr ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05357__B (.DIODE(\u_spi2wb.reg_rd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05365__A1 (.DIODE(wbm_cyc_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__05365__A2 (.DIODE(wbm_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__05365__A3 (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05365__B1 (.DIODE(_01739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05366__A1 (.DIODE(_01731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05367__A (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05370__A (.DIODE(\wb_dat_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05372__A (.DIODE(\wb_dat_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05374__A (.DIODE(\wb_dat_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05376__A (.DIODE(\wb_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05379__A (.DIODE(\wb_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05381__A (.DIODE(\wb_dat_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05383__A (.DIODE(\wb_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05385__A (.DIODE(\wb_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05389__A (.DIODE(\wb_dat_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05391__A (.DIODE(\wb_dat_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05393__A (.DIODE(\wb_dat_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05395__A (.DIODE(\wb_dat_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05398__A (.DIODE(\wb_dat_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05400__A (.DIODE(\wb_dat_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05402__A (.DIODE(\wb_dat_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05404__A (.DIODE(\wb_dat_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05407__A (.DIODE(\wb_dat_o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05409__A (.DIODE(\wb_dat_o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05411__A (.DIODE(\wb_dat_o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05413__A (.DIODE(\wb_dat_o[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05416__A (.DIODE(\wb_dat_o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05418__A (.DIODE(\wb_dat_o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05420__A (.DIODE(\wb_dat_o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05422__A (.DIODE(\wb_dat_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05426__A (.DIODE(_01775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05428__A (.DIODE(\wb_dat_o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05430__A (.DIODE(\wb_dat_o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05432__A (.DIODE(\wb_dat_o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05434__A (.DIODE(\wb_dat_o[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05437__A (.DIODE(\wb_dat_o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05439__A (.DIODE(\wb_dat_o[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05441__A (.DIODE(\wb_dat_o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05443__A (.DIODE(\wb_dat_o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05446__A (.DIODE(_01787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05454__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__05456__A (.DIODE(_01794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05458__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__05462__A (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05462__B (.DIODE(\u_reg.cfg_glb_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05488__A (.DIODE(_01511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05513__A (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05515__B2 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05516__C_N (.DIODE(\u_spi2wb.reg_rd ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05520__A0 (.DIODE(\wb_dat_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05520__A1 (.DIODE(_01841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05520__S (.DIODE(wb_ack_o1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05526__A0 (.DIODE(\u_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05527__A0 (.DIODE(\wb_dat_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05527__A1 (.DIODE(_01847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05527__S (.DIODE(wb_ack_o1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05532__A0 (.DIODE(\wb_dat_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05532__A1 (.DIODE(_01850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05535__A (.DIODE(_01787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05537__A0 (.DIODE(\wb_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05541__A0 (.DIODE(\wb_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05541__A1 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05546__A0 (.DIODE(\wb_dat_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05546__A1 (.DIODE(_01862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05552__A0 (.DIODE(\wb_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05552__A1 (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05555__A (.DIODE(_01787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05557__A0 (.DIODE(\wb_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05557__A1 (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05561__A0 (.DIODE(\wb_dat_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05561__A1 (.DIODE(_01874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05566__A0 (.DIODE(\wb_dat_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05566__A1 (.DIODE(_01878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05571__A0 (.DIODE(\wb_dat_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05571__A1 (.DIODE(_01881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05574__A (.DIODE(_01479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05576__A1 (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05576__S (.DIODE(_01886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05577__A0 (.DIODE(\wb_dat_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05577__A1 (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05580__S (.DIODE(_01886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05581__A0 (.DIODE(\wb_dat_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05581__A1 (.DIODE(_01890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05585__S (.DIODE(_01886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05586__A0 (.DIODE(\wb_dat_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05586__A1 (.DIODE(_01894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05589__S (.DIODE(_01886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05591__A0 (.DIODE(\wb_dat_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05591__A1 (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05596__A0 (.DIODE(\wb_dat_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05596__A1 (.DIODE(_01902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05600__A0 (.DIODE(\wb_dat_o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05600__A1 (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05605__A0 (.DIODE(\wb_dat_o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05605__A1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05610__A0 (.DIODE(\wb_dat_o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05610__A1 (.DIODE(_01912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05615__A0 (.DIODE(\wb_dat_o[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05615__A1 (.DIODE(_01917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05619__A0 (.DIODE(\wb_dat_o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05619__A1 (.DIODE(_01920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05624__A0 (.DIODE(\wb_dat_o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05624__A1 (.DIODE(_01924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05629__A0 (.DIODE(\wb_dat_o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05629__A1 (.DIODE(_01927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05634__A0 (.DIODE(\wb_dat_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05638__A0 (.DIODE(\wb_dat_o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05642__A0 (.DIODE(\u_reg.reg_rdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05643__A0 (.DIODE(\wb_dat_o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05648__A0 (.DIODE(\wb_dat_o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05651__A (.DIODE(_01479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05652__A0 (.DIODE(\u_reg.reg_rdata[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05653__A0 (.DIODE(\wb_dat_o[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05656__A0 (.DIODE(\u_reg.reg_rdata[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05657__A0 (.DIODE(\wb_dat_o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05661__A0 (.DIODE(\wb_dat_o[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05665__A0 (.DIODE(\wb_dat_o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05668__S (.DIODE(_01787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05669__A0 (.DIODE(\wb_dat_o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05688__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__05690__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__05775__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05776__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05782__A0 (.DIODE(\u_spi2wb.reg_be[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05784__A (.DIODE(_02048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05785__A1 (.DIODE(\u_spi2wb.reg_be[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05794__A (.DIODE(_02059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05796__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05831__A (.DIODE(_02059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05841__A (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05843__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05878__A (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05939__A0 (.DIODE(_01794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05941__B1 (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05946__A (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05947__A1 (.DIODE(wbm_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05947__A2 (.DIODE(_01775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05948__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__05952__B2 (.DIODE(wbm_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05953__A (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05954__B1 (.DIODE(wbm_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05956__A (.DIODE(_02161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05958__A1 (.DIODE(wbm_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05959__A (.DIODE(_02164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05960__B1 (.DIODE(wbm_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05962__A (.DIODE(_02167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05964__C_N (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05966__A (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05966__B (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05968__A0 (.DIODE(\u_reg.cfg_glb_ctrl[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05973__B1 (.DIODE(wbm_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05975__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__05977__A1 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05980__B1 (.DIODE(wbm_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05982__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__05984__A1 (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05986__A (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05987__A1 (.DIODE(wbm_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05987__A2 (.DIODE(_01775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05988__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__05996__A1 (.DIODE(wbm_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__05997__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__06003__A1 (.DIODE(wbm_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06004__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06008__B1 (.DIODE(wbm_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06010__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__06015__A (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06016__A1 (.DIODE(wbm_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06016__A2 (.DIODE(_02213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06017__A (.DIODE(_02215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06021__A (.DIODE(wb_req));
 sky130_fd_sc_hd__diode_2 ANTENNA__06021__B (.DIODE(_01476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06023__B (.DIODE(_01485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06023__C (.DIODE(_02220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06024__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06027__A (.DIODE(\u_async_wb.m_cmd_wr_data[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06029__A1 (.DIODE(wbm_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06030__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__06032__A1 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06034__A (.DIODE(\u_async_wb.m_cmd_wr_data[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06036__A1 (.DIODE(wbm_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06036__A2 (.DIODE(_02213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06037__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__06038__A1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06040__A (.DIODE(\u_async_wb.m_cmd_wr_data[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06042__A1 (.DIODE(wbm_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06043__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06044__A (.DIODE(_02238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06047__A (.DIODE(\u_async_wb.m_cmd_wr_data[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06050__A1 (.DIODE(wbm_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06051__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__06053__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06054__A1 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06054__S (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06056__A (.DIODE(\u_async_wb.m_cmd_wr_data[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06058__B1 (.DIODE(wbm_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06060__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__06062__A1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06062__S (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06064__B1 (.DIODE(wbm_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06066__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__06068__A1 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06068__S (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06073__A1 (.DIODE(wbm_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06074__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06076__A1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06076__S (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06079__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06088__A (.DIODE(\u_async_wb.m_cmd_wr_data[65] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06092__A (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06093__S (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06095__A (.DIODE(\u_async_wb.m_cmd_wr_data[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06096__S (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06100__A1 (.DIODE(wbm_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06101__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__06103__A1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06103__S (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06105__A_N (.DIODE(_02164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06105__B (.DIODE(_02167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06105__C (.DIODE(_02161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06106__B (.DIODE(_01484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06106__C (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06107__A (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06109__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__06109__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__06110__A0 (.DIODE(strap_sticky[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06110__S (.DIODE(_01794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06112__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__06112__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06113__A0 (.DIODE(strap_sticky[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06113__S (.DIODE(_01794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06115__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__06117__A0 (.DIODE(strap_sticky[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06119__A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__06119__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__06120__A0 (.DIODE(strap_sticky[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06123__A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__06123__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__06124__A0 (.DIODE(strap_sticky[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06126__A0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__06126__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06127__A0 (.DIODE(strap_sticky[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06129__A0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__06129__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__06130__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06132__A0 (.DIODE(strap_sticky[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06134__A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__06134__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__06135__A0 (.DIODE(strap_sticky[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06138__A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__06138__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__06139__A0 (.DIODE(strap_sticky[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06141__A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__06141__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__06142__A0 (.DIODE(strap_sticky[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06144__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__06144__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__06146__A0 (.DIODE(strap_sticky[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06148__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__06148__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__06149__A0 (.DIODE(strap_sticky[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06152__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__06152__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__06153__A0 (.DIODE(strap_sticky[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06155__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__06155__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06156__A0 (.DIODE(strap_sticky[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06158__A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__06160__A0 (.DIODE(strap_sticky[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__A1 (.DIODE(_02215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06163__A0 (.DIODE(strap_sticky[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06166__A1 (.DIODE(wbm_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06167__A (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06169__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__06169__A1 (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06170__A0 (.DIODE(strap_sticky[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06174__A1 (.DIODE(wbm_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06175__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__06175__A1 (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06176__A0 (.DIODE(strap_sticky[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06180__A1 (.DIODE(wbm_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06181__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__06181__A1 (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06183__A0 (.DIODE(strap_sticky[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06186__B1 (.DIODE(wbm_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06188__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__06188__A1 (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06189__A0 (.DIODE(strap_sticky[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06191__B1 (.DIODE(wbm_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06194__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__06194__A1 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06195__A0 (.DIODE(strap_sticky[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06198__A1 (.DIODE(wbm_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06199__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__06199__A1 (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06200__A0 (.DIODE(strap_sticky[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06202__B1 (.DIODE(wbm_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06204__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__06204__A1 (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06205__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06206__A0 (.DIODE(strap_sticky[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06209__A1 (.DIODE(wbm_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06210__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__06210__A1 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06211__A0 (.DIODE(strap_sticky[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06214__B1 (.DIODE(wbm_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06217__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__06217__A1 (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06218__A0 (.DIODE(strap_sticky[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06221__B1 (.DIODE(wbm_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06223__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__06223__A1 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06224__A0 (.DIODE(strap_sticky[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06227__B1 (.DIODE(wbm_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06229__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__06229__A1 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06230__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06231__A0 (.DIODE(strap_sticky[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06234__A1 (.DIODE(wbm_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06234__A2 (.DIODE(_02213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06234__B1 (.DIODE(_01739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06235__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__06235__A1 (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06236__A0 (.DIODE(strap_sticky[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06238__B1 (.DIODE(wbm_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06241__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__06241__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06242__A0 (.DIODE(strap_sticky[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06245__A1 (.DIODE(wbm_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06245__A2 (.DIODE(_02213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06245__B1 (.DIODE(_01739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06246__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__06246__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__A0 (.DIODE(strap_sticky[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06249__B1 (.DIODE(wbm_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06251__A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__06251__A1 (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06252__A0 (.DIODE(strap_sticky[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06254__A1 (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06254__B1 (.DIODE(wbm_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06259__A (.DIODE(\u_async_wb.m_cmd_wr_data[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06260__S (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06262__A (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06265__B2 (.DIODE(wbm_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06266__B (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06266__C (.DIODE(_02415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06267__A (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06268__A1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06268__A2 (.DIODE(_02415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06268__B1 (.DIODE(_01107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06269__A (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06271__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06272__B (.DIODE(strap_sticky[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06273__A1 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06273__B2 (.DIODE(\u_reg.cfg_clk_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06274__A (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06276__B (.DIODE(strap_sticky[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06277__A1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06277__B2 (.DIODE(\u_reg.cfg_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06278__A (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06280__B (.DIODE(strap_sticky[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06281__A1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06282__A (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06284__B (.DIODE(strap_sticky[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06285__A1 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06286__A (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06288__A (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06289__A (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06290__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06291__B (.DIODE(strap_sticky[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06292__A1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06292__B2 (.DIODE(\u_reg.cfg_clk_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06293__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06295__B (.DIODE(strap_sticky[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06296__A1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06296__B2 (.DIODE(\u_reg.cfg_clk_ctrl[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06297__A (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06299__B (.DIODE(strap_sticky[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06300__A1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06301__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06303__B (.DIODE(strap_sticky[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06304__A1 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06305__A_N (.DIODE(_02167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06305__B (.DIODE(_02164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06305__C (.DIODE(_02161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06306__B (.DIODE(_01485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06306__C (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06309__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__06309__S (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06310__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__06313__A (.DIODE(_01479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06313__B (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06313__C_N (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06315__A (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06317__A (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06318__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__06321__A1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06322__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__06322__S (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06323__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__06325__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__06325__S (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06326__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__06328__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06329__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06331__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__06334__A1 (.DIODE(_02238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06337__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__06339__A1 (.DIODE(_02473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06340__A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__06340__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__06343__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__06345__A1 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06346__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__06349__A (.DIODE(_01107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06351__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__06354__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__06355__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__06356__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06357__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__06360__A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__06363__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__06363__A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__06366__A (.DIODE(_02215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06367__A (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06368__A (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06372__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__06373__A1 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06374__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__06375__A1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06376__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__06377__A1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06378__A (.DIODE(_01107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06380__A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__06380__S (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06381__A (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06383__A (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06384__A (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06385__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__06387__A1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06388__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__06389__A1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06390__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__06391__A1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06392__A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__06392__S (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06393__A (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06395__A (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06396__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__06397__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06398__A (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06400__A (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06401__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__06404__A1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06405__A (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06406__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__06407__A1 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06408__A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__06408__A1 (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06408__S (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06409__A (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06411__A (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06412__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__06413__A1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06414__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06414__S (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06415__A (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06417__A (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06418__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__06419__A1 (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06420__A (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06421__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__06421__B (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06422__A1 (.DIODE(_02531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06422__A2 (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06422__C1 (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06423__B (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06427__A (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06430__B (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06431__A (.DIODE(_02540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06433__A (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06434__A (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06436__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06438__A (.DIODE(_02220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06439__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06440__B1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06441__B1 (.DIODE(_02547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__C1 (.DIODE(_02551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06446__A (.DIODE(_02540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__06448__A (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06449__A (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06450__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06452__A1 (.DIODE(\u_reg.cfg_glb_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06452__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__06454__A (.DIODE(_02547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06455__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__06458__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06458__A3 (.DIODE(_02564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06458__B2 (.DIODE(\u_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06461__A (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06462__B1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06463__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__06467__B1 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06468__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__06470__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06470__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__06471__A2 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06471__A3 (.DIODE(_02577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06472__A (.DIODE(_02547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06473__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06473__B1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06474__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__06475__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__06476__B1 (.DIODE(_02580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06477__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06477__B1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06478__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__06479__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__06480__B1 (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06481__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__A (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__A2 (.DIODE(_02588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__A3 (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__06489__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__06490__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__06491__B1 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06492__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__06498__A1 (.DIODE(\u_reg.cfg_glb_ctrl[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06499__A2 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06499__A3 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06500__B2 (.DIODE(\u_async_wb.m_cmd_wr_data[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06503__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__06504__B1 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06505__A2 (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06505__B2 (.DIODE(\u_async_wb.m_cmd_wr_data[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__B1 (.DIODE(_02606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06510__A (.DIODE(_02540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06511__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__06513__A (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06514__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__06514__A2 (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06514__B1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06517__A3 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06518__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__06519__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[65] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__A3 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06522__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__06523__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__06523__A2 (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06523__B1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06525__A3 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__A2 (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__06529__B1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06530__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__06531__A2 (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06531__B1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06533__A2 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06533__A3 (.DIODE(_02627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06534__A (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__A1 (.DIODE(\u_reg.cfg_clk_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__A2 (.DIODE(_02557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__B1 (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__B2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__06536__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__06536__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__06539__A (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__A1 (.DIODE(\u_reg.cfg_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__B1 (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__B2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__06541__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__06541__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__06544__A (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06545__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__A1 (.DIODE(\u_reg.cfg_clk_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__A (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06552__A1 (.DIODE(\u_reg.cfg_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06552__B2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__06553__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__06553__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__06556__A1 (.DIODE(\u_reg.cfg_clk_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06556__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__06557__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__06557__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__06560__A1 (.DIODE(\u_reg.cfg_clk_ctrl[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06560__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06560__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__06564__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06564__B2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__06565__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__06565__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__06569__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__06569__B1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06569__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__06574__A (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06575__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__06575__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__A (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__06579__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__A1 (.DIODE(\u_reg.reg_rdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__B2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__A (.DIODE(_02547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06589__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__06589__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__06591__A1 (.DIODE(\u_reg.reg_rdata[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__06594__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__06594__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__06595__A1 (.DIODE(\u_reg.reg_rdata[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06596__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__06596__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__06603__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__06605__A (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06612__B (.DIODE(strap_sticky[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06613__A2 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06613__B2 (.DIODE(strap_sticky[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06614__C_N (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06615__B (.DIODE(_02690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06617__A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__06619__B (.DIODE(_02690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__B (.DIODE(_02690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__B2 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06625__B (.DIODE(_02690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__B (.DIODE(strap_sticky[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__C_N (.DIODE(strap_sticky[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__B2 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06629__B (.DIODE(strap_sticky[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06630__A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06630__B2 (.DIODE(strap_sticky[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06631__A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__06633__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__06633__B2 (.DIODE(_02473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06634__B (.DIODE(strap_sticky[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06634__C_N (.DIODE(strap_sticky[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__B2 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06639__A (.DIODE(strap_sticky[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06640__B (.DIODE(strap_sticky[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06642__B2 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06643__B2 (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06648__C_N (.DIODE(strap_sticky[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06649__B2 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06650__B (.DIODE(strap_sticky[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06651__A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06651__B2 (.DIODE(strap_sticky[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06655__A (.DIODE(strap_sticky[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06656__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06656__C (.DIODE(strap_sticky[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06658__A (.DIODE(strap_sticky[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06659__A2 (.DIODE(strap_sticky[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06659__B1 (.DIODE(_01799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__B2 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__A1 (.DIODE(strap_sticky[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__A2 (.DIODE(strap_sticky[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__B1 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06662__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__06662__B2 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A1 (.DIODE(strap_sticky[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A2 (.DIODE(strap_sticky[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__B2 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__B (.DIODE(strap_sticky[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__C_N (.DIODE(strap_sticky[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__B2 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06668__B (.DIODE(strap_sticky[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06668__C (.DIODE(strap_sticky[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06669__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__06669__B2 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__A1 (.DIODE(strap_sticky[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__A2 (.DIODE(strap_sticky[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__B2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__A (.DIODE(strap_sticky[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06673__B (.DIODE(strap_sticky[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__B2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06676__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__06676__B2 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__A (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__B (.DIODE(strap_sticky[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__C (.DIODE(strap_sticky[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__B2 (.DIODE(_02733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__B1 (.DIODE(wbs_ack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__C_N (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__A1 (.DIODE(wbs_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__A1 (.DIODE(wbs_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06693__A1 (.DIODE(wbs_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__A1 (.DIODE(wbs_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__A1 (.DIODE(wbs_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06701__A1 (.DIODE(wbs_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06703__A1 (.DIODE(wbs_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__A1 (.DIODE(wbs_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06708__A1 (.DIODE(wbs_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__A1 (.DIODE(wbs_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06712__A1 (.DIODE(wbs_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06716__A1 (.DIODE(wbs_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__A1 (.DIODE(wbs_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__A1 (.DIODE(wbs_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__A1 (.DIODE(wbs_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06725__A1 (.DIODE(wbs_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06727__A1 (.DIODE(wbs_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06729__A1 (.DIODE(wbs_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06731__A1 (.DIODE(wbs_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06734__A1 (.DIODE(wbs_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__A1 (.DIODE(wbs_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06738__A1 (.DIODE(wbs_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__A1 (.DIODE(wbs_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06743__A1 (.DIODE(wbs_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__A1 (.DIODE(wbs_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06747__A1 (.DIODE(wbs_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06749__A1 (.DIODE(wbs_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__A1 (.DIODE(wbs_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06754__A1 (.DIODE(wbs_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__A1 (.DIODE(wbs_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__A1 (.DIODE(wbs_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__A1 (.DIODE(wbs_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__A1 (.DIODE(wbs_err_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06765__A (.DIODE(wbs_ack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__06768__A (.DIODE(_01530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06769__A (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__A (.DIODE(wbs_ack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__A1 (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__A (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__A (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__A (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A (.DIODE(\u_async_wb.u_cmd_if.grey_wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__A (.DIODE(_02807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06795__A (.DIODE(\u_async_wb.u_cmd_if.grey_wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__A0 (.DIODE(wbs_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06801__A0 (.DIODE(wbs_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06803__A0 (.DIODE(wbs_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__A0 (.DIODE(wbs_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06808__A0 (.DIODE(wbs_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06810__A0 (.DIODE(wbs_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__A0 (.DIODE(wbs_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__A0 (.DIODE(wbs_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__A0 (.DIODE(wbs_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__A0 (.DIODE(wbs_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06821__A0 (.DIODE(wbs_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06823__A0 (.DIODE(wbs_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__A0 (.DIODE(wbs_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__A0 (.DIODE(wbs_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06831__A0 (.DIODE(wbs_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__A0 (.DIODE(wbs_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06836__A0 (.DIODE(wbs_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06838__A0 (.DIODE(wbs_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06840__A0 (.DIODE(wbs_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__A0 (.DIODE(wbs_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06845__A0 (.DIODE(wbs_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__A0 (.DIODE(wbs_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__A0 (.DIODE(wbs_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__A0 (.DIODE(wbs_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06854__A0 (.DIODE(wbs_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06856__A0 (.DIODE(wbs_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__A0 (.DIODE(wbs_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__A0 (.DIODE(wbs_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A0 (.DIODE(wbs_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__A0 (.DIODE(wbs_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__A0 (.DIODE(wbs_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06869__A0 (.DIODE(wbs_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__A0 (.DIODE(wbs_err_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__B (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__A (.DIODE(wbm_cyc_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__A1 (.DIODE(wbm_cyc_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__A2 (.DIODE(wbm_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__A2 (.DIODE(_01731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__B2 (.DIODE(_01731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__B (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__A3 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__A (.DIODE(_02930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__B1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__B (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__B1 (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__D1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__B1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__A (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A2 (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__C1 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07009__B1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__A (.DIODE(_02930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__A (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__B (.DIODE(_02996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__B1 (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__A2 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__A2 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__A2 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__B1 (.DIODE(_02996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__A2 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__B (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A2 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A2 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__B1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__A2 (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__B2 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__B (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A2 (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__A2 (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__C (.DIODE(_03079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__B1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__B1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A (.DIODE(_03091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__B1 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__B2 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A2 (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__C (.DIODE(_03079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__A2 (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__A (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__B1 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A2 (.DIODE(_03132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A2 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A2 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__A (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A2 (.DIODE(_03139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__C (.DIODE(_03079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__B1 (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A2 (.DIODE(_02953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A2 (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B2 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A2 (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__C (.DIODE(_03079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__B1 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A (.DIODE(_03091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__A2 (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__B2 (.DIODE(wbm_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A (.DIODE(_03178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__A (.DIODE(_02415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A2 (.DIODE(\u_spi2wb.reg_be[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__B1 (.DIODE(wbm_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A0 (.DIODE(_03185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__A0 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__A0 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A0 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__A (.DIODE(_02807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A (.DIODE(_03191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A (.DIODE(_03192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A0 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A0 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A0 (.DIODE(_02473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07298__A (.DIODE(_03192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A0 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A0 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__A0 (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__A (.DIODE(_03192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__A0 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__A (.DIODE(_03192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A0 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__A0 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A0 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__A (.DIODE(_02807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A0 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A0 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A0 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A0 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A0 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07338__A0 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__A0 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__A0 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A0 (.DIODE(_02733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A0 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07349__A (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A0 (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__A0 (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__A0 (.DIODE(_02531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__A (.DIODE(_01485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A1 (.DIODE(wbm_adr_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__A0 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A1 (.DIODE(wbm_adr_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A0 (.DIODE(_03241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A (.DIODE(_02807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A (.DIODE(_01775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__A1 (.DIODE(wbm_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__A0 (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__A1 (.DIODE(wbm_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A0 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__A1 (.DIODE(wbm_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__A0 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07399__A (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A1 (.DIODE(_01731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__B1 (.DIODE(wbm_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__A0 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A1 (.DIODE(wbm_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__A0 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__A (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__B1 (.DIODE(wbm_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A0 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__B1 (.DIODE(wbm_adr_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__A0 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__B1 (.DIODE(wbm_adr_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__A0 (.DIODE(_03283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07424__A (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__B1 (.DIODE(wbm_adr_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__A0 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A1 (.DIODE(wbm_adr_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A0 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__B1 (.DIODE(wbm_adr_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07436__A0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__B1 (.DIODE(wbm_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A0 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__A1 (.DIODE(wbm_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__B1 (.DIODE(wbm_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__A (.DIODE(_03191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__A0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A (.DIODE(_03191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A (.DIODE(_03191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__A1 (.DIODE(_03185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__A1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A (.DIODE(_03338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__A (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__A (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A (.DIODE(_03338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A1 (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A1 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__A1 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A1 (.DIODE(_02733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__A (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A1 (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__A1 (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__A (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A1 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07570__A1 (.DIODE(_03241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__A (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A1 (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A1 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07585__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__A1 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A1 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__A1 (.DIODE(_03283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__A1 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A1 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A1 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A1 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__A1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A (.DIODE(_03338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A (.DIODE(_03338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__S (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__S (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__S (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__A (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__A0 (.DIODE(_03185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__A0 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__A0 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__A0 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__A0 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__A0 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A0 (.DIODE(_02473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__A (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07666__A (.DIODE(_03427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__A0 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__A0 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__A0 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A0 (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__A (.DIODE(_03427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A0 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A (.DIODE(_03427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A (.DIODE(_03427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__A0 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A (.DIODE(_03448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__A0 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__A0 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A0 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A0 (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A (.DIODE(_03448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__A0 (.DIODE(_02733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__A0 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__A0 (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__A0 (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07721__A (.DIODE(_03448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__A0 (.DIODE(_02531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A0 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A0 (.DIODE(_03241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__A (.DIODE(_03448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A0 (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__A0 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07743__A0 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A0 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__A0 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__A0 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A0 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07754__A0 (.DIODE(_03283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__A0 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A0 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A0 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A (.DIODE(_03502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__A1 (.DIODE(_03185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A1 (.DIODE(_02238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A (.DIODE(_03502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__A (.DIODE(_03520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__A (.DIODE(_03520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07847__A (.DIODE(_03520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A (.DIODE(_03520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__A (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07867__A1 (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__A1 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__A1 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A1 (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A1 (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A1 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A1 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A1 (.DIODE(_03241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A1 (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__A1 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A (.DIODE(_03502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A1 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__A1 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A1 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A1 (.DIODE(_03279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A1 (.DIODE(_03283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A1 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A1 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A1 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A1 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__A (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A (.DIODE(_03519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__A1 (.DIODE(\u_async_wb.m_cmd_wr_data[65] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__B2 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__A2 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__B1 (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__B2 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__B2 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A2 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__B1 (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__B2 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__A2 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__B1 (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__B2 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__B2 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__B (.DIODE(_01739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__A1 (.DIODE(\wb_dat_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__A1 (.DIODE(\wb_dat_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__A1 (.DIODE(\wb_dat_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A1 (.DIODE(\wb_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A1 (.DIODE(\wb_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__A1 (.DIODE(\wb_dat_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A1 (.DIODE(\wb_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__A (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__A1 (.DIODE(\wb_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__A1 (.DIODE(\wb_dat_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__A1 (.DIODE(\wb_dat_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A1 (.DIODE(\wb_dat_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__A1 (.DIODE(\wb_dat_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__A1 (.DIODE(\wb_dat_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__A1 (.DIODE(\wb_dat_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08031__A1 (.DIODE(\wb_dat_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__A (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A1 (.DIODE(\wb_dat_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__A1 (.DIODE(\wb_dat_o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__A1 (.DIODE(\wb_dat_o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__A1 (.DIODE(\wb_dat_o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__A (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A1 (.DIODE(\wb_dat_o[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__A (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__A1 (.DIODE(\wb_dat_o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A1 (.DIODE(\wb_dat_o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__A1 (.DIODE(\wb_dat_o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A1 (.DIODE(\wb_dat_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__A1 (.DIODE(\wb_dat_o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__A1 (.DIODE(\wb_dat_o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__A1 (.DIODE(\wb_dat_o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A1 (.DIODE(\wb_dat_o[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__A (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__A1 (.DIODE(\wb_dat_o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A1 (.DIODE(\wb_dat_o[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A1 (.DIODE(\wb_dat_o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A1 (.DIODE(\wb_dat_o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__B1 (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A1 (.DIODE(_01511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A (.DIODE(_01511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A (.DIODE(\u_uart2wb.auto_rx_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__S (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__S (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__S (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__S (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__A1 (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__S (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A1 (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__S (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__A1 (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__S (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__A1 (.DIODE(_03711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__S (.DIODE(_03712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__S (.DIODE(_03712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__A1 (.DIODE(_03716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__S (.DIODE(_03712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08161__S (.DIODE(_03712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__A (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__A (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__A (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__A1 (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__B1 (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__A1 (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__B1 (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__A (.DIODE(_03711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A1 (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__B1 (.DIODE(_03711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__A (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__B1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__B1 (.DIODE(_03716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A1 (.DIODE(_03716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__A1 (.DIODE(\u_uart2wb.auto_baud_16x[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A1 (.DIODE(\u_uart2wb.auto_baud_16x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__D1 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__A (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__A (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A (.DIODE(_03804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__A (.DIODE(_03876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B (.DIODE(la_data_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__C_N (.DIODE(la_data_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__A1 (.DIODE(\u_uart2wb.tx_data_avail ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__A (.DIODE(\u_uart2wb.u_core.si_ss ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08427__A_N (.DIODE(_01163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A (.DIODE(_01149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A (.DIODE(la_data_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__A (.DIODE(\u_uart2wb.auto_rx_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__C1 (.DIODE(\u_uart2wb.u_core.si_ss ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__A1 (.DIODE(\u_uart2wb.u_core.si_ss ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__A1 (.DIODE(\u_uart2wb.u_core.si_ss ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08458__B (.DIODE(_01149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__B (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__A1 (.DIODE(la_data_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__B2 (.DIODE(\u_uart2wb.auto_baud_16x[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__A (.DIODE(strap_uartm[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08546__A (.DIODE(la_data_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__A (.DIODE(strap_uartm[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__A (.DIODE(la_data_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__A (.DIODE(la_data_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__B_N (.DIODE(strap_uartm[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A1 (.DIODE(la_data_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__B (.DIODE(la_data_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A1 (.DIODE(la_data_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A2 (.DIODE(la_data_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__A1 (.DIODE(la_data_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__A1 (.DIODE(la_data_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__B1 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__A1 (.DIODE(la_data_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__B1 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__A1 (.DIODE(la_data_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__B1 (.DIODE(_01436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__B2 (.DIODE(\u_uart2wb.auto_baud_16x[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__08696__A (.DIODE(_04170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__A (.DIODE(_04170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08714__A (.DIODE(_04170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__A1 (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__A1 (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__A1 (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__A1 (.DIODE(_03711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A (.DIODE(_04170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08724__A1 (.DIODE(_03714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__A1 (.DIODE(_03716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__A1 (.DIODE(_02930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__A2 (.DIODE(_02940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08768__A (.DIODE(_03132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__A2 (.DIODE(_03139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__A2 (.DIODE(_03139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__B1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__B2 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A2 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__B1 (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__B2 (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__B2 (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__B2 (.DIODE(_02531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__A (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__B (.DIODE(_03178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08830__A0 (.DIODE(\u_reg.cfg_glb_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__A1 (.DIODE(_02238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08900__A1 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__A (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__B (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__B1 (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__B2 (.DIODE(_04339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__B2 (.DIODE(_04340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08940__B1 (.DIODE(_04341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__A (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08968__A (.DIODE(_04352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08970__A (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__B (.DIODE(_04352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__A (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__B2 (.DIODE(_04333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__B2 (.DIODE(_04339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__B2 (.DIODE(_04340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__B2 (.DIODE(_04341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A (.DIODE(_04352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__A (.DIODE(_04356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__B1 (.DIODE(\u_uart2wb.tx_data_avail ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09044__A (.DIODE(_03091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A2 (.DIODE(_03132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__A2 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09053__A2 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__B1 (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__C (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__B1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A2 (.DIODE(_03065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A2_N (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__A (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__A1 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A2 (.DIODE(_03132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__B1_N (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09128__C (.DIODE(_04453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A2 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__C1 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__A2 (.DIODE(_03139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__B1 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__A2 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__A (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__A1 (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__B (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__A (.DIODE(_03091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__B1 (.DIODE(_02952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__C1 (.DIODE(_02996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A2 (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__B2 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__C (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__B1 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__B1 (.DIODE(_03145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__B1 (.DIODE(_02930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__B (.DIODE(_02996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__A_N (.DIODE(\u_spi2wb.u_if.sck_l1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__A1 (.DIODE(\wb_dat_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__A1 (.DIODE(\wb_dat_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A1 (.DIODE(\wb_dat_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__A (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A1 (.DIODE(\wb_dat_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09260__A1 (.DIODE(\wb_dat_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A1 (.DIODE(\wb_dat_o[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__A1 (.DIODE(\wb_dat_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__A (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A1 (.DIODE(\wb_dat_o[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09274__A1 (.DIODE(\wb_dat_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__A1 (.DIODE(\wb_dat_o[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__A1 (.DIODE(\wb_dat_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A1 (.DIODE(\wb_dat_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A1 (.DIODE(\wb_dat_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__A1 (.DIODE(\wb_dat_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A1 (.DIODE(\wb_dat_o[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__A (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A1 (.DIODE(\wb_dat_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__A1 (.DIODE(\wb_dat_o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A1 (.DIODE(\wb_dat_o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A1 (.DIODE(\wb_dat_o[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A1 (.DIODE(\wb_dat_o[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__A1 (.DIODE(\wb_dat_o[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__A1 (.DIODE(\wb_dat_o[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A1 (.DIODE(\wb_dat_o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A1 (.DIODE(\wb_dat_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__A1 (.DIODE(\wb_dat_o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__A1 (.DIODE(\wb_dat_o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A1 (.DIODE(\wb_dat_o[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__A1 (.DIODE(\wb_dat_o[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__A1 (.DIODE(\wb_dat_o[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__A1 (.DIODE(\wb_dat_o[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__A1 (.DIODE(\wb_dat_o[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A1 (.DIODE(\wb_dat_o[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__S (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__A1 (.DIODE(\u_spi2wb.u_if.ssn_l1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A (.DIODE(_01835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__B1 (.DIODE(\u_spi2wb.reg_wr ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__RESET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__09367__RESET_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__RESET_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__RESET_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__RESET_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__RESET_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__RESET_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__RESET_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__RESET_B (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09391__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09394__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__D (.DIODE(sclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__SET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__D (.DIODE(ssn));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__RESET_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__RESET_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__RESET_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__RESET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__RESET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__RESET_B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__RESET_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09462__RESET_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__RESET_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__RESET_B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09465__RESET_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__RESET_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__RESET_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__RESET_B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__RESET_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__RESET_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__RESET_B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__RESET_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__RESET_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__D (.DIODE(strap_sticky[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__RESET_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__RESET_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__RESET_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__RESET_B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__RESET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__RESET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__RESET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__RESET_B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__RESET_B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__RESET_B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__RESET_B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__RESET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__RESET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__RESET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__SET_B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__RESET_B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__RESET_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__RESET_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__RESET_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__RESET_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__RESET_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__RESET_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__RESET_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__RESET_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__RESET_B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09624__RESET_B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09682__RESET_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__RESET_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__RESET_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__D (.DIODE(\u_async_wb.u_cmd_if.grey_wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09694__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09696__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__RESET_B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09740__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09742__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__RESET_B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__D (.DIODE(wbs_ack_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__RESET_B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__RESET_B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__D (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__SET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__RESET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__RESET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__RESET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__RESET_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__RESET_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__RESET_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__D (.DIODE(wb_ack_o1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__RESET_B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__D (.DIODE(wb_err_o1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__RESET_B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__RESET_B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__RESET_B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__RESET_B (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__RESET_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__RESET_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__RESET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__10119__RESET_B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__RESET_B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__RESET_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__RESET_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__RESET_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__RESET_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__RESET_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__RESET_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__RESET_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__RESET_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__RESET_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__RESET_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__RESET_B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__RESET_B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__RESET_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10169__RESET_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10170__RESET_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__RESET_B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__RESET_B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__RESET_B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__RESET_B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__RESET_B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__RESET_B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__RESET_B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__RESET_B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__RESET_B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__10193__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__D (.DIODE(uartm_rxd));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__SET_B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__RESET_B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__RESET_B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__RESET_B (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__RESET_B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__RESET_B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__RESET_B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__RESET_B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__RESET_B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__RESET_B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__RESET_B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__RESET_B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__RESET_B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__RESET_B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__RESET_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__RESET_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__RESET_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__RESET_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__RESET_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10257__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10266__RESET_B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__RESET_B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__RESET_B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__RESET_B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__RESET_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__RESET_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__D (.DIODE(uartm_rxd));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__SET_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__RESET_B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__CLK (.DIODE(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__RESET_B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__RESET_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__RESET_B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__RESET_B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__RESET_B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__RESET_B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__RESET_B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__RESET_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__RESET_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__RESET_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__RESET_B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10392__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10395__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10399__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__RESET_B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__RESET_B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__RESET_B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__RESET_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__RESET_B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__RESET_B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__RESET_B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__CLK (.DIODE(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__RESET_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__RESET_B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__RESET_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__RESET_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__RESET_B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__RESET_B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__RESET_B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__SET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__RESET_B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_0_u_async_wb.u_cmd_if.rd_clk_A  (.DIODE(\u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_0_u_uart2wb.baud_clk_16x_A  (.DIODE(\u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_wbm_clk_i_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_1_0__f_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_0_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_1_1__f_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_0_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_0__f_u_async_wb.u_cmd_if.rd_clk_A  (.DIODE(\clknet_0_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_wbm_clk_i_A (.DIODE(clknet_0_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_1__f_u_async_wb.u_cmd_if.rd_clk_A  (.DIODE(\clknet_0_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_wbm_clk_i_A (.DIODE(clknet_0_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_2__f_u_async_wb.u_cmd_if.rd_clk_A  (.DIODE(\clknet_0_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_wbm_clk_i_A (.DIODE(clknet_0_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_3__f_u_async_wb.u_cmd_if.rd_clk_A  (.DIODE(\clknet_0_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_wbm_clk_i_A (.DIODE(clknet_0_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_4__f_u_async_wb.u_cmd_if.rd_clk_A  (.DIODE(\clknet_0_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_wbm_clk_i_A (.DIODE(clknet_0_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_5__f_u_async_wb.u_cmd_if.rd_clk_A  (.DIODE(\clknet_0_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_wbm_clk_i_A (.DIODE(clknet_0_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_6__f_u_async_wb.u_cmd_if.rd_clk_A  (.DIODE(\clknet_0_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_wbm_clk_i_A (.DIODE(clknet_0_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_3_7__f_u_async_wb.u_cmd_if.rd_clk_A  (.DIODE(\clknet_0_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_wbm_clk_i_A (.DIODE(clknet_0_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_0_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_10_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_11_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_12_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_13_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_14_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_15_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_16_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_17_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_18_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_19_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_1_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_20_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_21_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_22_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_23_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_24_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_25_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_26_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_27_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_2_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wbm_clk_i_A (.DIODE(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_3_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_wbm_clk_i_A (.DIODE(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_4_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_wbm_clk_i_A (.DIODE(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_wbm_clk_i_A (.DIODE(clknet_3_7__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_wbm_clk_i_A (.DIODE(clknet_3_7__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_wbm_clk_i_A (.DIODE(clknet_3_7__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_wbm_clk_i_A (.DIODE(clknet_3_7__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_5_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_wbm_clk_i_A (.DIODE(clknet_3_7__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_wbm_clk_i_A (.DIODE(clknet_3_7__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_wbm_clk_i_A (.DIODE(clknet_3_7__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_wbm_clk_i_A (.DIODE(clknet_3_7__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_6_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_wbm_clk_i_A (.DIODE(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_7_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_wbm_clk_i_A (.DIODE(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_8_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_wbm_clk_i_A (.DIODE(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_leaf_9_u_uart2wb.baud_clk_16x_A  (.DIODE(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wbm_clk_i_A (.DIODE(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold15_A (.DIODE(wbm_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold21_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(\u_spi2wb.u_if.sck_l1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold47_A (.DIODE(wbm_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold48_A (.DIODE(\u_spi2wb.u_if.ssn_l1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output10_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_output11_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_output12_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_output13_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_output14_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_output153_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_output154_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_output17_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_output188_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_output18_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_output190_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output196_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_output197_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_output198_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_output199_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_output19_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_output200_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_output201_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_output202_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_output204_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_output209_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_output20_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_output210_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_output211_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_output212_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_output213_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_output214_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_output24_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output8_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_output9_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_clkgate.u_gate_CLK  (.DIODE(wbs_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_reg.u_fastsim_buf.u_buf_A  (.DIODE(\u_reg.cfg_glb_ctrl[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_clkbuf_in.u_buf_A  (.DIODE(wbd_clk_int));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_00.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_01.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_02.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_03.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_04.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_05.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_06.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_07.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_10.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_11.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_12.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_13.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_20.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[2]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_21.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[2]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_wh.u_mux_level_30.genblk1.u_mux_S  (.DIODE(cfg_cska_wh[3]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_uart2wb.u_arst_sync.u_buf.genblk1.u_mux_A1  (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_uart2wb.u_core.u_line_rst.u_buf.genblk1.u_mux_A1  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1_A (.DIODE(wbm_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire306_A (.DIODE(user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire307_A (.DIODE(user_clock1));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire308_A (.DIODE(sdin));
 sky130_fd_sc_hd__decap_4 FILLER_0_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 _04631_ (.A(\u_uart2wb.u_core.u_txfsm.divcnt[0] ),
    .X(_01105_));
 sky130_fd_sc_hd__clkinv_2 _04632_ (.A(_01105_),
    .Y(_00032_));
 sky130_fd_sc_hd__inv_2 _04633_ (.A(net286),
    .Y(_01106_));
 sky130_fd_sc_hd__clkbuf_2 _04634_ (.A(_01106_),
    .X(_01107_));
 sky130_fd_sc_hd__buf_2 _04635_ (.A(_01107_),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04636_ (.A(\u_uart2wb.u_core.u_rxfsm.offset[0] ),
    .X(_01108_));
 sky130_fd_sc_hd__clkinv_2 _04637_ (.A(_01108_),
    .Y(_00028_));
 sky130_fd_sc_hd__inv_2 _04638_ (.A(\u_spi2wb.u_if.ssn_l1 ),
    .Y(_01109_));
 sky130_fd_sc_hd__clkbuf_1 _04639_ (.A(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__clkbuf_1 _04640_ (.A(\u_spi2wb.u_if.spi_if_st[0] ),
    .X(_01111_));
 sky130_fd_sc_hd__clkbuf_1 _04641_ (.A(\u_spi2wb.u_if.spi_if_st[1] ),
    .X(_01112_));
 sky130_fd_sc_hd__or2b_2 _04642_ (.A(\u_spi2wb.u_if.sck_l2 ),
    .B_N(\u_spi2wb.u_if.sck_l1 ),
    .X(_01113_));
 sky130_fd_sc_hd__and3_1 _04643_ (.A(\u_spi2wb.u_if.bitcnt[1] ),
    .B(\u_spi2wb.u_if.bitcnt[0] ),
    .C(\u_spi2wb.u_if.bitcnt[2] ),
    .X(_01114_));
 sky130_fd_sc_hd__inv_2 _04644_ (.A(_01114_),
    .Y(_01115_));
 sky130_fd_sc_hd__or4_1 _04645_ (.A(\u_spi2wb.u_if.bitcnt[3] ),
    .B(\u_spi2wb.u_if.bitcnt[5] ),
    .C(\u_spi2wb.u_if.bitcnt[4] ),
    .D(_01115_),
    .X(_01116_));
 sky130_fd_sc_hd__or2_1 _04646_ (.A(_01113_),
    .B(_01116_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _04647_ (.A0(_01112_),
    .A1(\u_spi2wb.u_if.cmd_phase ),
    .S(_01117_),
    .X(_01118_));
 sky130_fd_sc_hd__or2_1 _04648_ (.A(_01111_),
    .B(_01118_),
    .X(_01119_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04649_ (.A(\u_spi2wb.u_if.rd_phase ),
    .X(_01120_));
 sky130_fd_sc_hd__nor4b_1 _04650_ (.A(\u_spi2wb.u_if.cmd_reg[5] ),
    .B(\u_spi2wb.u_if.cmd_reg[7] ),
    .C(\u_spi2wb.u_if.cmd_reg[6] ),
    .D_N(\u_spi2wb.u_if.cmd_reg[4] ),
    .Y(_01121_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04651_ (.A(\u_spi2wb.u_if.adr_phase ),
    .X(_01122_));
 sky130_fd_sc_hd__or4b_1 _04652_ (.A(\u_spi2wb.u_if.cmd_reg[4] ),
    .B(\u_spi2wb.u_if.cmd_reg[7] ),
    .C(\u_spi2wb.u_if.cmd_reg[6] ),
    .D_N(\u_spi2wb.u_if.cmd_reg[5] ),
    .X(_01123_));
 sky130_fd_sc_hd__and3b_1 _04653_ (.A_N(_01121_),
    .B(_01122_),
    .C(_01123_),
    .X(_01124_));
 sky130_fd_sc_hd__and2_1 _04654_ (.A(\u_spi2wb.u_if.bitcnt[3] ),
    .B(_01114_),
    .X(_01125_));
 sky130_fd_sc_hd__nand2_1 _04655_ (.A(\u_spi2wb.u_if.bitcnt[4] ),
    .B(_01125_),
    .Y(_01126_));
 sky130_fd_sc_hd__clkbuf_1 _04656_ (.A(_01126_),
    .X(_01127_));
 sky130_fd_sc_hd__clkbuf_1 _04657_ (.A(\u_spi2wb.u_if.bitcnt[5] ),
    .X(_01128_));
 sky130_fd_sc_hd__and2b_1 _04658_ (.A_N(\u_spi2wb.u_if.sck_l2 ),
    .B(\u_spi2wb.u_if.sck_l1 ),
    .X(_01129_));
 sky130_fd_sc_hd__clkbuf_1 _04659_ (.A(_01129_),
    .X(_01130_));
 sky130_fd_sc_hd__and4bb_1 _04660_ (.A_N(_01127_),
    .B_N(_01128_),
    .C(_01110_),
    .D(_01130_),
    .X(_01131_));
 sky130_fd_sc_hd__clkbuf_1 _04661_ (.A(_01131_),
    .X(_01132_));
 sky130_fd_sc_hd__o21a_1 _04662_ (.A1(_01120_),
    .A2(_01124_),
    .B1(_01132_),
    .X(_01133_));
 sky130_fd_sc_hd__a21o_1 _04663_ (.A1(_01110_),
    .A2(_01119_),
    .B1(_01133_),
    .X(_00005_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04664_ (.A(\u_uart2wb.u_core.u_txfsm.divcnt[1] ),
    .X(_01134_));
 sky130_fd_sc_hd__nor4_2 _04665_ (.A(\u_uart2wb.u_core.u_txfsm.divcnt[0] ),
    .B(_01134_),
    .C(\u_uart2wb.u_core.u_txfsm.divcnt[3] ),
    .D(\u_uart2wb.u_core.u_txfsm.divcnt[2] ),
    .Y(_01135_));
 sky130_fd_sc_hd__clkbuf_1 _04666_ (.A(\u_uart2wb.u_core.u_txfsm.cnt[2] ),
    .X(_01136_));
 sky130_fd_sc_hd__clkbuf_1 _04667_ (.A(\u_uart2wb.u_core.u_txfsm.txstate[3] ),
    .X(_01137_));
 sky130_fd_sc_hd__or4_2 _04668_ (.A(\u_uart2wb.u_core.u_txfsm.divcnt[0] ),
    .B(\u_uart2wb.u_core.u_txfsm.divcnt[1] ),
    .C(\u_uart2wb.u_core.u_txfsm.divcnt[3] ),
    .D(\u_uart2wb.u_core.u_txfsm.divcnt[2] ),
    .X(_01138_));
 sky130_fd_sc_hd__clkbuf_1 _04669_ (.A(\u_uart2wb.u_core.u_txfsm.cnt[1] ),
    .X(_01139_));
 sky130_fd_sc_hd__clkbuf_1 _04670_ (.A(\u_uart2wb.u_core.u_txfsm.cnt[0] ),
    .X(_01140_));
 sky130_fd_sc_hd__nand2_1 _04671_ (.A(_01139_),
    .B(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_1 _04672_ (.A(_01138_),
    .B(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__and3_1 _04673_ (.A(_01136_),
    .B(_01137_),
    .C(_01142_),
    .X(_01143_));
 sky130_fd_sc_hd__clkbuf_1 _04674_ (.A(strap_uartm[1]),
    .X(_01144_));
 sky130_fd_sc_hd__and2_1 _04675_ (.A(strap_uartm[0]),
    .B(_01144_),
    .X(_01145_));
 sky130_fd_sc_hd__clkbuf_1 _04676_ (.A(_01145_),
    .X(_01146_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04677_ (.A(_01146_),
    .X(_01147_));
 sky130_fd_sc_hd__or2_1 _04678_ (.A(la_data_in[16]),
    .B(la_data_in[17]),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_1 _04679_ (.A(_01147_),
    .B(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__and2_1 _04680_ (.A(\u_uart2wb.u_core.u_txfsm.txstate[4] ),
    .B(_01138_),
    .X(_01150_));
 sky130_fd_sc_hd__a221o_1 _04681_ (.A1(\u_uart2wb.u_core.u_txfsm.txstate[2] ),
    .A2(_01135_),
    .B1(_01143_),
    .B2(_01149_),
    .C1(_01150_),
    .X(_00019_));
 sky130_fd_sc_hd__inv_2 _04682_ (.A(_01137_),
    .Y(_01151_));
 sky130_fd_sc_hd__a21o_1 _04683_ (.A1(_01136_),
    .A2(_01142_),
    .B1(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__clkbuf_1 _04684_ (.A(strap_uartm[0]),
    .X(_01153_));
 sky130_fd_sc_hd__clkbuf_1 _04685_ (.A(_01153_),
    .X(_01154_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04686_ (.A(_01144_),
    .X(_01155_));
 sky130_fd_sc_hd__nand2_2 _04687_ (.A(_01154_),
    .B(_01155_),
    .Y(_01156_));
 sky130_fd_sc_hd__or2_2 _04688_ (.A(_01154_),
    .B(_01155_),
    .X(_01157_));
 sky130_fd_sc_hd__o22a_1 _04689_ (.A1(la_data_in[1]),
    .A2(_01156_),
    .B1(_01157_),
    .B2(\u_uart2wb.auto_rx_enb ),
    .X(_01158_));
 sky130_fd_sc_hd__clkbuf_1 _04690_ (.A(_01158_),
    .X(_01159_));
 sky130_fd_sc_hd__nand4_1 _04691_ (.A(\u_uart2wb.tx_data_avail ),
    .B(\u_uart2wb.u_core.u_txfsm.txstate[0] ),
    .C(_01135_),
    .D(_01159_),
    .Y(_01160_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04692_ (.A(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__nand2_1 _04693_ (.A(_01152_),
    .B(_01161_),
    .Y(_00018_));
 sky130_fd_sc_hd__clkbuf_1 _04694_ (.A(_01138_),
    .X(_01162_));
 sky130_fd_sc_hd__a32o_1 _04695_ (.A1(_01147_),
    .A2(_01148_),
    .A3(_01143_),
    .B1(_01162_),
    .B2(\u_uart2wb.u_core.u_txfsm.txstate[2] ),
    .X(_00017_));
 sky130_fd_sc_hd__nor2_2 _04696_ (.A(la_data_in[3]),
    .B(_01156_),
    .Y(_01163_));
 sky130_fd_sc_hd__nor2_1 _04697_ (.A(_01162_),
    .B(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__a22o_1 _04698_ (.A1(\u_uart2wb.u_core.u_txfsm.txstate[1] ),
    .A2(_01162_),
    .B1(_01164_),
    .B2(\u_uart2wb.u_core.u_txfsm.txstate[4] ),
    .X(_00016_));
 sky130_fd_sc_hd__or2b_1 _04699_ (.A(\u_uart2wb.u_aut_det.rxd_sync[2] ),
    .B_N(\u_uart2wb.u_aut_det.rxd_sync[1] ),
    .X(_01165_));
 sky130_fd_sc_hd__clkbuf_1 _04700_ (.A(_01165_),
    .X(_01166_));
 sky130_fd_sc_hd__and2_1 _04701_ (.A(\u_uart2wb.u_aut_det.clk_cnt[18] ),
    .B(\u_uart2wb.u_aut_det.clk_cnt[19] ),
    .X(_01167_));
 sky130_fd_sc_hd__and3_1 _04702_ (.A(\u_uart2wb.u_aut_det.clk_cnt[1] ),
    .B(\u_uart2wb.u_aut_det.clk_cnt[0] ),
    .C(\u_uart2wb.u_aut_det.clk_cnt[2] ),
    .X(_01168_));
 sky130_fd_sc_hd__and3_1 _04703_ (.A(\u_uart2wb.u_aut_det.clk_cnt[3] ),
    .B(\u_uart2wb.u_aut_det.clk_cnt[4] ),
    .C(_01168_),
    .X(_01169_));
 sky130_fd_sc_hd__and4_1 _04704_ (.A(\u_uart2wb.u_aut_det.clk_cnt[5] ),
    .B(\u_uart2wb.u_aut_det.clk_cnt[7] ),
    .C(\u_uart2wb.u_aut_det.clk_cnt[6] ),
    .D(_01169_),
    .X(_01170_));
 sky130_fd_sc_hd__and3_1 _04705_ (.A(\u_uart2wb.u_aut_det.clk_cnt[9] ),
    .B(\u_uart2wb.u_aut_det.clk_cnt[8] ),
    .C(_01170_),
    .X(_01171_));
 sky130_fd_sc_hd__and3_1 _04706_ (.A(\u_uart2wb.u_aut_det.clk_cnt[11] ),
    .B(\u_uart2wb.u_aut_det.clk_cnt[10] ),
    .C(\u_uart2wb.u_aut_det.clk_cnt[12] ),
    .X(_01172_));
 sky130_fd_sc_hd__and3_1 _04707_ (.A(\u_uart2wb.u_aut_det.clk_cnt[13] ),
    .B(_01171_),
    .C(_01172_),
    .X(_01173_));
 sky130_fd_sc_hd__and4_1 _04708_ (.A(\u_uart2wb.u_aut_det.clk_cnt[15] ),
    .B(\u_uart2wb.u_aut_det.clk_cnt[14] ),
    .C(\u_uart2wb.u_aut_det.clk_cnt[16] ),
    .D(_01173_),
    .X(_01174_));
 sky130_fd_sc_hd__nand3_1 _04709_ (.A(\u_uart2wb.u_aut_det.clk_cnt[17] ),
    .B(_01167_),
    .C(_01174_),
    .Y(_01175_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04710_ (.A(_01175_),
    .X(_01176_));
 sky130_fd_sc_hd__clkbuf_1 _04711_ (.A(_01176_),
    .X(_01177_));
 sky130_fd_sc_hd__and2b_1 _04712_ (.A_N(\u_uart2wb.u_aut_det.rxd_sync[1] ),
    .B(\u_uart2wb.u_aut_det.rxd_sync[2] ),
    .X(_01178_));
 sky130_fd_sc_hd__and2_1 _04713_ (.A(\u_uart2wb.u_aut_det.state[2] ),
    .B(_01178_),
    .X(_01179_));
 sky130_fd_sc_hd__clkbuf_2 _04714_ (.A(_01179_),
    .X(_01180_));
 sky130_fd_sc_hd__a31o_1 _04715_ (.A1(\u_uart2wb.u_aut_det.state[6] ),
    .A2(_01166_),
    .A3(_01177_),
    .B1(_01180_),
    .X(_00013_));
 sky130_fd_sc_hd__and2b_1 _04716_ (.A_N(\u_uart2wb.u_aut_det.rxd_sync[2] ),
    .B(\u_uart2wb.u_aut_det.rxd_sync[1] ),
    .X(_01181_));
 sky130_fd_sc_hd__and2_1 _04717_ (.A(\u_uart2wb.u_aut_det.state[3] ),
    .B(_01181_),
    .X(_01182_));
 sky130_fd_sc_hd__or2_1 _04718_ (.A(\u_uart2wb.u_aut_det.state[7] ),
    .B(_01182_),
    .X(_01183_));
 sky130_fd_sc_hd__clkbuf_1 _04719_ (.A(_01183_),
    .X(_00014_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04720_ (.A(\u_uart2wb.u_core.u_txfsm.txstate[0] ),
    .X(_01184_));
 sky130_fd_sc_hd__a21boi_1 _04721_ (.A1(\u_uart2wb.tx_data_avail ),
    .A2(_01159_),
    .B1_N(\u_uart2wb.u_core.u_txfsm.txstate[0] ),
    .Y(_01185_));
 sky130_fd_sc_hd__or2_1 _04722_ (.A(\u_uart2wb.u_core.u_txfsm.txstate[4] ),
    .B(\u_uart2wb.u_core.u_txfsm.txstate[1] ),
    .X(_01186_));
 sky130_fd_sc_hd__o211a_1 _04723_ (.A1(\u_uart2wb.u_core.u_txfsm.txstate[1] ),
    .A2(_01163_),
    .B1(_01186_),
    .C1(_01135_),
    .X(_01187_));
 sky130_fd_sc_hd__a211o_1 _04724_ (.A1(_01184_),
    .A2(_01162_),
    .B1(_01185_),
    .C1(_01187_),
    .X(_00015_));
 sky130_fd_sc_hd__xnor2_1 _04725_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[4] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[4] ),
    .Y(_01188_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04726_ (.A(_01188_),
    .X(_01189_));
 sky130_fd_sc_hd__xor2_2 _04727_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[3] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[3] ),
    .X(_01190_));
 sky130_fd_sc_hd__xor2_1 _04728_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[2] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[2] ),
    .X(_01191_));
 sky130_fd_sc_hd__nor2_1 _04729_ (.A(_01190_),
    .B(_01191_),
    .Y(_01192_));
 sky130_fd_sc_hd__clkbuf_1 _04730_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[1] ),
    .X(_01193_));
 sky130_fd_sc_hd__clkbuf_1 _04731_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[1] ),
    .X(_01194_));
 sky130_fd_sc_hd__or2b_1 _04732_ (.A(_01193_),
    .B_N(_01194_),
    .X(_01195_));
 sky130_fd_sc_hd__or2b_1 _04733_ (.A(_01194_),
    .B_N(_01193_),
    .X(_01196_));
 sky130_fd_sc_hd__nand3b_1 _04734_ (.A_N(\u_uart2wb.u_aut_det.ref1_cnt[0] ),
    .B(_01196_),
    .C(\u_uart2wb.u_aut_det.ref2_cnt[0] ),
    .Y(_01197_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04735_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[2] ),
    .X(_01198_));
 sky130_fd_sc_hd__inv_2 _04736_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[2] ),
    .Y(_01199_));
 sky130_fd_sc_hd__clkbuf_1 _04737_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[3] ),
    .X(_01200_));
 sky130_fd_sc_hd__clkbuf_1 _04738_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[3] ),
    .X(_01201_));
 sky130_fd_sc_hd__and2b_1 _04739_ (.A_N(_01200_),
    .B(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__or2b_1 _04740_ (.A(_01201_),
    .B_N(_01200_),
    .X(_01203_));
 sky130_fd_sc_hd__o31ai_1 _04741_ (.A1(_01198_),
    .A2(_01199_),
    .A3(_01202_),
    .B1(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__a31o_1 _04742_ (.A1(_01192_),
    .A2(_01195_),
    .A3(_01197_),
    .B1(_01204_),
    .X(_01205_));
 sky130_fd_sc_hd__clkbuf_1 _04743_ (.A(_01205_),
    .X(_01206_));
 sky130_fd_sc_hd__nand3b_1 _04744_ (.A_N(\u_uart2wb.u_aut_det.ref2_cnt[0] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[0] ),
    .C(_01195_),
    .Y(_01207_));
 sky130_fd_sc_hd__a31o_1 _04745_ (.A1(_01198_),
    .A2(_01199_),
    .A3(_01203_),
    .B1(_01202_),
    .X(_01208_));
 sky130_fd_sc_hd__a31o_1 _04746_ (.A1(_01192_),
    .A2(_01196_),
    .A3(_01207_),
    .B1(_01208_),
    .X(_01209_));
 sky130_fd_sc_hd__and2b_1 _04747_ (.A_N(\u_uart2wb.u_aut_det.ref1_cnt[7] ),
    .B(\u_uart2wb.u_aut_det.ref2_cnt[7] ),
    .X(_01210_));
 sky130_fd_sc_hd__or2b_1 _04748_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[7] ),
    .B_N(\u_uart2wb.u_aut_det.ref1_cnt[7] ),
    .X(_01211_));
 sky130_fd_sc_hd__and2b_1 _04749_ (.A_N(_01210_),
    .B(_01211_),
    .X(_01212_));
 sky130_fd_sc_hd__xnor2_1 _04750_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[6] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[6] ),
    .Y(_01213_));
 sky130_fd_sc_hd__clkbuf_1 _04751_ (.A(_01213_),
    .X(_01214_));
 sky130_fd_sc_hd__xor2_1 _04752_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[5] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[5] ),
    .X(_01215_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04753_ (.A(_01215_),
    .X(_01216_));
 sky130_fd_sc_hd__and2b_1 _04754_ (.A_N(_01216_),
    .B(_01189_),
    .X(_01217_));
 sky130_fd_sc_hd__and3_1 _04755_ (.A(_01212_),
    .B(_01214_),
    .C(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__clkbuf_1 _04756_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[5] ),
    .X(_01219_));
 sky130_fd_sc_hd__clkbuf_1 _04757_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[5] ),
    .X(_01220_));
 sky130_fd_sc_hd__and2b_1 _04758_ (.A_N(_01219_),
    .B(_01220_),
    .X(_01221_));
 sky130_fd_sc_hd__clkbuf_1 _04759_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[4] ),
    .X(_01222_));
 sky130_fd_sc_hd__clkbuf_1 _04760_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[4] ),
    .X(_01223_));
 sky130_fd_sc_hd__and2b_1 _04761_ (.A_N(_01222_),
    .B(_01223_),
    .X(_01224_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04762_ (.A(_01212_),
    .X(_01225_));
 sky130_fd_sc_hd__or2b_1 _04763_ (.A(_01220_),
    .B_N(_01219_),
    .X(_01226_));
 sky130_fd_sc_hd__o2111a_1 _04764_ (.A1(_01221_),
    .A2(_01224_),
    .B1(_01225_),
    .C1(_01214_),
    .D1(_01226_),
    .X(_01227_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04765_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[6] ),
    .X(_01228_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04766_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[6] ),
    .X(_01229_));
 sky130_fd_sc_hd__inv_2 _04767_ (.A(_01229_),
    .Y(_01230_));
 sky130_fd_sc_hd__a31o_1 _04768_ (.A1(_01228_),
    .A2(_01230_),
    .A3(_01211_),
    .B1(_01210_),
    .X(_01231_));
 sky130_fd_sc_hd__a211oi_2 _04769_ (.A1(_01209_),
    .A2(_01218_),
    .B1(_01227_),
    .C1(_01231_),
    .Y(_01232_));
 sky130_fd_sc_hd__xor2_1 _04770_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[14] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[14] ),
    .X(_01233_));
 sky130_fd_sc_hd__xor2_2 _04771_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[15] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[15] ),
    .X(_01234_));
 sky130_fd_sc_hd__clkbuf_2 _04772_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[12] ),
    .X(_01235_));
 sky130_fd_sc_hd__xor2_4 _04773_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[12] ),
    .B(_01235_),
    .X(_01236_));
 sky130_fd_sc_hd__xnor2_1 _04774_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[13] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[13] ),
    .Y(_01237_));
 sky130_fd_sc_hd__inv_2 _04775_ (.A(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__or4_1 _04776_ (.A(_01233_),
    .B(_01234_),
    .C(_01236_),
    .D(_01238_),
    .X(_01239_));
 sky130_fd_sc_hd__xnor2_1 _04777_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[11] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[11] ),
    .Y(_01240_));
 sky130_fd_sc_hd__clkbuf_1 _04778_ (.A(_01240_),
    .X(_01241_));
 sky130_fd_sc_hd__xnor2_1 _04779_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[10] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[10] ),
    .Y(_01242_));
 sky130_fd_sc_hd__nand2_1 _04780_ (.A(_01241_),
    .B(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__xnor2_1 _04781_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[8] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[8] ),
    .Y(_01244_));
 sky130_fd_sc_hd__clkbuf_1 _04782_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[9] ),
    .X(_01245_));
 sky130_fd_sc_hd__clkbuf_1 _04783_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[9] ),
    .X(_01246_));
 sky130_fd_sc_hd__xnor2_1 _04784_ (.A(_01245_),
    .B(_01246_),
    .Y(_01247_));
 sky130_fd_sc_hd__nand2_1 _04785_ (.A(_01244_),
    .B(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__or2_1 _04786_ (.A(_01243_),
    .B(_01248_),
    .X(_01249_));
 sky130_fd_sc_hd__or2_1 _04787_ (.A(_01239_),
    .B(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__clkbuf_1 _04788_ (.A(_01233_),
    .X(_01251_));
 sky130_fd_sc_hd__nor2_1 _04789_ (.A(_01251_),
    .B(_01234_),
    .Y(_01252_));
 sky130_fd_sc_hd__xnor2_1 _04790_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[12] ),
    .B(_01235_),
    .Y(_01253_));
 sky130_fd_sc_hd__clkbuf_1 _04791_ (.A(_01237_),
    .X(_01254_));
 sky130_fd_sc_hd__and3_1 _04792_ (.A(_01252_),
    .B(_01253_),
    .C(_01254_),
    .X(_01255_));
 sky130_fd_sc_hd__clkbuf_1 _04793_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[11] ),
    .X(_01256_));
 sky130_fd_sc_hd__inv_2 _04794_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[11] ),
    .Y(_01257_));
 sky130_fd_sc_hd__and2_1 _04795_ (.A(_01256_),
    .B(_01257_),
    .X(_01258_));
 sky130_fd_sc_hd__and2b_1 _04796_ (.A_N(\u_uart2wb.u_aut_det.ref1_cnt[8] ),
    .B(\u_uart2wb.u_aut_det.ref2_cnt[8] ),
    .X(_01259_));
 sky130_fd_sc_hd__and2b_1 _04797_ (.A_N(\u_uart2wb.u_aut_det.ref1_cnt[9] ),
    .B(\u_uart2wb.u_aut_det.ref2_cnt[9] ),
    .X(_01260_));
 sky130_fd_sc_hd__or2b_1 _04798_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[9] ),
    .B_N(\u_uart2wb.u_aut_det.ref1_cnt[9] ),
    .X(_01261_));
 sky130_fd_sc_hd__o2111a_1 _04799_ (.A1(_01259_),
    .A2(_01260_),
    .B1(_01261_),
    .C1(_01242_),
    .D1(_01241_),
    .X(_01262_));
 sky130_fd_sc_hd__inv_2 _04800_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[10] ),
    .Y(_01263_));
 sky130_fd_sc_hd__and3_1 _04801_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[10] ),
    .B(_01263_),
    .C(_01240_),
    .X(_01264_));
 sky130_fd_sc_hd__or3_1 _04802_ (.A(_01258_),
    .B(_01262_),
    .C(_01264_),
    .X(_01265_));
 sky130_fd_sc_hd__inv_2 _04803_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[14] ),
    .Y(_01266_));
 sky130_fd_sc_hd__and2b_1 _04804_ (.A_N(\u_uart2wb.u_aut_det.ref1_cnt[15] ),
    .B(\u_uart2wb.u_aut_det.ref2_cnt[15] ),
    .X(_01267_));
 sky130_fd_sc_hd__clkbuf_1 _04805_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[15] ),
    .X(_01268_));
 sky130_fd_sc_hd__clkbuf_1 _04806_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[15] ),
    .X(_01269_));
 sky130_fd_sc_hd__and2b_1 _04807_ (.A_N(_01268_),
    .B(_01269_),
    .X(_01270_));
 sky130_fd_sc_hd__nor2_1 _04808_ (.A(_01267_),
    .B(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hd__and3_1 _04809_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[14] ),
    .B(_01266_),
    .C(_01271_),
    .X(_01272_));
 sky130_fd_sc_hd__clkbuf_1 _04810_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[13] ),
    .X(_01273_));
 sky130_fd_sc_hd__clkbuf_1 _04811_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[13] ),
    .X(_01274_));
 sky130_fd_sc_hd__and2b_1 _04812_ (.A_N(_01273_),
    .B(_01274_),
    .X(_01275_));
 sky130_fd_sc_hd__inv_2 _04813_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[12] ),
    .Y(_01276_));
 sky130_fd_sc_hd__and3_1 _04814_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[12] ),
    .B(_01276_),
    .C(_01254_),
    .X(_01277_));
 sky130_fd_sc_hd__o21a_1 _04815_ (.A1(_01275_),
    .A2(_01277_),
    .B1(_01252_),
    .X(_01278_));
 sky130_fd_sc_hd__a2111oi_1 _04816_ (.A1(_01255_),
    .A2(_01265_),
    .B1(_01272_),
    .C1(_01278_),
    .D1(_01267_),
    .Y(_01279_));
 sky130_fd_sc_hd__o21ai_1 _04817_ (.A1(_01232_),
    .A2(_01250_),
    .B1(_01279_),
    .Y(_01280_));
 sky130_fd_sc_hd__and2b_1 _04818_ (.A_N(\u_uart2wb.u_aut_det.ref1_cnt[18] ),
    .B(\u_uart2wb.u_aut_det.ref2_cnt[18] ),
    .X(_01281_));
 sky130_fd_sc_hd__clkbuf_1 _04819_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[18] ),
    .X(_01282_));
 sky130_fd_sc_hd__clkbuf_1 _04820_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[18] ),
    .X(_01283_));
 sky130_fd_sc_hd__and2b_1 _04821_ (.A_N(_01282_),
    .B(_01283_),
    .X(_01284_));
 sky130_fd_sc_hd__nor2_1 _04822_ (.A(_01281_),
    .B(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__xnor2_1 _04823_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[19] ),
    .B(\u_uart2wb.u_aut_det.ref2_cnt[19] ),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _04824_ (.A(_01285_),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__clkbuf_2 _04825_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[16] ),
    .X(_01288_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04826_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[16] ),
    .X(_01289_));
 sky130_fd_sc_hd__xnor2_2 _04827_ (.A(_01288_),
    .B(_01289_),
    .Y(_01290_));
 sky130_fd_sc_hd__xnor2_1 _04828_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[17] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[17] ),
    .Y(_01291_));
 sky130_fd_sc_hd__clkbuf_1 _04829_ (.A(_01291_),
    .X(_01292_));
 sky130_fd_sc_hd__nand2_1 _04830_ (.A(_01290_),
    .B(_01292_),
    .Y(_01293_));
 sky130_fd_sc_hd__nor2_1 _04831_ (.A(_01287_),
    .B(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__inv_2 _04832_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[19] ),
    .Y(_01295_));
 sky130_fd_sc_hd__clkbuf_1 _04833_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[17] ),
    .X(_01296_));
 sky130_fd_sc_hd__inv_2 _04834_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[17] ),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_1 _04835_ (.A(_01296_),
    .B(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__inv_2 _04836_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[16] ),
    .Y(_01299_));
 sky130_fd_sc_hd__nand3_1 _04837_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[16] ),
    .B(_01299_),
    .C(_01291_),
    .Y(_01300_));
 sky130_fd_sc_hd__a21oi_1 _04838_ (.A1(_01298_),
    .A2(_01300_),
    .B1(_01287_),
    .Y(_01301_));
 sky130_fd_sc_hd__o21a_1 _04839_ (.A1(_01295_),
    .A2(\u_uart2wb.u_aut_det.ref2_cnt[19] ),
    .B1(_01281_),
    .X(_01302_));
 sky130_fd_sc_hd__a211o_1 _04840_ (.A1(_01295_),
    .A2(\u_uart2wb.u_aut_det.ref2_cnt[19] ),
    .B1(_01301_),
    .C1(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__a21o_1 _04841_ (.A1(_01280_),
    .A2(_01294_),
    .B1(_01303_),
    .X(_01304_));
 sky130_fd_sc_hd__clkbuf_1 _04842_ (.A(_01304_),
    .X(_01305_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04843_ (.A(_01305_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _04844_ (.A0(_01206_),
    .A1(_01209_),
    .S(_01306_),
    .X(_01307_));
 sky130_fd_sc_hd__xor2_1 _04845_ (.A(_01189_),
    .B(_01307_),
    .X(_01308_));
 sky130_fd_sc_hd__a21bo_1 _04846_ (.A1(_01217_),
    .A2(_01206_),
    .B1_N(_01305_),
    .X(_01309_));
 sky130_fd_sc_hd__or2b_1 _04847_ (.A(_01223_),
    .B_N(_01222_),
    .X(_01310_));
 sky130_fd_sc_hd__a21oi_1 _04848_ (.A1(_01226_),
    .A2(_01310_),
    .B1(_01221_),
    .Y(_01311_));
 sky130_fd_sc_hd__a21oi_1 _04849_ (.A1(_01217_),
    .A2(_01206_),
    .B1(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__clkbuf_1 _04850_ (.A(_01214_),
    .X(_01313_));
 sky130_fd_sc_hd__and2b_1 _04851_ (.A_N(_01312_),
    .B(_01313_),
    .X(_01314_));
 sky130_fd_sc_hd__and2b_1 _04852_ (.A_N(_01313_),
    .B(_01312_),
    .X(_01315_));
 sky130_fd_sc_hd__or2_1 _04853_ (.A(_01314_),
    .B(_01315_),
    .X(_01316_));
 sky130_fd_sc_hd__inv_2 _04854_ (.A(_01228_),
    .Y(_01317_));
 sky130_fd_sc_hd__a21oi_1 _04855_ (.A1(_01317_),
    .A2(_01229_),
    .B1(_01314_),
    .Y(_01318_));
 sky130_fd_sc_hd__xnor2_1 _04856_ (.A(_01225_),
    .B(_01318_),
    .Y(_01319_));
 sky130_fd_sc_hd__a21oi_1 _04857_ (.A1(_01309_),
    .A2(_01316_),
    .B1(_01319_),
    .Y(_01320_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04858_ (.A(_01253_),
    .X(_01321_));
 sky130_fd_sc_hd__clkbuf_1 _04859_ (.A(_01260_),
    .X(_01322_));
 sky130_fd_sc_hd__and2b_1 _04860_ (.A_N(_01245_),
    .B(_01246_),
    .X(_01323_));
 sky130_fd_sc_hd__or2_1 _04861_ (.A(_01322_),
    .B(_01323_),
    .X(_01324_));
 sky130_fd_sc_hd__clkbuf_1 _04862_ (.A(_01324_),
    .X(_01325_));
 sky130_fd_sc_hd__and3_1 _04863_ (.A(_01225_),
    .B(_01214_),
    .C(_01311_),
    .X(_01326_));
 sky130_fd_sc_hd__a21oi_1 _04864_ (.A1(_01218_),
    .A2(_01205_),
    .B1(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__o31a_1 _04865_ (.A1(_01228_),
    .A2(_01230_),
    .A3(_01210_),
    .B1(_01211_),
    .X(_01328_));
 sky130_fd_sc_hd__a21bo_1 _04866_ (.A1(_01327_),
    .A2(_01328_),
    .B1_N(_01244_),
    .X(_01329_));
 sky130_fd_sc_hd__clkbuf_1 _04867_ (.A(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__clkbuf_1 _04868_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[8] ),
    .X(_01331_));
 sky130_fd_sc_hd__clkbuf_1 _04869_ (.A(\u_uart2wb.u_aut_det.ref1_cnt[8] ),
    .X(_01332_));
 sky130_fd_sc_hd__or2b_1 _04870_ (.A(_01331_),
    .B_N(_01332_),
    .X(_01333_));
 sky130_fd_sc_hd__a21o_1 _04871_ (.A1(_01333_),
    .A2(_01261_),
    .B1(_01322_),
    .X(_01334_));
 sky130_fd_sc_hd__clkbuf_1 _04872_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[10] ),
    .X(_01335_));
 sky130_fd_sc_hd__or3_1 _04873_ (.A(_01335_),
    .B(_01263_),
    .C(_01258_),
    .X(_01336_));
 sky130_fd_sc_hd__o221a_1 _04874_ (.A1(_01256_),
    .A2(_01257_),
    .B1(_01243_),
    .B2(_01334_),
    .C1(_01336_),
    .X(_01337_));
 sky130_fd_sc_hd__o31a_1 _04875_ (.A1(_01243_),
    .A2(_01325_),
    .A3(_01330_),
    .B1(_01337_),
    .X(_01338_));
 sky130_fd_sc_hd__xnor2_1 _04876_ (.A(_01321_),
    .B(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04877_ (.A(_01289_),
    .X(_01340_));
 sky130_fd_sc_hd__xor2_1 _04878_ (.A(_01288_),
    .B(_01340_),
    .X(_01341_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04879_ (.A(_01341_),
    .X(_01342_));
 sky130_fd_sc_hd__clkbuf_1 _04880_ (.A(_01288_),
    .X(_01343_));
 sky130_fd_sc_hd__a21o_1 _04881_ (.A1(_01343_),
    .A2(_01299_),
    .B1(_01292_),
    .X(_01344_));
 sky130_fd_sc_hd__and2_1 _04882_ (.A(_01300_),
    .B(_01344_),
    .X(_01345_));
 sky130_fd_sc_hd__clkbuf_1 _04883_ (.A(_01244_),
    .X(_01346_));
 sky130_fd_sc_hd__clkbuf_1 _04884_ (.A(_01346_),
    .X(_01347_));
 sky130_fd_sc_hd__clkbuf_1 _04885_ (.A(_01232_),
    .X(_01348_));
 sky130_fd_sc_hd__nor2_1 _04886_ (.A(_01347_),
    .B(_01348_),
    .Y(_01349_));
 sky130_fd_sc_hd__and2_1 _04887_ (.A(_01347_),
    .B(_01348_),
    .X(_01350_));
 sky130_fd_sc_hd__a211o_1 _04888_ (.A1(_01342_),
    .A2(_01345_),
    .B1(_01349_),
    .C1(_01350_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _04889_ (.A0(_01339_),
    .A1(_01351_),
    .S(_01306_),
    .X(_01352_));
 sky130_fd_sc_hd__a21o_1 _04890_ (.A1(_01327_),
    .A2(_01328_),
    .B1(_01250_),
    .X(_01353_));
 sky130_fd_sc_hd__or2b_1 _04891_ (.A(_01274_),
    .B_N(_01273_),
    .X(_01354_));
 sky130_fd_sc_hd__clkbuf_1 _04892_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[12] ),
    .X(_01355_));
 sky130_fd_sc_hd__or3_1 _04893_ (.A(_01355_),
    .B(_01276_),
    .C(_01275_),
    .X(_01356_));
 sky130_fd_sc_hd__a21bo_1 _04894_ (.A1(_01354_),
    .A2(_01356_),
    .B1_N(_01252_),
    .X(_01357_));
 sky130_fd_sc_hd__inv_2 _04895_ (.A(_01269_),
    .Y(_01358_));
 sky130_fd_sc_hd__clkbuf_1 _04896_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[14] ),
    .X(_01359_));
 sky130_fd_sc_hd__or3_1 _04897_ (.A(_01359_),
    .B(_01266_),
    .C(_01267_),
    .X(_01360_));
 sky130_fd_sc_hd__o221a_1 _04898_ (.A1(_01268_),
    .A2(_01358_),
    .B1(_01239_),
    .B2(_01337_),
    .C1(_01360_),
    .X(_01361_));
 sky130_fd_sc_hd__a31o_1 _04899_ (.A1(_01353_),
    .A2(_01357_),
    .A3(_01361_),
    .B1(_01341_),
    .X(_01362_));
 sky130_fd_sc_hd__nand4_1 _04900_ (.A(_01342_),
    .B(_01353_),
    .C(_01357_),
    .D(_01361_),
    .Y(_01363_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04901_ (.A(_01304_),
    .X(_01364_));
 sky130_fd_sc_hd__a21o_1 _04902_ (.A1(_01362_),
    .A2(_01363_),
    .B1(_01364_),
    .X(_01365_));
 sky130_fd_sc_hd__clkbuf_1 _04903_ (.A(_01304_),
    .X(_01366_));
 sky130_fd_sc_hd__xnor2_1 _04904_ (.A(_01290_),
    .B(_01280_),
    .Y(_01367_));
 sky130_fd_sc_hd__nand2_1 _04905_ (.A(_01366_),
    .B(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__a21oi_1 _04906_ (.A1(_01342_),
    .A2(_01303_),
    .B1(_01345_),
    .Y(_01369_));
 sky130_fd_sc_hd__clkbuf_1 _04907_ (.A(_01329_),
    .X(_01370_));
 sky130_fd_sc_hd__a21oi_1 _04908_ (.A1(_01333_),
    .A2(_01370_),
    .B1(_01325_),
    .Y(_01371_));
 sky130_fd_sc_hd__and3_1 _04909_ (.A(_01333_),
    .B(_01325_),
    .C(_01330_),
    .X(_01372_));
 sky130_fd_sc_hd__o211a_1 _04910_ (.A1(_01371_),
    .A2(_01372_),
    .B1(_01364_),
    .C1(_01370_),
    .X(_01373_));
 sky130_fd_sc_hd__a211oi_1 _04911_ (.A1(_01366_),
    .A2(_01370_),
    .B1(_01371_),
    .C1(_01372_),
    .Y(_01374_));
 sky130_fd_sc_hd__a2111o_1 _04912_ (.A1(_01365_),
    .A2(_01368_),
    .B1(_01369_),
    .C1(_01373_),
    .D1(_01374_),
    .X(_01375_));
 sky130_fd_sc_hd__clkbuf_1 _04913_ (.A(_01242_),
    .X(_01376_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04914_ (.A(_01376_),
    .X(_01377_));
 sky130_fd_sc_hd__nor2_1 _04915_ (.A(_01259_),
    .B(_01322_),
    .Y(_01378_));
 sky130_fd_sc_hd__o22a_1 _04916_ (.A1(_01248_),
    .A2(_01348_),
    .B1(_01378_),
    .B2(_01323_),
    .X(_01379_));
 sky130_fd_sc_hd__xnor2_1 _04917_ (.A(_01377_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__and3b_1 _04918_ (.A_N(_01347_),
    .B(_01327_),
    .C(_01328_),
    .X(_01381_));
 sky130_fd_sc_hd__nor2_1 _04919_ (.A(_01306_),
    .B(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hd__a22o_1 _04920_ (.A1(_01306_),
    .A2(_01380_),
    .B1(_01382_),
    .B2(_01370_),
    .X(_01383_));
 sky130_fd_sc_hd__or4_1 _04921_ (.A(_01320_),
    .B(_01352_),
    .C(_01375_),
    .D(_01383_),
    .X(_01384_));
 sky130_fd_sc_hd__clkbuf_1 _04922_ (.A(_01305_),
    .X(_01385_));
 sky130_fd_sc_hd__a31o_1 _04923_ (.A1(_01353_),
    .A2(_01357_),
    .A3(_01361_),
    .B1(_01293_),
    .X(_01386_));
 sky130_fd_sc_hd__clkbuf_1 _04924_ (.A(_01386_),
    .X(_01387_));
 sky130_fd_sc_hd__nand2_1 _04925_ (.A(_01385_),
    .B(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__or2_1 _04926_ (.A(_01281_),
    .B(_01284_),
    .X(_01389_));
 sky130_fd_sc_hd__nand2_1 _04927_ (.A(_01340_),
    .B(_01298_),
    .Y(_01390_));
 sky130_fd_sc_hd__o22a_1 _04928_ (.A1(_01296_),
    .A2(_01297_),
    .B1(_01343_),
    .B2(_01390_),
    .X(_01391_));
 sky130_fd_sc_hd__nand3_1 _04929_ (.A(_01389_),
    .B(_01387_),
    .C(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__a21o_1 _04930_ (.A1(_01387_),
    .A2(_01391_),
    .B1(_01389_),
    .X(_01393_));
 sky130_fd_sc_hd__o211a_1 _04931_ (.A1(_01325_),
    .A2(_01330_),
    .B1(_01334_),
    .C1(_01377_),
    .X(_01394_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04932_ (.A(_01286_),
    .X(_01395_));
 sky130_fd_sc_hd__inv_2 _04933_ (.A(_01215_),
    .Y(_01396_));
 sky130_fd_sc_hd__a21bo_1 _04934_ (.A1(_01189_),
    .A2(_01206_),
    .B1_N(_01310_),
    .X(_01397_));
 sky130_fd_sc_hd__xnor2_1 _04935_ (.A(_01396_),
    .B(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__o21ai_1 _04936_ (.A1(_01281_),
    .A2(_01395_),
    .B1(_01398_),
    .Y(_01399_));
 sky130_fd_sc_hd__a311o_1 _04937_ (.A1(_01333_),
    .A2(_01261_),
    .A3(_01330_),
    .B1(_01322_),
    .C1(_01376_),
    .X(_01400_));
 sky130_fd_sc_hd__or4b_1 _04938_ (.A(_01305_),
    .B(_01394_),
    .C(_01399_),
    .D_N(_01400_),
    .X(_01401_));
 sky130_fd_sc_hd__nor2_1 _04939_ (.A(_01348_),
    .B(_01249_),
    .Y(_01402_));
 sky130_fd_sc_hd__clkbuf_1 _04940_ (.A(_01236_),
    .X(_01403_));
 sky130_fd_sc_hd__o21ai_1 _04941_ (.A1(_01402_),
    .A2(_01265_),
    .B1(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__a21oi_1 _04942_ (.A1(_01310_),
    .A2(_01209_),
    .B1(_01224_),
    .Y(_01405_));
 sky130_fd_sc_hd__xnor2_1 _04943_ (.A(_01216_),
    .B(_01405_),
    .Y(_01406_));
 sky130_fd_sc_hd__o32a_1 _04944_ (.A1(_01236_),
    .A2(_01402_),
    .A3(_01265_),
    .B1(_01284_),
    .B2(_01395_),
    .X(_01407_));
 sky130_fd_sc_hd__nand4_1 _04945_ (.A(_01385_),
    .B(_01404_),
    .C(_01406_),
    .D(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__a32o_1 _04946_ (.A1(_01388_),
    .A2(_01392_),
    .A3(_01393_),
    .B1(_01401_),
    .B2(_01408_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _04947_ (.A0(_01316_),
    .A1(_01319_),
    .S(_01309_),
    .X(_01410_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04948_ (.A(_01254_),
    .X(_01411_));
 sky130_fd_sc_hd__a21oi_1 _04949_ (.A1(_01355_),
    .A2(_01276_),
    .B1(_01411_),
    .Y(_01412_));
 sky130_fd_sc_hd__o211ai_1 _04950_ (.A1(_01277_),
    .A2(_01412_),
    .B1(_01385_),
    .C1(_01403_),
    .Y(_01413_));
 sky130_fd_sc_hd__a211o_1 _04951_ (.A1(_01403_),
    .A2(_01364_),
    .B1(_01412_),
    .C1(_01277_),
    .X(_01414_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04952_ (.A(_01251_),
    .X(_01415_));
 sky130_fd_sc_hd__a21oi_1 _04953_ (.A1(_01359_),
    .A2(_01266_),
    .B1(_01271_),
    .Y(_01416_));
 sky130_fd_sc_hd__nor2_1 _04954_ (.A(_01272_),
    .B(_01416_),
    .Y(_01417_));
 sky130_fd_sc_hd__and3_1 _04955_ (.A(_01415_),
    .B(_01364_),
    .C(_01417_),
    .X(_01418_));
 sky130_fd_sc_hd__a21oi_1 _04956_ (.A1(_01415_),
    .A2(_01385_),
    .B1(_01417_),
    .Y(_01419_));
 sky130_fd_sc_hd__a211o_1 _04957_ (.A1(_01413_),
    .A2(_01414_),
    .B1(_01418_),
    .C1(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__and3_1 _04958_ (.A(_01285_),
    .B(_01386_),
    .C(_01391_),
    .X(_01421_));
 sky130_fd_sc_hd__a21oi_1 _04959_ (.A1(_01387_),
    .A2(_01391_),
    .B1(_01285_),
    .Y(_01422_));
 sky130_fd_sc_hd__clkbuf_1 _04960_ (.A(_01241_),
    .X(_01423_));
 sky130_fd_sc_hd__a21oi_1 _04961_ (.A1(_01335_),
    .A2(_01263_),
    .B1(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__a211oi_1 _04962_ (.A1(_01323_),
    .A2(_01366_),
    .B1(_01424_),
    .C1(_01264_),
    .Y(_01425_));
 sky130_fd_sc_hd__o211a_1 _04963_ (.A1(_01264_),
    .A2(_01424_),
    .B1(_01366_),
    .C1(_01323_),
    .X(_01426_));
 sky130_fd_sc_hd__o32a_1 _04964_ (.A1(_01388_),
    .A2(_01421_),
    .A3(_01422_),
    .B1(_01425_),
    .B2(_01426_),
    .X(_01427_));
 sky130_fd_sc_hd__or4b_1 _04965_ (.A(_01409_),
    .B(_01410_),
    .C(_01420_),
    .D_N(_01427_),
    .X(_01428_));
 sky130_fd_sc_hd__inv_2 _04966_ (.A(_01415_),
    .Y(_01429_));
 sky130_fd_sc_hd__o311a_1 _04967_ (.A1(_01403_),
    .A2(_01238_),
    .A3(_01338_),
    .B1(_01356_),
    .C1(_01354_),
    .X(_01430_));
 sky130_fd_sc_hd__xnor2_1 _04968_ (.A(_01429_),
    .B(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__xnor2_1 _04969_ (.A(_01339_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor4b_2 _04970_ (.A(_01308_),
    .B(_01384_),
    .C(_01428_),
    .D_N(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__a32o_1 _04971_ (.A1(\u_uart2wb.u_aut_det.state[3] ),
    .A2(_01166_),
    .A3(_01177_),
    .B1(_01433_),
    .B2(\u_uart2wb.u_aut_det.state[5] ),
    .X(_00011_));
 sky130_fd_sc_hd__nor2_1 _04972_ (.A(_01153_),
    .B(_01144_),
    .Y(_01434_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04973_ (.A(_01434_),
    .X(_01435_));
 sky130_fd_sc_hd__clkbuf_2 _04974_ (.A(_01435_),
    .X(_01436_));
 sky130_fd_sc_hd__and3_1 _04975_ (.A(\u_uart2wb.u_aut_det.state[0] ),
    .B(_01436_),
    .C(_01178_),
    .X(_01437_));
 sky130_fd_sc_hd__a31o_1 _04976_ (.A1(\u_uart2wb.u_aut_det.state[4] ),
    .A2(_01166_),
    .A3(_01177_),
    .B1(_01437_),
    .X(_00012_));
 sky130_fd_sc_hd__or2b_1 _04977_ (.A(\u_uart2wb.u_aut_det.rxd_sync[1] ),
    .B_N(\u_uart2wb.u_aut_det.rxd_sync[2] ),
    .X(_01438_));
 sky130_fd_sc_hd__clkbuf_1 _04978_ (.A(_01438_),
    .X(_01439_));
 sky130_fd_sc_hd__a32o_1 _04979_ (.A1(\u_uart2wb.u_aut_det.state[2] ),
    .A2(_01439_),
    .A3(_01177_),
    .B1(_01181_),
    .B2(\u_uart2wb.u_aut_det.state[4] ),
    .X(_00010_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04980_ (.A(_01175_),
    .X(_01440_));
 sky130_fd_sc_hd__a32o_1 _04981_ (.A1(\u_uart2wb.u_aut_det.state[1] ),
    .A2(_01439_),
    .A3(_01440_),
    .B1(_01181_),
    .B2(\u_uart2wb.u_aut_det.state[6] ),
    .X(_00009_));
 sky130_fd_sc_hd__and3_1 _04982_ (.A(\u_uart2wb.u_aut_det.clk_cnt[17] ),
    .B(_01167_),
    .C(_01174_),
    .X(_01441_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _04983_ (.A(_01441_),
    .X(_01442_));
 sky130_fd_sc_hd__or2_1 _04984_ (.A(\u_uart2wb.u_aut_det.state[2] ),
    .B(\u_uart2wb.u_aut_det.state[1] ),
    .X(_01443_));
 sky130_fd_sc_hd__or2_1 _04985_ (.A(\u_uart2wb.u_aut_det.state[6] ),
    .B(\u_uart2wb.u_aut_det.state[4] ),
    .X(_01444_));
 sky130_fd_sc_hd__or2_1 _04986_ (.A(\u_uart2wb.u_aut_det.state[3] ),
    .B(_01444_),
    .X(_01445_));
 sky130_fd_sc_hd__a22o_1 _04987_ (.A1(_01439_),
    .A2(_01443_),
    .B1(_01445_),
    .B2(_01166_),
    .X(_01446_));
 sky130_fd_sc_hd__o21a_1 _04988_ (.A1(_01157_),
    .A2(_01438_),
    .B1(\u_uart2wb.u_aut_det.state[0] ),
    .X(_01447_));
 sky130_fd_sc_hd__and2b_1 _04989_ (.A_N(_01433_),
    .B(\u_uart2wb.u_aut_det.state[5] ),
    .X(_01448_));
 sky130_fd_sc_hd__a211o_1 _04990_ (.A1(_01442_),
    .A2(_01446_),
    .B1(_01447_),
    .C1(_01448_),
    .X(_00008_));
 sky130_fd_sc_hd__and2_1 _04991_ (.A(\u_spi2wb.u_if.wr_phase ),
    .B(_01131_),
    .X(_01449_));
 sky130_fd_sc_hd__a31o_1 _04992_ (.A1(_01110_),
    .A2(_01112_),
    .A3(_01117_),
    .B1(_01449_),
    .X(_00002_));
 sky130_fd_sc_hd__clkbuf_1 _04993_ (.A(\u_spi2wb.u_if.spi_if_st[5] ),
    .X(_01450_));
 sky130_fd_sc_hd__nor2_1 _04994_ (.A(\u_spi2wb.u_if.ssn_l1 ),
    .B(_01117_),
    .Y(_01451_));
 sky130_fd_sc_hd__nand2_1 _04995_ (.A(_01450_),
    .B(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__o31a_1 _04996_ (.A1(\u_spi2wb.u_if.bitcnt[5] ),
    .A2(_01113_),
    .A3(_01126_),
    .B1(_01109_),
    .X(_01453_));
 sky130_fd_sc_hd__nand2_1 _04997_ (.A(_01120_),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__nand2_1 _04998_ (.A(_01452_),
    .B(_01454_),
    .Y(_00004_));
 sky130_fd_sc_hd__inv_2 _04999_ (.A(_01122_),
    .Y(_01455_));
 sky130_fd_sc_hd__nor2_1 _05000_ (.A(_01455_),
    .B(_01123_),
    .Y(_01456_));
 sky130_fd_sc_hd__and2_1 _05001_ (.A(\u_spi2wb.u_if.wr_phase ),
    .B(_01453_),
    .X(_01457_));
 sky130_fd_sc_hd__a21o_1 _05002_ (.A1(_01132_),
    .A2(_01456_),
    .B1(_01457_),
    .X(_00007_));
 sky130_fd_sc_hd__clkbuf_1 _05003_ (.A(_01122_),
    .X(_01458_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05004_ (.A(\u_spi2wb.u_if.ssn_l1 ),
    .X(_01459_));
 sky130_fd_sc_hd__nand2_1 _05005_ (.A(_01450_),
    .B(_01117_),
    .Y(_01460_));
 sky130_fd_sc_hd__nor2_1 _05006_ (.A(_01459_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__a31o_1 _05007_ (.A1(_01458_),
    .A2(_01121_),
    .A3(_01132_),
    .B1(_01461_),
    .X(_00006_));
 sky130_fd_sc_hd__a22o_1 _05008_ (.A1(\u_spi2wb.u_if.cmd_phase ),
    .A2(_01451_),
    .B1(_01453_),
    .B2(_01458_),
    .X(_00003_));
 sky130_fd_sc_hd__xnor2_1 _05009_ (.A(\u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ),
    .B(net332),
    .Y(_01462_));
 sky130_fd_sc_hd__xor2_1 _05010_ (.A(\u_async_wb.u_cmd_if.rd_ptr[0] ),
    .B(\u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ),
    .X(_01463_));
 sky130_fd_sc_hd__xnor2_1 _05011_ (.A(_01462_),
    .B(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__xnor2_1 _05012_ (.A(\u_async_wb.u_cmd_if.rd_ptr[1] ),
    .B(\u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ),
    .Y(_01465_));
 sky130_fd_sc_hd__nor2_1 _05013_ (.A(net332),
    .B(_01465_),
    .Y(_01466_));
 sky130_fd_sc_hd__mux2_1 _05014_ (.A0(net332),
    .A1(_01465_),
    .S(\u_async_wb.u_cmd_if.grey_rd_ptr[2] ),
    .X(_01467_));
 sky130_fd_sc_hd__or3_4 _05015_ (.A(_01464_),
    .B(_01466_),
    .C(net333),
    .X(_01468_));
 sky130_fd_sc_hd__mux4_1 _05016_ (.A0(\u_async_wb.u_cmd_if.mem[0][36] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][36] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][36] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][36] ),
    .S0(\u_async_wb.u_cmd_if.rd_ptr[0] ),
    .S1(net336),
    .X(_01469_));
 sky130_fd_sc_hd__and2_1 _05017_ (.A(net334),
    .B(net337),
    .X(_01470_));
 sky130_fd_sc_hd__clkbuf_2 _05018_ (.A(_01470_),
    .X(net214));
 sky130_fd_sc_hd__inv_2 _05019_ (.A(wbm_rst_i),
    .Y(\u_wbm_rst.arst_n ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05020_ (.A(\u_arb.gnt[1] ),
    .X(_01471_));
 sky130_fd_sc_hd__inv_2 _05021_ (.A(\u_arb.gnt[0] ),
    .Y(_01472_));
 sky130_fd_sc_hd__nor2_1 _05022_ (.A(_01472_),
    .B(\u_arb.gnt[1] ),
    .Y(_01473_));
 sky130_fd_sc_hd__nor2_1 _05023_ (.A(\u_arb.gnt[0] ),
    .B(\u_arb.gnt[1] ),
    .Y(_01474_));
 sky130_fd_sc_hd__and2_1 _05024_ (.A(wbm_adr_i[19]),
    .B(_01474_),
    .X(_01475_));
 sky130_fd_sc_hd__a221o_4 _05025_ (.A1(_01471_),
    .A2(\u_spi2wb.reg_addr[19] ),
    .B1(_01473_),
    .B2(\u_uart2wb.reg_addr[19] ),
    .C1(_01475_),
    .X(_01476_));
 sky130_fd_sc_hd__nand2_1 _05026_ (.A(wb_req),
    .B(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05027_ (.A(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__clkbuf_2 _05028_ (.A(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05029_ (.A(_01473_),
    .X(_01480_));
 sky130_fd_sc_hd__clkbuf_1 _05030_ (.A(\u_arb.gnt[1] ),
    .X(_01481_));
 sky130_fd_sc_hd__clkbuf_1 _05031_ (.A(_01474_),
    .X(_01482_));
 sky130_fd_sc_hd__a22o_1 _05032_ (.A1(_01481_),
    .A2(\u_spi2wb.reg_wr ),
    .B1(wbm_we_i),
    .B2(_01482_),
    .X(_01483_));
 sky130_fd_sc_hd__a21o_4 _05033_ (.A1(\u_uart2wb.reg_wr ),
    .A2(_01480_),
    .B1(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05034_ (.A(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__clkinv_2 _05035_ (.A(wb_req),
    .Y(_01486_));
 sky130_fd_sc_hd__or2_1 _05036_ (.A(_01486_),
    .B(_01476_),
    .X(_01487_));
 sky130_fd_sc_hd__xnor2_1 _05037_ (.A(\u_async_wb.u_cmd_if.sync_rd_ptr_1[1] ),
    .B(\u_async_wb.u_cmd_if.sync_rd_ptr[2] ),
    .Y(_01488_));
 sky130_fd_sc_hd__clkbuf_1 _05038_ (.A(\u_async_wb.u_cmd_if.wr_ptr[0] ),
    .X(_01489_));
 sky130_fd_sc_hd__clkbuf_1 _05039_ (.A(\u_async_wb.u_cmd_if.wr_ptr[1] ),
    .X(_01490_));
 sky130_fd_sc_hd__nor2_1 _05040_ (.A(_01489_),
    .B(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__and3b_1 _05041_ (.A_N(\u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ),
    .B(\u_async_wb.u_cmd_if.wr_ptr[1] ),
    .C(\u_async_wb.u_cmd_if.wr_ptr[0] ),
    .X(_01492_));
 sky130_fd_sc_hd__xnor2_1 _05042_ (.A(\u_async_wb.u_cmd_if.sync_rd_ptr[2] ),
    .B(\u_async_wb.u_cmd_if.grey_wr_ptr[2] ),
    .Y(_01493_));
 sky130_fd_sc_hd__mux2_1 _05043_ (.A0(_01491_),
    .A1(_01492_),
    .S(_01493_),
    .X(_01494_));
 sky130_fd_sc_hd__and2_1 _05044_ (.A(\u_async_wb.u_cmd_if.wr_ptr[0] ),
    .B(\u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ),
    .X(_01495_));
 sky130_fd_sc_hd__o21ai_1 _05045_ (.A1(_01488_),
    .A2(_01495_),
    .B1(_01490_),
    .Y(_01496_));
 sky130_fd_sc_hd__inv_2 _05046_ (.A(_01493_),
    .Y(_01497_));
 sky130_fd_sc_hd__o211a_1 _05047_ (.A1(_01490_),
    .A2(_01495_),
    .B1(_01496_),
    .C1(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__a211o_1 _05048_ (.A1(_01488_),
    .A2(_01494_),
    .B1(_01498_),
    .C1(\u_async_wb.PendingRd ),
    .X(_01499_));
 sky130_fd_sc_hd__nor2_1 _05049_ (.A(_01487_),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__clkbuf_1 _05050_ (.A(_01500_),
    .X(_01501_));
 sky130_fd_sc_hd__nand2_1 _05051_ (.A(_01485_),
    .B(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__and2_1 _05052_ (.A(\u_async_wb.u_resp_if.rd_ptr[1] ),
    .B(\u_async_wb.u_resp_if.sync_wr_ptr_1[1] ),
    .X(_01503_));
 sky130_fd_sc_hd__nor2_1 _05053_ (.A(\u_async_wb.u_resp_if.rd_ptr[1] ),
    .B(\u_async_wb.u_resp_if.sync_wr_ptr_1[1] ),
    .Y(_01504_));
 sky130_fd_sc_hd__xor2_1 _05054_ (.A(\u_async_wb.u_resp_if.rd_ptr[1] ),
    .B(\u_async_wb.u_resp_if.rd_ptr[0] ),
    .X(_01505_));
 sky130_fd_sc_hd__xnor2_1 _05055_ (.A(\u_async_wb.u_resp_if.sync_wr_ptr_1[0] ),
    .B(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__o21a_1 _05056_ (.A1(_01503_),
    .A2(_01504_),
    .B1(_01506_),
    .X(_01507_));
 sky130_fd_sc_hd__or3_1 _05057_ (.A(_01484_),
    .B(_01487_),
    .C(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__nor2_2 _05058_ (.A(\u_reg.reg_ack ),
    .B(_01478_),
    .Y(_00020_));
 sky130_fd_sc_hd__a31oi_4 _05059_ (.A1(_01479_),
    .A2(_01502_),
    .A3(_01508_),
    .B1(_00020_),
    .Y(_01509_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05060_ (.A(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__buf_2 _05061_ (.A(_01510_),
    .X(wb_ack_o1));
 sky130_fd_sc_hd__clkbuf_2 _05062_ (.A(wb_ack_o),
    .X(_01511_));
 sky130_fd_sc_hd__nor3b_1 _05063_ (.A(_01511_),
    .B(wb_ack_o1),
    .C_N(\u_delay2_stb2.X ),
    .Y(_00000_));
 sky130_fd_sc_hd__mux4_1 _05064_ (.A0(net307),
    .A1(net306),
    .A2(int_pll_clock),
    .A3(xtal_clk),
    .S0(\u_reg.cfg_clk_ctrl[0] ),
    .S1(\u_reg.cfg_clk_ctrl[1] ),
    .X(_01512_));
 sky130_fd_sc_hd__clkbuf_1 _05065_ (.A(_01512_),
    .X(\u_reg.u_wbs_ref_clkbuf.A ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05066_ (.A(\u_reg.cfg_clk_ctrl[3] ),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _05067_ (.A0(\u_reg.u_wbclk.clk_div_4 ),
    .A1(\u_reg.u_wbclk.clk_div_8 ),
    .S(\u_reg.cfg_clk_ctrl[2] ),
    .X(_01514_));
 sky130_fd_sc_hd__and2_1 _05068_ (.A(_01513_),
    .B(_01514_),
    .X(_01515_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05069_ (.A(\u_reg.cfg_clk_ctrl[2] ),
    .X(_01516_));
 sky130_fd_sc_hd__inv_2 _05070_ (.A(_01513_),
    .Y(_01517_));
 sky130_fd_sc_hd__and3b_1 _05071_ (.A_N(_01516_),
    .B(_01517_),
    .C(\u_reg.u_wbclk.mclk ),
    .X(_01518_));
 sky130_fd_sc_hd__a31o_1 _05072_ (.A1(_01516_),
    .A2(_01517_),
    .A3(\u_reg.u_wbclk.clk_div_2 ),
    .B1(\u_reg.force_refclk ),
    .X(_01519_));
 sky130_fd_sc_hd__inv_2 _05073_ (.A(\u_reg.force_refclk ),
    .Y(_01520_));
 sky130_fd_sc_hd__o32a_1 _05074_ (.A1(_01515_),
    .A2(_01518_),
    .A3(_01519_),
    .B1(_01520_),
    .B2(net307),
    .X(\u_reg.u_clkgate_wbs.CLK ));
 sky130_fd_sc_hd__mux4_1 _05075_ (.A0(net307),
    .A1(net306),
    .A2(int_pll_clock),
    .A3(xtal_clk),
    .S0(\u_reg.cfg_clk_ctrl[4] ),
    .S1(\u_reg.cfg_clk_ctrl[5] ),
    .X(_01521_));
 sky130_fd_sc_hd__clkbuf_1 _05076_ (.A(_01521_),
    .X(\u_reg.cpu_ref_clk_int ));
 sky130_fd_sc_hd__mux4_1 _05077_ (.A0(\u_reg.cpu_ref_clk ),
    .A1(\u_reg.cpu_ref_clk_div_2 ),
    .A2(\u_reg.cpu_ref_clk_div_4 ),
    .A3(\u_reg.cpu_ref_clk_div_8 ),
    .S0(_01516_),
    .S1(_01513_),
    .X(_01522_));
 sky130_fd_sc_hd__clkbuf_1 _05078_ (.A(_01522_),
    .X(\u_reg.cpu_clk_div ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05079_ (.A(net334),
    .X(_01523_));
 sky130_fd_sc_hd__clkbuf_2 _05080_ (.A(_01523_),
    .X(_01524_));
 sky130_fd_sc_hd__clkbuf_1 _05081_ (.A(_01524_),
    .X(_01525_));
 sky130_fd_sc_hd__clkbuf_2 _05082_ (.A(net340),
    .X(_01526_));
 sky130_fd_sc_hd__clkbuf_2 _05083_ (.A(_01526_),
    .X(_01527_));
 sky130_fd_sc_hd__clkbuf_2 _05084_ (.A(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__clkbuf_2 _05085_ (.A(net336),
    .X(_01529_));
 sky130_fd_sc_hd__clkbuf_2 _05086_ (.A(_01529_),
    .X(_01530_));
 sky130_fd_sc_hd__clkbuf_2 _05087_ (.A(_01530_),
    .X(_01531_));
 sky130_fd_sc_hd__mux4_1 _05088_ (.A0(\u_async_wb.u_cmd_if.mem[0][0] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][0] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][0] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][0] ),
    .S0(_01528_),
    .S1(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__and2_1 _05089_ (.A(_01525_),
    .B(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__clkbuf_2 _05090_ (.A(_01533_),
    .X(net209));
 sky130_fd_sc_hd__mux4_1 _05091_ (.A0(\u_async_wb.u_cmd_if.mem[0][1] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][1] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][1] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][1] ),
    .S0(_01528_),
    .S1(_01531_),
    .X(_01534_));
 sky130_fd_sc_hd__and2_1 _05092_ (.A(_01525_),
    .B(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05093_ (.A(_01535_),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 _05094_ (.A(_01527_),
    .X(_01536_));
 sky130_fd_sc_hd__mux4_1 _05095_ (.A0(\u_async_wb.u_cmd_if.mem[0][2] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][2] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][2] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][2] ),
    .S0(_01536_),
    .S1(_01531_),
    .X(_01537_));
 sky130_fd_sc_hd__and2_1 _05096_ (.A(_01525_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05097_ (.A(_01538_),
    .X(net211));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05098_ (.A(_01530_),
    .X(_01539_));
 sky130_fd_sc_hd__mux4_1 _05099_ (.A0(\u_async_wb.u_cmd_if.mem[0][3] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][3] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][3] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][3] ),
    .S0(_01536_),
    .S1(_01539_),
    .X(_01540_));
 sky130_fd_sc_hd__and2_1 _05100_ (.A(_01525_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__clkbuf_2 _05101_ (.A(_01541_),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 _05102_ (.A(_01524_),
    .X(_01542_));
 sky130_fd_sc_hd__mux4_1 _05103_ (.A0(\u_async_wb.u_cmd_if.mem[0][4] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][4] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][4] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][4] ),
    .S0(_01536_),
    .S1(_01539_),
    .X(_01543_));
 sky130_fd_sc_hd__and2_1 _05104_ (.A(_01542_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__clkbuf_1 _05105_ (.A(_01544_),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 _05106_ (.A0(\u_async_wb.u_cmd_if.mem[0][5] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][5] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][5] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][5] ),
    .S0(_01536_),
    .S1(_01539_),
    .X(_01545_));
 sky130_fd_sc_hd__and2_1 _05107_ (.A(_01542_),
    .B(_01545_),
    .X(_01546_));
 sky130_fd_sc_hd__clkbuf_1 _05108_ (.A(_01546_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 _05109_ (.A(_01526_),
    .X(_01547_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05110_ (.A(_01547_),
    .X(_01548_));
 sky130_fd_sc_hd__clkbuf_2 _05111_ (.A(_01548_),
    .X(_01549_));
 sky130_fd_sc_hd__mux4_1 _05112_ (.A0(\u_async_wb.u_cmd_if.mem[0][6] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][6] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][6] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][6] ),
    .S0(_01549_),
    .S1(_01539_),
    .X(_01550_));
 sky130_fd_sc_hd__and2_1 _05113_ (.A(_01542_),
    .B(_01550_),
    .X(_01551_));
 sky130_fd_sc_hd__clkbuf_1 _05114_ (.A(_01551_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 _05115_ (.A(_01529_),
    .X(_01552_));
 sky130_fd_sc_hd__clkbuf_2 _05116_ (.A(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05117_ (.A(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__mux4_1 _05118_ (.A0(\u_async_wb.u_cmd_if.mem[0][7] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][7] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][7] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][7] ),
    .S0(_01549_),
    .S1(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__and2_1 _05119_ (.A(_01542_),
    .B(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__clkbuf_1 _05120_ (.A(_01556_),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 _05121_ (.A(_01524_),
    .X(_01557_));
 sky130_fd_sc_hd__mux4_1 _05122_ (.A0(\u_async_wb.u_cmd_if.mem[0][8] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][8] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][8] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][8] ),
    .S0(_01549_),
    .S1(_01554_),
    .X(_01558_));
 sky130_fd_sc_hd__and2_1 _05123_ (.A(_01557_),
    .B(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__clkbuf_1 _05124_ (.A(_01559_),
    .X(net203));
 sky130_fd_sc_hd__mux4_2 _05125_ (.A0(\u_async_wb.u_cmd_if.mem[0][9] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][9] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][9] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][9] ),
    .S0(_01549_),
    .S1(_01554_),
    .X(_01560_));
 sky130_fd_sc_hd__and2_1 _05126_ (.A(_01557_),
    .B(_01560_),
    .X(_01561_));
 sky130_fd_sc_hd__clkbuf_1 _05127_ (.A(_01561_),
    .X(net204));
 sky130_fd_sc_hd__buf_2 _05128_ (.A(_01548_),
    .X(_01562_));
 sky130_fd_sc_hd__mux4_1 _05129_ (.A0(\u_async_wb.u_cmd_if.mem[0][10] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][10] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][10] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][10] ),
    .S0(_01562_),
    .S1(_01554_),
    .X(_01563_));
 sky130_fd_sc_hd__and2_1 _05130_ (.A(_01557_),
    .B(_01563_),
    .X(_01564_));
 sky130_fd_sc_hd__clkbuf_1 _05131_ (.A(_01564_),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 _05132_ (.A(_01553_),
    .X(_01565_));
 sky130_fd_sc_hd__mux4_1 _05133_ (.A0(\u_async_wb.u_cmd_if.mem[0][11] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][11] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][11] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][11] ),
    .S0(_01562_),
    .S1(_01565_),
    .X(_01566_));
 sky130_fd_sc_hd__and2_1 _05134_ (.A(_01557_),
    .B(_01566_),
    .X(_01567_));
 sky130_fd_sc_hd__clkbuf_1 _05135_ (.A(_01567_),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 _05136_ (.A(_01524_),
    .X(_01568_));
 sky130_fd_sc_hd__mux4_2 _05137_ (.A0(\u_async_wb.u_cmd_if.mem[0][12] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][12] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][12] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][12] ),
    .S0(_01562_),
    .S1(_01565_),
    .X(_01569_));
 sky130_fd_sc_hd__and2_1 _05138_ (.A(_01568_),
    .B(_01569_),
    .X(_01570_));
 sky130_fd_sc_hd__clkbuf_1 _05139_ (.A(_01570_),
    .X(net207));
 sky130_fd_sc_hd__mux4_2 _05140_ (.A0(\u_async_wb.u_cmd_if.mem[0][13] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][13] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][13] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][13] ),
    .S0(_01562_),
    .S1(_01565_),
    .X(_01571_));
 sky130_fd_sc_hd__and2_1 _05141_ (.A(_01568_),
    .B(_01571_),
    .X(_01572_));
 sky130_fd_sc_hd__clkbuf_1 _05142_ (.A(_01572_),
    .X(net208));
 sky130_fd_sc_hd__buf_2 _05143_ (.A(_01548_),
    .X(_01573_));
 sky130_fd_sc_hd__mux4_2 _05144_ (.A0(\u_async_wb.u_cmd_if.mem[0][14] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][14] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][14] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][14] ),
    .S0(_01573_),
    .S1(_01565_),
    .X(_01574_));
 sky130_fd_sc_hd__and2_1 _05145_ (.A(_01568_),
    .B(_01574_),
    .X(_01575_));
 sky130_fd_sc_hd__clkbuf_1 _05146_ (.A(_01575_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 _05147_ (.A(_01553_),
    .X(_01576_));
 sky130_fd_sc_hd__mux4_1 _05148_ (.A0(\u_async_wb.u_cmd_if.mem[0][15] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][15] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][15] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][15] ),
    .S0(_01573_),
    .S1(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__and2_1 _05149_ (.A(_01568_),
    .B(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__clkbuf_1 _05150_ (.A(_01578_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 _05151_ (.A(_01523_),
    .X(_01579_));
 sky130_fd_sc_hd__clkbuf_1 _05152_ (.A(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__mux4_2 _05153_ (.A0(\u_async_wb.u_cmd_if.mem[0][16] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][16] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][16] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][16] ),
    .S0(_01573_),
    .S1(_01576_),
    .X(_01581_));
 sky130_fd_sc_hd__and2_1 _05154_ (.A(_01580_),
    .B(_01581_),
    .X(_01582_));
 sky130_fd_sc_hd__clkbuf_1 _05155_ (.A(_01582_),
    .X(net180));
 sky130_fd_sc_hd__mux4_2 _05156_ (.A0(\u_async_wb.u_cmd_if.mem[0][17] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][17] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][17] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][17] ),
    .S0(_01573_),
    .S1(_01576_),
    .X(_01583_));
 sky130_fd_sc_hd__and2_1 _05157_ (.A(_01580_),
    .B(_01583_),
    .X(_01584_));
 sky130_fd_sc_hd__clkbuf_1 _05158_ (.A(_01584_),
    .X(net181));
 sky130_fd_sc_hd__buf_2 _05159_ (.A(_01548_),
    .X(_01585_));
 sky130_fd_sc_hd__mux4_2 _05160_ (.A0(\u_async_wb.u_cmd_if.mem[0][18] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][18] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][18] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][18] ),
    .S0(_01585_),
    .S1(_01576_),
    .X(_01586_));
 sky130_fd_sc_hd__and2_1 _05161_ (.A(_01580_),
    .B(_01586_),
    .X(_01587_));
 sky130_fd_sc_hd__clkbuf_1 _05162_ (.A(_01587_),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 _05163_ (.A(_01553_),
    .X(_01588_));
 sky130_fd_sc_hd__mux4_2 _05164_ (.A0(\u_async_wb.u_cmd_if.mem[0][19] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][19] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][19] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][19] ),
    .S0(_01585_),
    .S1(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__and2_1 _05165_ (.A(_01580_),
    .B(_01589_),
    .X(_01590_));
 sky130_fd_sc_hd__clkbuf_1 _05166_ (.A(_01590_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 _05167_ (.A(_01579_),
    .X(_01591_));
 sky130_fd_sc_hd__mux4_1 _05168_ (.A0(\u_async_wb.u_cmd_if.mem[0][20] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][20] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][20] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][20] ),
    .S0(_01585_),
    .S1(_01588_),
    .X(_01592_));
 sky130_fd_sc_hd__and2_1 _05169_ (.A(_01591_),
    .B(_01592_),
    .X(_01593_));
 sky130_fd_sc_hd__clkbuf_1 _05170_ (.A(_01593_),
    .X(net184));
 sky130_fd_sc_hd__mux4_1 _05171_ (.A0(\u_async_wb.u_cmd_if.mem[0][21] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][21] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][21] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][21] ),
    .S0(_01585_),
    .S1(_01588_),
    .X(_01594_));
 sky130_fd_sc_hd__and2_1 _05172_ (.A(_01591_),
    .B(_01594_),
    .X(_01595_));
 sky130_fd_sc_hd__clkbuf_1 _05173_ (.A(_01595_),
    .X(net185));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05174_ (.A(_01526_),
    .X(_01596_));
 sky130_fd_sc_hd__clkbuf_2 _05175_ (.A(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__mux4_1 _05176_ (.A0(\u_async_wb.u_cmd_if.mem[0][22] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][22] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][22] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][22] ),
    .S0(_01597_),
    .S1(_01588_),
    .X(_01598_));
 sky130_fd_sc_hd__and2_1 _05177_ (.A(_01591_),
    .B(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__clkbuf_1 _05178_ (.A(_01599_),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 _05179_ (.A(_01529_),
    .X(_01600_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05180_ (.A(_01600_),
    .X(_01601_));
 sky130_fd_sc_hd__mux4_1 _05181_ (.A0(\u_async_wb.u_cmd_if.mem[0][23] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][23] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][23] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][23] ),
    .S0(_01597_),
    .S1(_01601_),
    .X(_01602_));
 sky130_fd_sc_hd__and2_1 _05182_ (.A(_01591_),
    .B(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__clkbuf_1 _05183_ (.A(_01603_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 _05184_ (.A(_01579_),
    .X(_01604_));
 sky130_fd_sc_hd__mux4_1 _05185_ (.A0(\u_async_wb.u_cmd_if.mem[0][24] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][24] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][24] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][24] ),
    .S0(_01597_),
    .S1(_01601_),
    .X(_01605_));
 sky130_fd_sc_hd__and2_1 _05186_ (.A(_01604_),
    .B(_01605_),
    .X(_01606_));
 sky130_fd_sc_hd__clkbuf_1 _05187_ (.A(_01606_),
    .X(net189));
 sky130_fd_sc_hd__mux4_1 _05188_ (.A0(\u_async_wb.u_cmd_if.mem[0][25] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][25] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][25] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][25] ),
    .S0(_01597_),
    .S1(_01601_),
    .X(_01607_));
 sky130_fd_sc_hd__and2_1 _05189_ (.A(_01604_),
    .B(_01607_),
    .X(_01608_));
 sky130_fd_sc_hd__clkbuf_1 _05190_ (.A(_01608_),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 _05191_ (.A(_01596_),
    .X(_01609_));
 sky130_fd_sc_hd__mux4_1 _05192_ (.A0(\u_async_wb.u_cmd_if.mem[0][26] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][26] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][26] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][26] ),
    .S0(_01609_),
    .S1(_01601_),
    .X(_01610_));
 sky130_fd_sc_hd__and2_1 _05193_ (.A(_01604_),
    .B(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__clkbuf_1 _05194_ (.A(_01611_),
    .X(net191));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05195_ (.A(_01600_),
    .X(_01612_));
 sky130_fd_sc_hd__mux4_1 _05196_ (.A0(\u_async_wb.u_cmd_if.mem[0][27] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][27] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][27] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][27] ),
    .S0(_01609_),
    .S1(_01612_),
    .X(_01613_));
 sky130_fd_sc_hd__and2_1 _05197_ (.A(_01604_),
    .B(_01613_),
    .X(_01614_));
 sky130_fd_sc_hd__clkbuf_1 _05198_ (.A(_01614_),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 _05199_ (.A(_01579_),
    .X(_01615_));
 sky130_fd_sc_hd__mux4_1 _05200_ (.A0(\u_async_wb.u_cmd_if.mem[0][28] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][28] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][28] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][28] ),
    .S0(_01609_),
    .S1(_01612_),
    .X(_01616_));
 sky130_fd_sc_hd__and2_1 _05201_ (.A(_01615_),
    .B(_01616_),
    .X(_01617_));
 sky130_fd_sc_hd__clkbuf_1 _05202_ (.A(_01617_),
    .X(net193));
 sky130_fd_sc_hd__mux4_1 _05203_ (.A0(\u_async_wb.u_cmd_if.mem[0][29] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][29] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][29] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][29] ),
    .S0(_01609_),
    .S1(_01612_),
    .X(_01618_));
 sky130_fd_sc_hd__and2_1 _05204_ (.A(_01615_),
    .B(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__clkbuf_1 _05205_ (.A(_01619_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 _05206_ (.A(_01596_),
    .X(_01620_));
 sky130_fd_sc_hd__mux4_1 _05207_ (.A0(\u_async_wb.u_cmd_if.mem[0][30] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][30] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][30] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][30] ),
    .S0(_01620_),
    .S1(_01612_),
    .X(_01621_));
 sky130_fd_sc_hd__and2_1 _05208_ (.A(_01615_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__clkbuf_1 _05209_ (.A(_01622_),
    .X(net195));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05210_ (.A(_01600_),
    .X(_01623_));
 sky130_fd_sc_hd__mux4_1 _05211_ (.A0(\u_async_wb.u_cmd_if.mem[0][31] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][31] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][31] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][31] ),
    .S0(_01620_),
    .S1(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__and2_1 _05212_ (.A(_01615_),
    .B(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__clkbuf_1 _05213_ (.A(_01625_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 _05214_ (.A(_01523_),
    .X(_01626_));
 sky130_fd_sc_hd__clkbuf_1 _05215_ (.A(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__mux4_1 _05216_ (.A0(\u_async_wb.u_cmd_if.mem[0][32] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][32] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][32] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][32] ),
    .S0(_01620_),
    .S1(_01623_),
    .X(_01628_));
 sky130_fd_sc_hd__and2_1 _05217_ (.A(_01627_),
    .B(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__clkbuf_1 _05218_ (.A(_01629_),
    .X(net197));
 sky130_fd_sc_hd__mux4_1 _05219_ (.A0(\u_async_wb.u_cmd_if.mem[0][33] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][33] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][33] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][33] ),
    .S0(_01620_),
    .S1(_01623_),
    .X(_01630_));
 sky130_fd_sc_hd__and2_1 _05220_ (.A(_01627_),
    .B(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__clkbuf_1 _05221_ (.A(_01631_),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 _05222_ (.A(_01596_),
    .X(_01632_));
 sky130_fd_sc_hd__mux4_1 _05223_ (.A0(\u_async_wb.u_cmd_if.mem[0][34] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][34] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][34] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][34] ),
    .S0(_01632_),
    .S1(_01623_),
    .X(_01633_));
 sky130_fd_sc_hd__and2_1 _05224_ (.A(_01627_),
    .B(_01633_),
    .X(_01634_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05225_ (.A(_01634_),
    .X(net200));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05226_ (.A(_01600_),
    .X(_01635_));
 sky130_fd_sc_hd__mux4_1 _05227_ (.A0(\u_async_wb.u_cmd_if.mem[0][35] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][35] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][35] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][35] ),
    .S0(_01632_),
    .S1(_01635_),
    .X(_01636_));
 sky130_fd_sc_hd__and2_1 _05228_ (.A(_01627_),
    .B(_01636_),
    .X(_01637_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05229_ (.A(_01637_),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 _05230_ (.A(_01626_),
    .X(_01638_));
 sky130_fd_sc_hd__mux4_1 _05231_ (.A0(\u_async_wb.u_cmd_if.mem[0][37] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][37] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][37] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][37] ),
    .S0(_01632_),
    .S1(_01635_),
    .X(_01639_));
 sky130_fd_sc_hd__and2_1 _05232_ (.A(_01638_),
    .B(_01639_),
    .X(_01640_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05233_ (.A(_01640_),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 _05234_ (.A0(\u_async_wb.u_cmd_if.mem[0][38] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][38] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][38] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][38] ),
    .S0(_01632_),
    .S1(_01635_),
    .X(_01641_));
 sky130_fd_sc_hd__and2_1 _05235_ (.A(_01638_),
    .B(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05236_ (.A(_01642_),
    .X(net154));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05237_ (.A(_01526_),
    .X(_01643_));
 sky130_fd_sc_hd__clkbuf_2 _05238_ (.A(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__mux4_1 _05239_ (.A0(\u_async_wb.u_cmd_if.mem[0][39] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][39] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][39] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][39] ),
    .S0(_01644_),
    .S1(_01635_),
    .X(_01645_));
 sky130_fd_sc_hd__and2_1 _05240_ (.A(_01638_),
    .B(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05241_ (.A(_01646_),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 _05242_ (.A(_01529_),
    .X(_01647_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05243_ (.A(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__mux4_1 _05244_ (.A0(\u_async_wb.u_cmd_if.mem[0][40] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][40] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][40] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][40] ),
    .S0(_01644_),
    .S1(_01648_),
    .X(_01649_));
 sky130_fd_sc_hd__and2_1 _05245_ (.A(_01638_),
    .B(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05246_ (.A(_01650_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 _05247_ (.A(_01626_),
    .X(_01651_));
 sky130_fd_sc_hd__mux4_1 _05248_ (.A0(\u_async_wb.u_cmd_if.mem[0][41] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][41] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][41] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][41] ),
    .S0(_01644_),
    .S1(_01648_),
    .X(_01652_));
 sky130_fd_sc_hd__and2_1 _05249_ (.A(_01651_),
    .B(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05250_ (.A(_01653_),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 _05251_ (.A0(\u_async_wb.u_cmd_if.mem[0][42] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][42] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][42] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][42] ),
    .S0(_01644_),
    .S1(_01648_),
    .X(_01654_));
 sky130_fd_sc_hd__and2_1 _05252_ (.A(_01651_),
    .B(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05253_ (.A(_01655_),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 _05254_ (.A(_01643_),
    .X(_01656_));
 sky130_fd_sc_hd__mux4_1 _05255_ (.A0(\u_async_wb.u_cmd_if.mem[0][43] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][43] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][43] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][43] ),
    .S0(_01656_),
    .S1(_01648_),
    .X(_01657_));
 sky130_fd_sc_hd__and2_1 _05256_ (.A(_01651_),
    .B(_01657_),
    .X(_01658_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05257_ (.A(_01658_),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 _05258_ (.A(_01647_),
    .X(_01659_));
 sky130_fd_sc_hd__mux4_2 _05259_ (.A0(\u_async_wb.u_cmd_if.mem[0][44] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][44] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][44] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][44] ),
    .S0(_01656_),
    .S1(_01659_),
    .X(_01660_));
 sky130_fd_sc_hd__and2_1 _05260_ (.A(_01651_),
    .B(_01660_),
    .X(_01661_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05261_ (.A(_01661_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 _05262_ (.A(_01626_),
    .X(_01662_));
 sky130_fd_sc_hd__mux4_2 _05263_ (.A0(\u_async_wb.u_cmd_if.mem[0][45] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][45] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][45] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][45] ),
    .S0(_01656_),
    .S1(_01659_),
    .X(_01663_));
 sky130_fd_sc_hd__and2_1 _05264_ (.A(_01662_),
    .B(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05265_ (.A(_01664_),
    .X(net173));
 sky130_fd_sc_hd__mux4_2 _05266_ (.A0(\u_async_wb.u_cmd_if.mem[0][46] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][46] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][46] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][46] ),
    .S0(_01656_),
    .S1(_01659_),
    .X(_01665_));
 sky130_fd_sc_hd__and2_1 _05267_ (.A(_01662_),
    .B(_01665_),
    .X(_01666_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05268_ (.A(_01666_),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 _05269_ (.A(_01643_),
    .X(_01667_));
 sky130_fd_sc_hd__mux4_2 _05270_ (.A0(\u_async_wb.u_cmd_if.mem[0][47] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][47] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][47] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][47] ),
    .S0(_01667_),
    .S1(_01659_),
    .X(_01668_));
 sky130_fd_sc_hd__and2_1 _05271_ (.A(_01662_),
    .B(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05272_ (.A(_01669_),
    .X(net144));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05273_ (.A(_01647_),
    .X(_01670_));
 sky130_fd_sc_hd__mux4_2 _05274_ (.A0(\u_async_wb.u_cmd_if.mem[0][48] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][48] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][48] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][48] ),
    .S0(_01667_),
    .S1(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__and2_1 _05275_ (.A(_01662_),
    .B(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05276_ (.A(_01672_),
    .X(net145));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05277_ (.A(net334),
    .X(_01673_));
 sky130_fd_sc_hd__clkbuf_1 _05278_ (.A(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_1 _05279_ (.A0(\u_async_wb.u_cmd_if.mem[0][49] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][49] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][49] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][49] ),
    .S0(_01667_),
    .S1(_01670_),
    .X(_01675_));
 sky130_fd_sc_hd__and2_1 _05280_ (.A(_01674_),
    .B(_01675_),
    .X(_01676_));
 sky130_fd_sc_hd__clkbuf_2 _05281_ (.A(_01676_),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 _05282_ (.A0(\u_async_wb.u_cmd_if.mem[0][50] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][50] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][50] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][50] ),
    .S0(_01667_),
    .S1(_01670_),
    .X(_01677_));
 sky130_fd_sc_hd__and2_1 _05283_ (.A(_01674_),
    .B(_01677_),
    .X(_01678_));
 sky130_fd_sc_hd__clkbuf_2 _05284_ (.A(_01678_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 _05285_ (.A(_01643_),
    .X(_01679_));
 sky130_fd_sc_hd__mux4_1 _05286_ (.A0(\u_async_wb.u_cmd_if.mem[0][51] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][51] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][51] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][51] ),
    .S0(_01679_),
    .S1(_01670_),
    .X(_01680_));
 sky130_fd_sc_hd__and2_1 _05287_ (.A(_01674_),
    .B(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__clkbuf_2 _05288_ (.A(_01681_),
    .X(net148));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05289_ (.A(_01647_),
    .X(_01682_));
 sky130_fd_sc_hd__mux4_1 _05290_ (.A0(\u_async_wb.u_cmd_if.mem[0][52] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][52] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][52] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][52] ),
    .S0(_01679_),
    .S1(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__and2_1 _05291_ (.A(_01674_),
    .B(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__clkbuf_2 _05292_ (.A(_01684_),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _05293_ (.A(_01673_),
    .X(_01685_));
 sky130_fd_sc_hd__mux4_1 _05294_ (.A0(\u_async_wb.u_cmd_if.mem[0][53] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][53] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][53] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][53] ),
    .S0(_01679_),
    .S1(_01682_),
    .X(_01686_));
 sky130_fd_sc_hd__and2_1 _05295_ (.A(_01685_),
    .B(_01686_),
    .X(_01687_));
 sky130_fd_sc_hd__clkbuf_1 _05296_ (.A(_01687_),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 _05297_ (.A0(\u_async_wb.u_cmd_if.mem[0][54] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][54] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][54] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][54] ),
    .S0(_01679_),
    .S1(_01682_),
    .X(_01688_));
 sky130_fd_sc_hd__and2_1 _05298_ (.A(_01685_),
    .B(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05299_ (.A(_01689_),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 _05300_ (.A(_01547_),
    .X(_01690_));
 sky130_fd_sc_hd__mux4_1 _05301_ (.A0(\u_async_wb.u_cmd_if.mem[0][55] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][55] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][55] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][55] ),
    .S0(_01690_),
    .S1(_01682_),
    .X(_01691_));
 sky130_fd_sc_hd__and2_1 _05302_ (.A(_01685_),
    .B(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05303_ (.A(_01692_),
    .X(net152));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05304_ (.A(_01552_),
    .X(_01693_));
 sky130_fd_sc_hd__mux4_1 _05305_ (.A0(\u_async_wb.u_cmd_if.mem[0][56] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][56] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][56] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][56] ),
    .S0(_01690_),
    .S1(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__and2_1 _05306_ (.A(_01685_),
    .B(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05307_ (.A(_01695_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _05308_ (.A(_01673_),
    .X(_01696_));
 sky130_fd_sc_hd__mux4_1 _05309_ (.A0(\u_async_wb.u_cmd_if.mem[0][57] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][57] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][57] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][57] ),
    .S0(_01690_),
    .S1(_01693_),
    .X(_01697_));
 sky130_fd_sc_hd__and2_1 _05310_ (.A(_01696_),
    .B(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__clkbuf_1 _05311_ (.A(_01698_),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 _05312_ (.A0(\u_async_wb.u_cmd_if.mem[0][58] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][58] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][58] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][58] ),
    .S0(_01690_),
    .S1(_01693_),
    .X(_01699_));
 sky130_fd_sc_hd__and2_1 _05313_ (.A(_01696_),
    .B(_01699_),
    .X(_01700_));
 sky130_fd_sc_hd__clkbuf_1 _05314_ (.A(_01700_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 _05315_ (.A(_01547_),
    .X(_01701_));
 sky130_fd_sc_hd__mux4_1 _05316_ (.A0(\u_async_wb.u_cmd_if.mem[0][59] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][59] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][59] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][59] ),
    .S0(_01701_),
    .S1(_01693_),
    .X(_01702_));
 sky130_fd_sc_hd__and2_1 _05317_ (.A(_01696_),
    .B(_01702_),
    .X(_01703_));
 sky130_fd_sc_hd__clkbuf_1 _05318_ (.A(_01703_),
    .X(net157));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05319_ (.A(_01552_),
    .X(_01704_));
 sky130_fd_sc_hd__mux4_1 _05320_ (.A0(\u_async_wb.u_cmd_if.mem[0][60] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][60] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][60] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][60] ),
    .S0(_01701_),
    .S1(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__and2_1 _05321_ (.A(_01696_),
    .B(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__clkbuf_1 _05322_ (.A(_01706_),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 _05323_ (.A(_01673_),
    .X(_01707_));
 sky130_fd_sc_hd__mux4_1 _05324_ (.A0(\u_async_wb.u_cmd_if.mem[0][61] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][61] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][61] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][61] ),
    .S0(_01701_),
    .S1(_01704_),
    .X(_01708_));
 sky130_fd_sc_hd__and2_1 _05325_ (.A(_01707_),
    .B(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__clkbuf_1 _05326_ (.A(_01709_),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 _05327_ (.A0(\u_async_wb.u_cmd_if.mem[0][62] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][62] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][62] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][62] ),
    .S0(_01701_),
    .S1(_01704_),
    .X(_01710_));
 sky130_fd_sc_hd__and2_1 _05328_ (.A(_01707_),
    .B(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__clkbuf_1 _05329_ (.A(_01711_),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 _05330_ (.A(_01547_),
    .X(_01712_));
 sky130_fd_sc_hd__mux4_1 _05331_ (.A0(\u_async_wb.u_cmd_if.mem[0][63] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][63] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][63] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][63] ),
    .S0(_01712_),
    .S1(_01704_),
    .X(_01713_));
 sky130_fd_sc_hd__and2_1 _05332_ (.A(_01707_),
    .B(_01713_),
    .X(_01714_));
 sky130_fd_sc_hd__clkbuf_1 _05333_ (.A(_01714_),
    .X(net161));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05334_ (.A(_01552_),
    .X(_01715_));
 sky130_fd_sc_hd__mux4_1 _05335_ (.A0(\u_async_wb.u_cmd_if.mem[0][64] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][64] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][64] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][64] ),
    .S0(_01712_),
    .S1(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__and2_1 _05336_ (.A(_01707_),
    .B(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__clkbuf_1 _05337_ (.A(_01717_),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 _05338_ (.A(_01523_),
    .X(_01718_));
 sky130_fd_sc_hd__mux4_1 _05339_ (.A0(\u_async_wb.u_cmd_if.mem[0][65] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][65] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][65] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][65] ),
    .S0(_01712_),
    .S1(_01715_),
    .X(_01719_));
 sky130_fd_sc_hd__and2_1 _05340_ (.A(_01718_),
    .B(_01719_),
    .X(_01720_));
 sky130_fd_sc_hd__clkbuf_1 _05341_ (.A(_01720_),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 _05342_ (.A0(\u_async_wb.u_cmd_if.mem[0][66] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][66] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][66] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][66] ),
    .S0(_01712_),
    .S1(_01715_),
    .X(_01721_));
 sky130_fd_sc_hd__and2_1 _05343_ (.A(_01718_),
    .B(_01721_),
    .X(_01722_));
 sky130_fd_sc_hd__clkbuf_1 _05344_ (.A(_01722_),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 _05345_ (.A0(\u_async_wb.u_cmd_if.mem[0][67] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][67] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][67] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][67] ),
    .S0(_01527_),
    .S1(_01715_),
    .X(_01723_));
 sky130_fd_sc_hd__and2_1 _05346_ (.A(_01718_),
    .B(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__clkbuf_1 _05347_ (.A(_01724_),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 _05348_ (.A0(\u_async_wb.u_cmd_if.mem[0][68] ),
    .A1(\u_async_wb.u_cmd_if.mem[1][68] ),
    .A2(\u_async_wb.u_cmd_if.mem[2][68] ),
    .A3(\u_async_wb.u_cmd_if.mem[3][68] ),
    .S0(_01527_),
    .S1(_01530_),
    .X(_01725_));
 sky130_fd_sc_hd__and2_1 _05349_ (.A(_01718_),
    .B(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__clkbuf_1 _05350_ (.A(_01726_),
    .X(net167));
 sky130_fd_sc_hd__and2b_1 _05351_ (.A_N(net330),
    .B(_01468_),
    .X(_01727_));
 sky130_fd_sc_hd__clkbuf_2 _05352_ (.A(net331),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 _05353_ (.A(_01481_),
    .X(_01728_));
 sky130_fd_sc_hd__clkbuf_1 _05354_ (.A(_01728_),
    .X(_01729_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05355_ (.A(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__clkbuf_2 _05356_ (.A(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__nor2_1 _05357_ (.A(\u_spi2wb.reg_wr ),
    .B(\u_spi2wb.reg_rd ),
    .Y(_01732_));
 sky130_fd_sc_hd__inv_2 _05358_ (.A(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__clkbuf_1 _05359_ (.A(_01482_),
    .X(_01734_));
 sky130_fd_sc_hd__clkbuf_1 _05360_ (.A(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__clkbuf_2 _05361_ (.A(_01735_),
    .X(_01736_));
 sky130_fd_sc_hd__clkbuf_1 _05362_ (.A(_01480_),
    .X(_01737_));
 sky130_fd_sc_hd__clkbuf_1 _05363_ (.A(_01737_),
    .X(_01738_));
 sky130_fd_sc_hd__clkbuf_2 _05364_ (.A(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__a32o_1 _05365_ (.A1(wbm_cyc_i),
    .A2(wbm_stb_i),
    .A3(_01736_),
    .B1(_01739_),
    .B2(\u_uart2wb.u_async_reg_bus.out_reg_cs ),
    .X(_01740_));
 sky130_fd_sc_hd__a21o_1 _05366_ (.A1(_01731_),
    .A2(_01733_),
    .B1(_01740_),
    .X(\u_delay1_stb0.A ));
 sky130_fd_sc_hd__clkbuf_1 _05367_ (.A(_01736_),
    .X(_01741_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05368_ (.A(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__clkbuf_1 _05369_ (.A(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__and2_1 _05370_ (.A(\wb_dat_o[0] ),
    .B(_01743_),
    .X(_01744_));
 sky130_fd_sc_hd__clkbuf_1 _05371_ (.A(_01744_),
    .X(net110));
 sky130_fd_sc_hd__and2_1 _05372_ (.A(\wb_dat_o[1] ),
    .B(_01743_),
    .X(_01745_));
 sky130_fd_sc_hd__clkbuf_1 _05373_ (.A(_01745_),
    .X(net121));
 sky130_fd_sc_hd__and2_1 _05374_ (.A(\wb_dat_o[2] ),
    .B(_01743_),
    .X(_01746_));
 sky130_fd_sc_hd__clkbuf_1 _05375_ (.A(_01746_),
    .X(net132));
 sky130_fd_sc_hd__and2_1 _05376_ (.A(\wb_dat_o[3] ),
    .B(_01743_),
    .X(_01747_));
 sky130_fd_sc_hd__clkbuf_1 _05377_ (.A(_01747_),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 _05378_ (.A(_01742_),
    .X(_01748_));
 sky130_fd_sc_hd__and2_1 _05379_ (.A(\wb_dat_o[4] ),
    .B(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__clkbuf_1 _05380_ (.A(_01749_),
    .X(net136));
 sky130_fd_sc_hd__and2_1 _05381_ (.A(\wb_dat_o[5] ),
    .B(_01748_),
    .X(_01750_));
 sky130_fd_sc_hd__clkbuf_1 _05382_ (.A(_01750_),
    .X(net137));
 sky130_fd_sc_hd__and2_1 _05383_ (.A(\wb_dat_o[6] ),
    .B(_01748_),
    .X(_01751_));
 sky130_fd_sc_hd__clkbuf_1 _05384_ (.A(_01751_),
    .X(net138));
 sky130_fd_sc_hd__and2_1 _05385_ (.A(\wb_dat_o[7] ),
    .B(_01748_),
    .X(_01752_));
 sky130_fd_sc_hd__clkbuf_1 _05386_ (.A(_01752_),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 _05387_ (.A(_01741_),
    .X(_01753_));
 sky130_fd_sc_hd__clkbuf_1 _05388_ (.A(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__and2_1 _05389_ (.A(\wb_dat_o[8] ),
    .B(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__clkbuf_1 _05390_ (.A(_01755_),
    .X(net140));
 sky130_fd_sc_hd__and2_1 _05391_ (.A(\wb_dat_o[9] ),
    .B(_01754_),
    .X(_01756_));
 sky130_fd_sc_hd__clkbuf_1 _05392_ (.A(_01756_),
    .X(net141));
 sky130_fd_sc_hd__and2_1 _05393_ (.A(\wb_dat_o[10] ),
    .B(_01754_),
    .X(_01757_));
 sky130_fd_sc_hd__clkbuf_1 _05394_ (.A(_01757_),
    .X(net111));
 sky130_fd_sc_hd__and2_1 _05395_ (.A(\wb_dat_o[11] ),
    .B(_01754_),
    .X(_01758_));
 sky130_fd_sc_hd__clkbuf_1 _05396_ (.A(_01758_),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 _05397_ (.A(_01753_),
    .X(_01759_));
 sky130_fd_sc_hd__and2_1 _05398_ (.A(\wb_dat_o[12] ),
    .B(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__clkbuf_1 _05399_ (.A(_01760_),
    .X(net113));
 sky130_fd_sc_hd__and2_1 _05400_ (.A(\wb_dat_o[13] ),
    .B(_01759_),
    .X(_01761_));
 sky130_fd_sc_hd__clkbuf_1 _05401_ (.A(_01761_),
    .X(net114));
 sky130_fd_sc_hd__and2_1 _05402_ (.A(\wb_dat_o[14] ),
    .B(_01759_),
    .X(_01762_));
 sky130_fd_sc_hd__clkbuf_1 _05403_ (.A(_01762_),
    .X(net115));
 sky130_fd_sc_hd__and2_1 _05404_ (.A(\wb_dat_o[15] ),
    .B(_01759_),
    .X(_01763_));
 sky130_fd_sc_hd__clkbuf_1 _05405_ (.A(_01763_),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 _05406_ (.A(_01753_),
    .X(_01764_));
 sky130_fd_sc_hd__and2_1 _05407_ (.A(\wb_dat_o[16] ),
    .B(_01764_),
    .X(_01765_));
 sky130_fd_sc_hd__clkbuf_1 _05408_ (.A(_01765_),
    .X(net117));
 sky130_fd_sc_hd__and2_1 _05409_ (.A(\wb_dat_o[17] ),
    .B(_01764_),
    .X(_01766_));
 sky130_fd_sc_hd__clkbuf_1 _05410_ (.A(_01766_),
    .X(net118));
 sky130_fd_sc_hd__and2_1 _05411_ (.A(\wb_dat_o[18] ),
    .B(_01764_),
    .X(_01767_));
 sky130_fd_sc_hd__clkbuf_1 _05412_ (.A(_01767_),
    .X(net119));
 sky130_fd_sc_hd__and2_1 _05413_ (.A(\wb_dat_o[19] ),
    .B(_01764_),
    .X(_01768_));
 sky130_fd_sc_hd__clkbuf_1 _05414_ (.A(_01768_),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 _05415_ (.A(_01753_),
    .X(_01769_));
 sky130_fd_sc_hd__and2_1 _05416_ (.A(\wb_dat_o[20] ),
    .B(_01769_),
    .X(_01770_));
 sky130_fd_sc_hd__clkbuf_1 _05417_ (.A(_01770_),
    .X(net122));
 sky130_fd_sc_hd__and2_1 _05418_ (.A(\wb_dat_o[21] ),
    .B(_01769_),
    .X(_01771_));
 sky130_fd_sc_hd__clkbuf_1 _05419_ (.A(_01771_),
    .X(net123));
 sky130_fd_sc_hd__and2_1 _05420_ (.A(\wb_dat_o[22] ),
    .B(_01769_),
    .X(_01772_));
 sky130_fd_sc_hd__clkbuf_1 _05421_ (.A(_01772_),
    .X(net124));
 sky130_fd_sc_hd__and2_1 _05422_ (.A(\wb_dat_o[23] ),
    .B(_01769_),
    .X(_01773_));
 sky130_fd_sc_hd__clkbuf_1 _05423_ (.A(_01773_),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 _05424_ (.A(_01734_),
    .X(_01774_));
 sky130_fd_sc_hd__clkbuf_2 _05425_ (.A(_01774_),
    .X(_01775_));
 sky130_fd_sc_hd__clkbuf_2 _05426_ (.A(_01775_),
    .X(_01776_));
 sky130_fd_sc_hd__clkbuf_1 _05427_ (.A(_01776_),
    .X(_01777_));
 sky130_fd_sc_hd__and2_1 _05428_ (.A(\wb_dat_o[24] ),
    .B(_01777_),
    .X(_01778_));
 sky130_fd_sc_hd__clkbuf_1 _05429_ (.A(_01778_),
    .X(net126));
 sky130_fd_sc_hd__and2_1 _05430_ (.A(\wb_dat_o[25] ),
    .B(_01777_),
    .X(_01779_));
 sky130_fd_sc_hd__clkbuf_1 _05431_ (.A(_01779_),
    .X(net127));
 sky130_fd_sc_hd__and2_1 _05432_ (.A(\wb_dat_o[26] ),
    .B(_01777_),
    .X(_01780_));
 sky130_fd_sc_hd__clkbuf_1 _05433_ (.A(_01780_),
    .X(net128));
 sky130_fd_sc_hd__and2_1 _05434_ (.A(\wb_dat_o[27] ),
    .B(_01777_),
    .X(_01781_));
 sky130_fd_sc_hd__clkbuf_1 _05435_ (.A(_01781_),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _05436_ (.A(_01776_),
    .X(_01782_));
 sky130_fd_sc_hd__and2_1 _05437_ (.A(\wb_dat_o[28] ),
    .B(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__clkbuf_1 _05438_ (.A(_01783_),
    .X(net130));
 sky130_fd_sc_hd__and2_1 _05439_ (.A(\wb_dat_o[29] ),
    .B(_01782_),
    .X(_01784_));
 sky130_fd_sc_hd__clkbuf_1 _05440_ (.A(_01784_),
    .X(net131));
 sky130_fd_sc_hd__and2_1 _05441_ (.A(\wb_dat_o[30] ),
    .B(_01782_),
    .X(_01785_));
 sky130_fd_sc_hd__clkbuf_1 _05442_ (.A(_01785_),
    .X(net133));
 sky130_fd_sc_hd__and2_1 _05443_ (.A(\wb_dat_o[31] ),
    .B(_01782_),
    .X(_01786_));
 sky130_fd_sc_hd__clkbuf_1 _05444_ (.A(_01786_),
    .X(net134));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05445_ (.A(_01478_),
    .X(_01787_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05446_ (.A(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05447_ (.A(\u_async_wb.u_resp_if.rd_ptr[0] ),
    .X(_01789_));
 sky130_fd_sc_hd__clkbuf_1 _05448_ (.A(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _05449_ (.A0(\u_async_wb.u_resp_if.mem[0][32] ),
    .A1(\u_async_wb.u_resp_if.mem[1][32] ),
    .S(_01790_),
    .X(_01791_));
 sky130_fd_sc_hd__and2_1 _05450_ (.A(_01788_),
    .B(_01791_),
    .X(_01792_));
 sky130_fd_sc_hd__clkbuf_4 _05451_ (.A(_01792_),
    .X(wb_err_o1));
 sky130_fd_sc_hd__clkinv_2 _05452_ (.A(\u_reg.u_wbclk.clk_div_2 ),
    .Y(_00025_));
 sky130_fd_sc_hd__clkinv_2 _05453_ (.A(\u_reg.cpu_ref_clk_div_2 ),
    .Y(_00022_));
 sky130_fd_sc_hd__clkbuf_1 _05454_ (.A(net304),
    .X(_01793_));
 sky130_fd_sc_hd__buf_2 _05455_ (.A(_01793_),
    .X(_01794_));
 sky130_fd_sc_hd__and2_1 _05456_ (.A(_01794_),
    .B(\u_reg.cfg_glb_ctrl[0] ),
    .X(_01795_));
 sky130_fd_sc_hd__clkbuf_1 _05457_ (.A(_01795_),
    .X(\u_reg.u_buf_wb_rst.A ));
 sky130_fd_sc_hd__clkbuf_1 _05458_ (.A(net291),
    .X(_01796_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05459_ (.A(_01796_),
    .X(_01797_));
 sky130_fd_sc_hd__clkbuf_1 _05460_ (.A(_01797_),
    .X(_01798_));
 sky130_fd_sc_hd__buf_2 _05461_ (.A(_01798_),
    .X(_01799_));
 sky130_fd_sc_hd__and2_1 _05462_ (.A(_01799_),
    .B(\u_reg.cfg_glb_ctrl[1] ),
    .X(_01800_));
 sky130_fd_sc_hd__clkbuf_1 _05463_ (.A(_01800_),
    .X(\u_reg.u_buf_pll_rst.A ));
 sky130_fd_sc_hd__and2_1 _05464_ (.A(\u_uart2wb.u_aut_det.state[1] ),
    .B(_01178_),
    .X(_01801_));
 sky130_fd_sc_hd__clkbuf_1 _05465_ (.A(_01801_),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_1 _05466_ (.A(\u_reg.u_wbclk.clk_div_4 ),
    .B(\u_reg.u_wbclk.clk_div_2 ),
    .Y(_01802_));
 sky130_fd_sc_hd__or2_1 _05467_ (.A(\u_reg.u_wbclk.clk_div_4 ),
    .B(\u_reg.u_wbclk.clk_div_2 ),
    .X(_01803_));
 sky130_fd_sc_hd__and2_1 _05468_ (.A(_01802_),
    .B(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__clkbuf_1 _05469_ (.A(_01804_),
    .X(_00026_));
 sky130_fd_sc_hd__xnor2_1 _05470_ (.A(\u_reg.u_wbclk.clk_div_8 ),
    .B(_01802_),
    .Y(_00027_));
 sky130_fd_sc_hd__xor2_1 _05471_ (.A(_01105_),
    .B(_01134_),
    .X(_00033_));
 sky130_fd_sc_hd__a21oi_1 _05472_ (.A1(_01105_),
    .A2(_01134_),
    .B1(\u_uart2wb.u_core.u_txfsm.divcnt[2] ),
    .Y(_01805_));
 sky130_fd_sc_hd__and3_1 _05473_ (.A(_01105_),
    .B(_01134_),
    .C(\u_uart2wb.u_core.u_txfsm.divcnt[2] ),
    .X(_01806_));
 sky130_fd_sc_hd__nor2_1 _05474_ (.A(_01805_),
    .B(_01806_),
    .Y(_00034_));
 sky130_fd_sc_hd__xor2_1 _05475_ (.A(\u_uart2wb.u_core.u_txfsm.divcnt[3] ),
    .B(_01806_),
    .X(_00035_));
 sky130_fd_sc_hd__nand2_1 _05476_ (.A(\u_reg.cpu_ref_clk_div_4 ),
    .B(\u_reg.cpu_ref_clk_div_2 ),
    .Y(_01807_));
 sky130_fd_sc_hd__or2_1 _05477_ (.A(\u_reg.cpu_ref_clk_div_4 ),
    .B(\u_reg.cpu_ref_clk_div_2 ),
    .X(_01808_));
 sky130_fd_sc_hd__and2_1 _05478_ (.A(_01807_),
    .B(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__clkbuf_1 _05479_ (.A(_01809_),
    .X(_00023_));
 sky130_fd_sc_hd__xnor2_1 _05480_ (.A(\u_reg.cpu_ref_clk_div_8 ),
    .B(_01807_),
    .Y(_00024_));
 sky130_fd_sc_hd__clkbuf_1 _05481_ (.A(\u_uart2wb.u_core.u_rxfsm.offset[1] ),
    .X(_01810_));
 sky130_fd_sc_hd__xor2_1 _05482_ (.A(_01108_),
    .B(_01810_),
    .X(_00029_));
 sky130_fd_sc_hd__and3_1 _05483_ (.A(\u_uart2wb.u_core.u_rxfsm.offset[0] ),
    .B(_01810_),
    .C(\u_uart2wb.u_core.u_rxfsm.offset[2] ),
    .X(_01811_));
 sky130_fd_sc_hd__a21oi_1 _05484_ (.A1(_01108_),
    .A2(_01810_),
    .B1(\u_uart2wb.u_core.u_rxfsm.offset[2] ),
    .Y(_01812_));
 sky130_fd_sc_hd__nor2_1 _05485_ (.A(_01811_),
    .B(_01812_),
    .Y(_00030_));
 sky130_fd_sc_hd__inv_2 _05486_ (.A(\u_uart2wb.u_core.u_rxfsm.offset[3] ),
    .Y(_01813_));
 sky130_fd_sc_hd__xnor2_1 _05487_ (.A(_01813_),
    .B(_01811_),
    .Y(_00031_));
 sky130_fd_sc_hd__and2_1 _05488_ (.A(_01511_),
    .B(_01742_),
    .X(_01814_));
 sky130_fd_sc_hd__clkbuf_1 _05489_ (.A(_01814_),
    .X(net109));
 sky130_fd_sc_hd__and2_1 _05490_ (.A(wb_err_o),
    .B(_01742_),
    .X(_01815_));
 sky130_fd_sc_hd__clkbuf_1 _05491_ (.A(_01815_),
    .X(net142));
 sky130_fd_sc_hd__or3_1 _05492_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[0] ),
    .B(\u_uart2wb.u_core.u_clk_ctl.low_count[1] ),
    .C(\u_uart2wb.u_core.u_clk_ctl.low_count[2] ),
    .X(_01816_));
 sky130_fd_sc_hd__or2_1 _05493_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[3] ),
    .B(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__or2_1 _05494_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[4] ),
    .B(_01817_),
    .X(_01818_));
 sky130_fd_sc_hd__or2_1 _05495_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[5] ),
    .B(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__or2_1 _05496_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[6] ),
    .B(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__or3_1 _05497_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[7] ),
    .B(\u_uart2wb.u_core.u_clk_ctl.low_count[8] ),
    .C(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__or2_1 _05498_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[9] ),
    .B(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__or3_1 _05499_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[11] ),
    .B(\u_uart2wb.u_core.u_clk_ctl.low_count[10] ),
    .C(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05500_ (.A(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05501_ (.A(_01824_),
    .X(_01825_));
 sky130_fd_sc_hd__or4_1 _05502_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[0] ),
    .B(\u_uart2wb.u_core.u_clk_ctl.high_count[1] ),
    .C(\u_uart2wb.u_core.u_clk_ctl.high_count[3] ),
    .D(\u_uart2wb.u_core.u_clk_ctl.high_count[2] ),
    .X(_01826_));
 sky130_fd_sc_hd__or3_1 _05503_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[5] ),
    .B(\u_uart2wb.u_core.u_clk_ctl.high_count[4] ),
    .C(_01826_),
    .X(_01827_));
 sky130_fd_sc_hd__or2_1 _05504_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[6] ),
    .B(_01827_),
    .X(_01828_));
 sky130_fd_sc_hd__or3_1 _05505_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[7] ),
    .B(\u_uart2wb.u_core.u_clk_ctl.high_count[8] ),
    .C(_01828_),
    .X(_01829_));
 sky130_fd_sc_hd__or2_1 _05506_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[9] ),
    .B(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__or2_1 _05507_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[10] ),
    .B(_01830_),
    .X(_01831_));
 sky130_fd_sc_hd__nor2_1 _05508_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[11] ),
    .B(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__clkbuf_1 _05509_ (.A(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05510_ (.A(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__o21ai_1 _05511_ (.A1(\u_uart2wb.u_core.line_clk_16x ),
    .A2(_01825_),
    .B1(_01834_),
    .Y(_00021_));
 sky130_fd_sc_hd__and3_2 _05512_ (.A(_01472_),
    .B(_01729_),
    .C(wb_ack_o),
    .X(_01835_));
 sky130_fd_sc_hd__clkbuf_1 _05513_ (.A(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__clkbuf_2 _05514_ (.A(_01836_),
    .X(_01837_));
 sky130_fd_sc_hd__o32a_1 _05515_ (.A1(_01458_),
    .A2(_01111_),
    .A3(_01450_),
    .B1(_01460_),
    .B2(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__nor3b_1 _05516_ (.A(_01459_),
    .B(_01838_),
    .C_N(\u_spi2wb.reg_rd ),
    .Y(_01839_));
 sky130_fd_sc_hd__a31o_1 _05517_ (.A1(_01458_),
    .A2(_01121_),
    .A3(_01132_),
    .B1(_01839_),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _05518_ (.A0(\u_async_wb.u_resp_if.mem[0][0] ),
    .A1(\u_async_wb.u_resp_if.mem[1][0] ),
    .S(_01790_),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_2 _05519_ (.A0(\u_reg.reg_rdata[0] ),
    .A1(_01840_),
    .S(_01788_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _05520_ (.A0(\wb_dat_o[0] ),
    .A1(_01841_),
    .S(wb_ack_o1),
    .X(_01842_));
 sky130_fd_sc_hd__clkbuf_1 _05521_ (.A(_01842_),
    .X(_00039_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05522_ (.A(\u_async_wb.u_resp_if.rd_ptr[0] ),
    .X(_01843_));
 sky130_fd_sc_hd__clkbuf_1 _05523_ (.A(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__clkbuf_2 _05524_ (.A(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _05525_ (.A0(\u_async_wb.u_resp_if.mem[0][1] ),
    .A1(\u_async_wb.u_resp_if.mem[1][1] ),
    .S(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_2 _05526_ (.A0(\u_reg.reg_rdata[1] ),
    .A1(_01846_),
    .S(_01788_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _05527_ (.A0(\wb_dat_o[1] ),
    .A1(_01847_),
    .S(wb_ack_o1),
    .X(_01848_));
 sky130_fd_sc_hd__clkbuf_1 _05528_ (.A(_01848_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _05529_ (.A0(\u_async_wb.u_resp_if.mem[0][2] ),
    .A1(\u_async_wb.u_resp_if.mem[1][2] ),
    .S(_01845_),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _05530_ (.A0(\u_reg.reg_rdata[2] ),
    .A1(_01849_),
    .S(_01788_),
    .X(_01850_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05531_ (.A(_01510_),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _05532_ (.A0(\wb_dat_o[2] ),
    .A1(_01850_),
    .S(_01851_),
    .X(_01852_));
 sky130_fd_sc_hd__clkbuf_1 _05533_ (.A(_01852_),
    .X(_00041_));
 sky130_fd_sc_hd__mux2_1 _05534_ (.A0(\u_async_wb.u_resp_if.mem[0][3] ),
    .A1(\u_async_wb.u_resp_if.mem[1][3] ),
    .S(_01845_),
    .X(_01853_));
 sky130_fd_sc_hd__clkbuf_2 _05535_ (.A(_01787_),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _05536_ (.A0(\u_reg.reg_rdata[3] ),
    .A1(_01853_),
    .S(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _05537_ (.A0(\wb_dat_o[3] ),
    .A1(_01855_),
    .S(_01851_),
    .X(_01856_));
 sky130_fd_sc_hd__clkbuf_1 _05538_ (.A(_01856_),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _05539_ (.A0(\u_async_wb.u_resp_if.mem[0][4] ),
    .A1(\u_async_wb.u_resp_if.mem[1][4] ),
    .S(_01845_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _05540_ (.A0(\u_reg.reg_rdata[4] ),
    .A1(_01857_),
    .S(_01854_),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _05541_ (.A0(\wb_dat_o[4] ),
    .A1(_01858_),
    .S(_01851_),
    .X(_01859_));
 sky130_fd_sc_hd__clkbuf_1 _05542_ (.A(_01859_),
    .X(_00043_));
 sky130_fd_sc_hd__clkbuf_2 _05543_ (.A(_01844_),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _05544_ (.A0(\u_async_wb.u_resp_if.mem[0][5] ),
    .A1(\u_async_wb.u_resp_if.mem[1][5] ),
    .S(_01860_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _05545_ (.A0(\u_reg.reg_rdata[5] ),
    .A1(_01861_),
    .S(_01854_),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _05546_ (.A0(\wb_dat_o[5] ),
    .A1(_01862_),
    .S(_01851_),
    .X(_01863_));
 sky130_fd_sc_hd__clkbuf_1 _05547_ (.A(_01863_),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _05548_ (.A0(\u_async_wb.u_resp_if.mem[0][6] ),
    .A1(\u_async_wb.u_resp_if.mem[1][6] ),
    .S(_01860_),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _05549_ (.A0(\u_reg.reg_rdata[6] ),
    .A1(_01864_),
    .S(_01854_),
    .X(_01865_));
 sky130_fd_sc_hd__clkbuf_1 _05550_ (.A(_01509_),
    .X(_01866_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05551_ (.A(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _05552_ (.A0(\wb_dat_o[6] ),
    .A1(_01865_),
    .S(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__clkbuf_1 _05553_ (.A(_01868_),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _05554_ (.A0(\u_async_wb.u_resp_if.mem[0][7] ),
    .A1(\u_async_wb.u_resp_if.mem[1][7] ),
    .S(_01860_),
    .X(_01869_));
 sky130_fd_sc_hd__clkbuf_2 _05555_ (.A(_01787_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_2 _05556_ (.A0(\u_reg.reg_rdata[7] ),
    .A1(_01869_),
    .S(_01870_),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _05557_ (.A0(\wb_dat_o[7] ),
    .A1(_01871_),
    .S(_01867_),
    .X(_01872_));
 sky130_fd_sc_hd__clkbuf_1 _05558_ (.A(_01872_),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _05559_ (.A0(\u_async_wb.u_resp_if.mem[0][8] ),
    .A1(\u_async_wb.u_resp_if.mem[1][8] ),
    .S(_01860_),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _05560_ (.A0(\u_reg.reg_rdata[8] ),
    .A1(_01873_),
    .S(_01870_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _05561_ (.A0(\wb_dat_o[8] ),
    .A1(_01874_),
    .S(_01867_),
    .X(_01875_));
 sky130_fd_sc_hd__clkbuf_1 _05562_ (.A(_01875_),
    .X(_00047_));
 sky130_fd_sc_hd__clkbuf_2 _05563_ (.A(_01844_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _05564_ (.A0(\u_async_wb.u_resp_if.mem[0][9] ),
    .A1(\u_async_wb.u_resp_if.mem[1][9] ),
    .S(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_2 _05565_ (.A0(\u_reg.reg_rdata[9] ),
    .A1(_01877_),
    .S(_01870_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _05566_ (.A0(\wb_dat_o[9] ),
    .A1(_01878_),
    .S(_01867_),
    .X(_01879_));
 sky130_fd_sc_hd__clkbuf_1 _05567_ (.A(_01879_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _05568_ (.A0(\u_async_wb.u_resp_if.mem[0][10] ),
    .A1(\u_async_wb.u_resp_if.mem[1][10] ),
    .S(_01876_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_2 _05569_ (.A0(\u_reg.reg_rdata[10] ),
    .A1(_01880_),
    .S(_01870_),
    .X(_01881_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05570_ (.A(_01866_),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _05571_ (.A0(\wb_dat_o[10] ),
    .A1(_01881_),
    .S(_01882_),
    .X(_01883_));
 sky130_fd_sc_hd__clkbuf_1 _05572_ (.A(_01883_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _05573_ (.A0(\u_async_wb.u_resp_if.mem[0][11] ),
    .A1(\u_async_wb.u_resp_if.mem[1][11] ),
    .S(_01876_),
    .X(_01884_));
 sky130_fd_sc_hd__clkbuf_1 _05574_ (.A(_01479_),
    .X(_01885_));
 sky130_fd_sc_hd__clkbuf_2 _05575_ (.A(_01885_),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _05576_ (.A0(\u_reg.reg_rdata[11] ),
    .A1(_01884_),
    .S(_01886_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _05577_ (.A0(\wb_dat_o[11] ),
    .A1(_01887_),
    .S(_01882_),
    .X(_01888_));
 sky130_fd_sc_hd__clkbuf_1 _05578_ (.A(_01888_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _05579_ (.A0(\u_async_wb.u_resp_if.mem[0][12] ),
    .A1(\u_async_wb.u_resp_if.mem[1][12] ),
    .S(_01876_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _05580_ (.A0(\u_reg.reg_rdata[12] ),
    .A1(_01889_),
    .S(_01886_),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _05581_ (.A0(\wb_dat_o[12] ),
    .A1(_01890_),
    .S(_01882_),
    .X(_01891_));
 sky130_fd_sc_hd__clkbuf_1 _05582_ (.A(_01891_),
    .X(_00051_));
 sky130_fd_sc_hd__clkbuf_2 _05583_ (.A(_01844_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _05584_ (.A0(\u_async_wb.u_resp_if.mem[0][13] ),
    .A1(\u_async_wb.u_resp_if.mem[1][13] ),
    .S(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__mux2_1 _05585_ (.A0(\u_reg.reg_rdata[13] ),
    .A1(_01893_),
    .S(_01886_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _05586_ (.A0(\wb_dat_o[13] ),
    .A1(_01894_),
    .S(_01882_),
    .X(_01895_));
 sky130_fd_sc_hd__clkbuf_1 _05587_ (.A(_01895_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _05588_ (.A0(\u_async_wb.u_resp_if.mem[0][14] ),
    .A1(\u_async_wb.u_resp_if.mem[1][14] ),
    .S(_01892_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_2 _05589_ (.A0(\u_reg.reg_rdata[14] ),
    .A1(_01896_),
    .S(_01886_),
    .X(_01897_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05590_ (.A(_01866_),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _05591_ (.A0(\wb_dat_o[14] ),
    .A1(_01897_),
    .S(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__clkbuf_1 _05592_ (.A(_01899_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _05593_ (.A0(\u_async_wb.u_resp_if.mem[0][15] ),
    .A1(\u_async_wb.u_resp_if.mem[1][15] ),
    .S(_01892_),
    .X(_01900_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05594_ (.A(_01885_),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_1 _05595_ (.A0(\u_reg.reg_rdata[15] ),
    .A1(_01900_),
    .S(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _05596_ (.A0(\wb_dat_o[15] ),
    .A1(_01902_),
    .S(_01898_),
    .X(_01903_));
 sky130_fd_sc_hd__clkbuf_1 _05597_ (.A(_01903_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _05598_ (.A0(\u_async_wb.u_resp_if.mem[0][16] ),
    .A1(\u_async_wb.u_resp_if.mem[1][16] ),
    .S(_01892_),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_1 _05599_ (.A0(\u_reg.reg_rdata[16] ),
    .A1(_01904_),
    .S(_01901_),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _05600_ (.A0(\wb_dat_o[16] ),
    .A1(_01905_),
    .S(_01898_),
    .X(_01906_));
 sky130_fd_sc_hd__clkbuf_1 _05601_ (.A(_01906_),
    .X(_00055_));
 sky130_fd_sc_hd__clkbuf_2 _05602_ (.A(_01843_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _05603_ (.A0(\u_async_wb.u_resp_if.mem[0][17] ),
    .A1(\u_async_wb.u_resp_if.mem[1][17] ),
    .S(_01907_),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _05604_ (.A0(\u_reg.reg_rdata[17] ),
    .A1(_01908_),
    .S(_01901_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _05605_ (.A0(\wb_dat_o[17] ),
    .A1(_01909_),
    .S(_01898_),
    .X(_01910_));
 sky130_fd_sc_hd__clkbuf_1 _05606_ (.A(_01910_),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _05607_ (.A0(\u_async_wb.u_resp_if.mem[0][18] ),
    .A1(\u_async_wb.u_resp_if.mem[1][18] ),
    .S(_01907_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _05608_ (.A0(\u_reg.reg_rdata[18] ),
    .A1(_01911_),
    .S(_01901_),
    .X(_01912_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05609_ (.A(_01866_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _05610_ (.A0(\wb_dat_o[18] ),
    .A1(_01912_),
    .S(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__clkbuf_1 _05611_ (.A(_01914_),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _05612_ (.A0(\u_async_wb.u_resp_if.mem[0][19] ),
    .A1(\u_async_wb.u_resp_if.mem[1][19] ),
    .S(_01907_),
    .X(_01915_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05613_ (.A(_01885_),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_1 _05614_ (.A0(\u_reg.reg_rdata[19] ),
    .A1(_01915_),
    .S(_01916_),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _05615_ (.A0(\wb_dat_o[19] ),
    .A1(_01917_),
    .S(_01913_),
    .X(_01918_));
 sky130_fd_sc_hd__clkbuf_1 _05616_ (.A(_01918_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _05617_ (.A0(\u_async_wb.u_resp_if.mem[0][20] ),
    .A1(\u_async_wb.u_resp_if.mem[1][20] ),
    .S(_01907_),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _05618_ (.A0(\u_reg.reg_rdata[20] ),
    .A1(_01919_),
    .S(_01916_),
    .X(_01920_));
 sky130_fd_sc_hd__mux2_1 _05619_ (.A0(\wb_dat_o[20] ),
    .A1(_01920_),
    .S(_01913_),
    .X(_01921_));
 sky130_fd_sc_hd__clkbuf_1 _05620_ (.A(_01921_),
    .X(_00059_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05621_ (.A(_01843_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _05622_ (.A0(\u_async_wb.u_resp_if.mem[0][21] ),
    .A1(\u_async_wb.u_resp_if.mem[1][21] ),
    .S(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__mux2_1 _05623_ (.A0(\u_reg.reg_rdata[21] ),
    .A1(_01923_),
    .S(_01916_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _05624_ (.A0(\wb_dat_o[21] ),
    .A1(_01924_),
    .S(_01913_),
    .X(_01925_));
 sky130_fd_sc_hd__clkbuf_1 _05625_ (.A(_01925_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _05626_ (.A0(\u_async_wb.u_resp_if.mem[0][22] ),
    .A1(\u_async_wb.u_resp_if.mem[1][22] ),
    .S(_01922_),
    .X(_01926_));
 sky130_fd_sc_hd__mux2_1 _05627_ (.A0(\u_reg.reg_rdata[22] ),
    .A1(_01926_),
    .S(_01916_),
    .X(_01927_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05628_ (.A(_01509_),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _05629_ (.A0(\wb_dat_o[22] ),
    .A1(_01927_),
    .S(_01928_),
    .X(_01929_));
 sky130_fd_sc_hd__clkbuf_1 _05630_ (.A(_01929_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _05631_ (.A0(\u_async_wb.u_resp_if.mem[0][23] ),
    .A1(\u_async_wb.u_resp_if.mem[1][23] ),
    .S(_01922_),
    .X(_01930_));
 sky130_fd_sc_hd__clkbuf_2 _05632_ (.A(_01885_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _05633_ (.A0(\u_reg.reg_rdata[23] ),
    .A1(_01930_),
    .S(_01931_),
    .X(_01932_));
 sky130_fd_sc_hd__mux2_1 _05634_ (.A0(\wb_dat_o[23] ),
    .A1(_01932_),
    .S(_01928_),
    .X(_01933_));
 sky130_fd_sc_hd__clkbuf_1 _05635_ (.A(_01933_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _05636_ (.A0(\u_async_wb.u_resp_if.mem[0][24] ),
    .A1(\u_async_wb.u_resp_if.mem[1][24] ),
    .S(_01922_),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_1 _05637_ (.A0(\u_reg.reg_rdata[24] ),
    .A1(_01934_),
    .S(_01931_),
    .X(_01935_));
 sky130_fd_sc_hd__mux2_1 _05638_ (.A0(\wb_dat_o[24] ),
    .A1(_01935_),
    .S(_01928_),
    .X(_01936_));
 sky130_fd_sc_hd__clkbuf_1 _05639_ (.A(_01936_),
    .X(_00063_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05640_ (.A(_01843_),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _05641_ (.A0(\u_async_wb.u_resp_if.mem[0][25] ),
    .A1(\u_async_wb.u_resp_if.mem[1][25] ),
    .S(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_1 _05642_ (.A0(\u_reg.reg_rdata[25] ),
    .A1(_01938_),
    .S(_01931_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _05643_ (.A0(\wb_dat_o[25] ),
    .A1(_01939_),
    .S(_01928_),
    .X(_01940_));
 sky130_fd_sc_hd__clkbuf_1 _05644_ (.A(_01940_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _05645_ (.A0(\u_async_wb.u_resp_if.mem[0][26] ),
    .A1(\u_async_wb.u_resp_if.mem[1][26] ),
    .S(_01937_),
    .X(_01941_));
 sky130_fd_sc_hd__mux2_1 _05646_ (.A0(\u_reg.reg_rdata[26] ),
    .A1(_01941_),
    .S(_01931_),
    .X(_01942_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05647_ (.A(_01509_),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_1 _05648_ (.A0(\wb_dat_o[26] ),
    .A1(_01942_),
    .S(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__clkbuf_1 _05649_ (.A(_01944_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _05650_ (.A0(\u_async_wb.u_resp_if.mem[0][27] ),
    .A1(\u_async_wb.u_resp_if.mem[1][27] ),
    .S(_01937_),
    .X(_01945_));
 sky130_fd_sc_hd__clkbuf_2 _05651_ (.A(_01479_),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _05652_ (.A0(\u_reg.reg_rdata[27] ),
    .A1(_01945_),
    .S(_01946_),
    .X(_01947_));
 sky130_fd_sc_hd__mux2_1 _05653_ (.A0(\wb_dat_o[27] ),
    .A1(_01947_),
    .S(_01943_),
    .X(_01948_));
 sky130_fd_sc_hd__clkbuf_1 _05654_ (.A(_01948_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _05655_ (.A0(\u_async_wb.u_resp_if.mem[0][28] ),
    .A1(\u_async_wb.u_resp_if.mem[1][28] ),
    .S(_01937_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _05656_ (.A0(\u_reg.reg_rdata[28] ),
    .A1(_01949_),
    .S(_01946_),
    .X(_01950_));
 sky130_fd_sc_hd__mux2_1 _05657_ (.A0(\wb_dat_o[28] ),
    .A1(_01950_),
    .S(_01943_),
    .X(_01951_));
 sky130_fd_sc_hd__clkbuf_1 _05658_ (.A(_01951_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _05659_ (.A0(\u_async_wb.u_resp_if.mem[0][29] ),
    .A1(\u_async_wb.u_resp_if.mem[1][29] ),
    .S(_01789_),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_1 _05660_ (.A0(\u_reg.reg_rdata[29] ),
    .A1(_01952_),
    .S(_01946_),
    .X(_01953_));
 sky130_fd_sc_hd__mux2_1 _05661_ (.A0(\wb_dat_o[29] ),
    .A1(_01953_),
    .S(_01943_),
    .X(_01954_));
 sky130_fd_sc_hd__clkbuf_1 _05662_ (.A(_01954_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _05663_ (.A0(\u_async_wb.u_resp_if.mem[0][30] ),
    .A1(\u_async_wb.u_resp_if.mem[1][30] ),
    .S(_01789_),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _05664_ (.A0(\u_reg.reg_rdata[30] ),
    .A1(_01955_),
    .S(_01946_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _05665_ (.A0(\wb_dat_o[30] ),
    .A1(_01956_),
    .S(_01510_),
    .X(_01957_));
 sky130_fd_sc_hd__clkbuf_1 _05666_ (.A(_01957_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _05667_ (.A0(\u_async_wb.u_resp_if.mem[0][31] ),
    .A1(\u_async_wb.u_resp_if.mem[1][31] ),
    .S(_01789_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _05668_ (.A0(\u_reg.reg_rdata[31] ),
    .A1(_01958_),
    .S(_01787_),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_1 _05669_ (.A0(\wb_dat_o[31] ),
    .A1(_01959_),
    .S(_01510_),
    .X(_01960_));
 sky130_fd_sc_hd__clkbuf_1 _05670_ (.A(_01960_),
    .X(_00070_));
 sky130_fd_sc_hd__inv_2 _05671_ (.A(\u_reset_fsm.state[1] ),
    .Y(_01961_));
 sky130_fd_sc_hd__clkbuf_1 _05672_ (.A(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__or2_1 _05673_ (.A(_01962_),
    .B(\u_reset_fsm.state[0] ),
    .X(_01963_));
 sky130_fd_sc_hd__nor2_1 _05674_ (.A(_01961_),
    .B(\u_reset_fsm.state[0] ),
    .Y(_01964_));
 sky130_fd_sc_hd__and3_1 _05675_ (.A(\u_reset_fsm.state[2] ),
    .B(\u_reset_fsm.boot_req_ss ),
    .C(_01964_),
    .X(_01965_));
 sky130_fd_sc_hd__nor2_1 _05676_ (.A(_01963_),
    .B(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__clkbuf_1 _05677_ (.A(\u_reset_fsm.state[2] ),
    .X(_01967_));
 sky130_fd_sc_hd__clkbuf_1 _05678_ (.A(\u_reset_fsm.clk_cnt[11] ),
    .X(_01968_));
 sky130_fd_sc_hd__or3_1 _05679_ (.A(\u_reset_fsm.clk_cnt[13] ),
    .B(\u_reset_fsm.clk_cnt[15] ),
    .C(\u_reset_fsm.clk_cnt[14] ),
    .X(_01969_));
 sky130_fd_sc_hd__or4b_1 _05680_ (.A(\u_reset_fsm.clk_cnt[9] ),
    .B(_01968_),
    .C(_01969_),
    .D_N(\u_reset_fsm.clk_cnt[2] ),
    .X(_01970_));
 sky130_fd_sc_hd__or3_1 _05681_ (.A(\u_reset_fsm.clk_cnt[4] ),
    .B(\u_reset_fsm.clk_cnt[8] ),
    .C(\u_reset_fsm.clk_cnt[10] ),
    .X(_01971_));
 sky130_fd_sc_hd__clkbuf_1 _05682_ (.A(\u_reset_fsm.clk_cnt[1] ),
    .X(_01972_));
 sky130_fd_sc_hd__clkbuf_1 _05683_ (.A(\u_reset_fsm.clk_cnt[0] ),
    .X(_01973_));
 sky130_fd_sc_hd__or2_1 _05684_ (.A(_01972_),
    .B(_01973_),
    .X(_01974_));
 sky130_fd_sc_hd__clkbuf_1 _05685_ (.A(\u_reset_fsm.clk_cnt[5] ),
    .X(_01975_));
 sky130_fd_sc_hd__or4bb_1 _05686_ (.A(\u_reset_fsm.clk_cnt[7] ),
    .B(\u_reset_fsm.clk_cnt[12] ),
    .C_N(\u_reset_fsm.clk_cnt[6] ),
    .D_N(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__and4b_1 _05687_ (.A_N(\u_reset_fsm.clk_cnt[2] ),
    .B(\u_reset_fsm.clk_cnt[9] ),
    .C(\u_reset_fsm.clk_cnt[13] ),
    .D(\u_reset_fsm.clk_cnt[15] ),
    .X(_01977_));
 sky130_fd_sc_hd__a31o_1 _05688_ (.A1(\u_reset_fsm.clk_cnt[11] ),
    .A2(\u_reset_fsm.clk_cnt[14] ),
    .A3(_01977_),
    .B1(net65),
    .X(_01978_));
 sky130_fd_sc_hd__or4b_1 _05689_ (.A(\u_reset_fsm.clk_cnt[3] ),
    .B(_01974_),
    .C(_01976_),
    .D_N(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__a211oi_2 _05690_ (.A1(net65),
    .A2(_01970_),
    .B1(_01971_),
    .C1(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__a21oi_1 _05691_ (.A1(_01961_),
    .A2(\u_reset_fsm.state[2] ),
    .B1(\u_reset_fsm.state[0] ),
    .Y(_01981_));
 sky130_fd_sc_hd__o21ai_1 _05692_ (.A1(_01967_),
    .A2(_01980_),
    .B1(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__inv_2 _05693_ (.A(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__nor2_1 _05694_ (.A(_01966_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__clkbuf_1 _05695_ (.A(_01966_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _05696_ (.A0(_01984_),
    .A1(_01985_),
    .S(_01973_),
    .X(_01986_));
 sky130_fd_sc_hd__clkbuf_1 _05697_ (.A(_01986_),
    .X(_00071_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05698_ (.A(_01963_),
    .X(_01987_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05699_ (.A(_01987_),
    .X(_01988_));
 sky130_fd_sc_hd__nand2_1 _05700_ (.A(_01972_),
    .B(_01973_),
    .Y(_01989_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05701_ (.A(_01985_),
    .X(_01990_));
 sky130_fd_sc_hd__a32o_1 _05702_ (.A1(_01988_),
    .A2(_01974_),
    .A3(_01989_),
    .B1(_01990_),
    .B2(_01972_),
    .X(_00072_));
 sky130_fd_sc_hd__o211a_1 _05703_ (.A1(_01987_),
    .A2(_01965_),
    .B1(_01972_),
    .C1(_01973_),
    .X(_01991_));
 sky130_fd_sc_hd__and3_1 _05704_ (.A(\u_reset_fsm.clk_cnt[1] ),
    .B(\u_reset_fsm.clk_cnt[0] ),
    .C(\u_reset_fsm.clk_cnt[2] ),
    .X(_01992_));
 sky130_fd_sc_hd__clkbuf_1 _05705_ (.A(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__nor2_1 _05706_ (.A(_01983_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__clkbuf_1 _05707_ (.A(_01966_),
    .X(_01995_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05708_ (.A(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__o22a_1 _05709_ (.A1(\u_reset_fsm.clk_cnt[2] ),
    .A2(_01991_),
    .B1(_01994_),
    .B2(_01996_),
    .X(_00073_));
 sky130_fd_sc_hd__clkbuf_1 _05710_ (.A(\u_reset_fsm.clk_cnt[3] ),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_1 _05711_ (.A(_01997_),
    .B(_01993_),
    .Y(_01998_));
 sky130_fd_sc_hd__or2_1 _05712_ (.A(_01997_),
    .B(_01993_),
    .X(_01999_));
 sky130_fd_sc_hd__a32o_1 _05713_ (.A1(_01988_),
    .A2(_01998_),
    .A3(_01999_),
    .B1(_01990_),
    .B2(_01997_),
    .X(_00074_));
 sky130_fd_sc_hd__nor2_1 _05714_ (.A(_01995_),
    .B(_01998_),
    .Y(_02000_));
 sky130_fd_sc_hd__clkbuf_1 _05715_ (.A(\u_reset_fsm.clk_cnt[9] ),
    .X(_02001_));
 sky130_fd_sc_hd__or4_1 _05716_ (.A(_01975_),
    .B(_02001_),
    .C(_01968_),
    .D(_01971_),
    .X(_02002_));
 sky130_fd_sc_hd__clkbuf_1 _05717_ (.A(\u_reset_fsm.clk_cnt[7] ),
    .X(_02003_));
 sky130_fd_sc_hd__clkbuf_1 _05718_ (.A(\u_reset_fsm.clk_cnt[6] ),
    .X(_02004_));
 sky130_fd_sc_hd__clkbuf_1 _05719_ (.A(\u_reset_fsm.clk_cnt[12] ),
    .X(_02005_));
 sky130_fd_sc_hd__or4_1 _05720_ (.A(_02003_),
    .B(_02004_),
    .C(_02005_),
    .D(_01969_),
    .X(_02006_));
 sky130_fd_sc_hd__nor3_1 _05721_ (.A(_01998_),
    .B(_02002_),
    .C(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05722_ (.A(_02007_),
    .X(_02008_));
 sky130_fd_sc_hd__inv_2 _05723_ (.A(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__and3_1 _05724_ (.A(_01997_),
    .B(\u_reset_fsm.clk_cnt[4] ),
    .C(_01993_),
    .X(_02010_));
 sky130_fd_sc_hd__inv_2 _05725_ (.A(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2_1 _05726_ (.A(\u_reset_fsm.state[2] ),
    .B(_01964_),
    .Y(_02012_));
 sky130_fd_sc_hd__o211a_1 _05727_ (.A1(_01981_),
    .A2(_02009_),
    .B1(_02011_),
    .C1(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__o22a_1 _05728_ (.A1(\u_reset_fsm.clk_cnt[4] ),
    .A2(_02000_),
    .B1(_02013_),
    .B2(_01996_),
    .X(_00075_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05729_ (.A(_01984_),
    .X(_02014_));
 sky130_fd_sc_hd__or2_1 _05730_ (.A(_01975_),
    .B(_02010_),
    .X(_02015_));
 sky130_fd_sc_hd__and2_1 _05731_ (.A(\u_reset_fsm.clk_cnt[3] ),
    .B(_01992_),
    .X(_02016_));
 sky130_fd_sc_hd__and3_1 _05732_ (.A(\u_reset_fsm.clk_cnt[4] ),
    .B(\u_reset_fsm.clk_cnt[5] ),
    .C(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__inv_2 _05733_ (.A(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__a32o_1 _05734_ (.A1(_02014_),
    .A2(_02015_),
    .A3(_02018_),
    .B1(_01990_),
    .B2(_01975_),
    .X(_00076_));
 sky130_fd_sc_hd__or2_1 _05735_ (.A(_02004_),
    .B(_02017_),
    .X(_02019_));
 sky130_fd_sc_hd__and2_1 _05736_ (.A(_02004_),
    .B(_02017_),
    .X(_02020_));
 sky130_fd_sc_hd__inv_2 _05737_ (.A(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__a32o_1 _05738_ (.A1(_02014_),
    .A2(_02019_),
    .A3(_02021_),
    .B1(_01990_),
    .B2(_02004_),
    .X(_00077_));
 sky130_fd_sc_hd__and3_1 _05739_ (.A(_02003_),
    .B(\u_reset_fsm.clk_cnt[6] ),
    .C(_02017_),
    .X(_02022_));
 sky130_fd_sc_hd__clkbuf_1 _05740_ (.A(_02022_),
    .X(_02023_));
 sky130_fd_sc_hd__o21ai_1 _05741_ (.A1(_02003_),
    .A2(_02020_),
    .B1(_01987_),
    .Y(_02024_));
 sky130_fd_sc_hd__a2bb2o_1 _05742_ (.A1_N(_02023_),
    .A2_N(_02024_),
    .B1(_02003_),
    .B2(_01996_),
    .X(_00078_));
 sky130_fd_sc_hd__clkbuf_1 _05743_ (.A(\u_reset_fsm.clk_cnt[8] ),
    .X(_02025_));
 sky130_fd_sc_hd__nand2_1 _05744_ (.A(_02025_),
    .B(_02023_),
    .Y(_02026_));
 sky130_fd_sc_hd__or2_1 _05745_ (.A(_02025_),
    .B(_02023_),
    .X(_02027_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05746_ (.A(_01985_),
    .X(_02028_));
 sky130_fd_sc_hd__a32o_1 _05747_ (.A1(_01988_),
    .A2(_02026_),
    .A3(_02027_),
    .B1(_02028_),
    .B2(_02025_),
    .X(_00079_));
 sky130_fd_sc_hd__and3_1 _05748_ (.A(_02001_),
    .B(\u_reset_fsm.clk_cnt[8] ),
    .C(_02022_),
    .X(_02029_));
 sky130_fd_sc_hd__inv_2 _05749_ (.A(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__a21o_1 _05750_ (.A1(_02025_),
    .A2(_02023_),
    .B1(_02001_),
    .X(_02031_));
 sky130_fd_sc_hd__a32o_1 _05751_ (.A1(_02014_),
    .A2(_02030_),
    .A3(_02031_),
    .B1(_02028_),
    .B2(_02001_),
    .X(_00080_));
 sky130_fd_sc_hd__clkbuf_1 _05752_ (.A(\u_reset_fsm.clk_cnt[10] ),
    .X(_02032_));
 sky130_fd_sc_hd__and2_1 _05753_ (.A(_02032_),
    .B(_02029_),
    .X(_02033_));
 sky130_fd_sc_hd__o21ai_1 _05754_ (.A1(_02032_),
    .A2(_02029_),
    .B1(_01987_),
    .Y(_02034_));
 sky130_fd_sc_hd__a2bb2o_1 _05755_ (.A1_N(_02033_),
    .A2_N(_02034_),
    .B1(_02032_),
    .B2(_01996_),
    .X(_00081_));
 sky130_fd_sc_hd__clkbuf_1 _05756_ (.A(_01968_),
    .X(_02035_));
 sky130_fd_sc_hd__nand2_1 _05757_ (.A(_02035_),
    .B(_02033_),
    .Y(_02036_));
 sky130_fd_sc_hd__or2_1 _05758_ (.A(_02035_),
    .B(_02033_),
    .X(_02037_));
 sky130_fd_sc_hd__a32o_1 _05759_ (.A1(_01984_),
    .A2(_02036_),
    .A3(_02037_),
    .B1(_02028_),
    .B2(_02035_),
    .X(_00082_));
 sky130_fd_sc_hd__a31o_1 _05760_ (.A1(_02035_),
    .A2(_02032_),
    .A3(_02029_),
    .B1(_02005_),
    .X(_02038_));
 sky130_fd_sc_hd__and3_1 _05761_ (.A(_01968_),
    .B(_02005_),
    .C(_02033_),
    .X(_02039_));
 sky130_fd_sc_hd__inv_2 _05762_ (.A(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__a32o_1 _05763_ (.A1(_01988_),
    .A2(_02038_),
    .A3(_02040_),
    .B1(_02028_),
    .B2(_02005_),
    .X(_00083_));
 sky130_fd_sc_hd__clkbuf_1 _05764_ (.A(\u_reset_fsm.clk_cnt[13] ),
    .X(_02041_));
 sky130_fd_sc_hd__nand2_1 _05765_ (.A(_02041_),
    .B(_02039_),
    .Y(_02042_));
 sky130_fd_sc_hd__or2_1 _05766_ (.A(_02041_),
    .B(_02039_),
    .X(_02043_));
 sky130_fd_sc_hd__a32o_1 _05767_ (.A1(_01984_),
    .A2(_02042_),
    .A3(_02043_),
    .B1(_01995_),
    .B2(_02041_),
    .X(_00084_));
 sky130_fd_sc_hd__nor2_1 _05768_ (.A(_01995_),
    .B(_02042_),
    .Y(_02044_));
 sky130_fd_sc_hd__nand3_1 _05769_ (.A(_02041_),
    .B(\u_reset_fsm.clk_cnt[14] ),
    .C(_02039_),
    .Y(_02045_));
 sky130_fd_sc_hd__a21o_1 _05770_ (.A1(_01982_),
    .A2(_02045_),
    .B1(_01985_),
    .X(_02046_));
 sky130_fd_sc_hd__o21a_1 _05771_ (.A1(\u_reset_fsm.clk_cnt[14] ),
    .A2(_02044_),
    .B1(_02046_),
    .X(_00085_));
 sky130_fd_sc_hd__nor2_1 _05772_ (.A(\u_reset_fsm.clk_cnt[15] ),
    .B(_02045_),
    .Y(_02047_));
 sky130_fd_sc_hd__a22o_1 _05773_ (.A1(\u_reset_fsm.clk_cnt[15] ),
    .A2(_02046_),
    .B1(_02047_),
    .B2(_02014_),
    .X(_00086_));
 sky130_fd_sc_hd__and2_2 _05774_ (.A(\u_spi2wb.u_if.cmd_phase ),
    .B(_01130_),
    .X(_02048_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05775_ (.A(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _05776_ (.A0(\u_spi2wb.reg_be[0] ),
    .A1(net308),
    .S(_02049_),
    .X(_02050_));
 sky130_fd_sc_hd__clkbuf_1 _05777_ (.A(_02050_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _05778_ (.A0(\u_spi2wb.reg_be[1] ),
    .A1(\u_spi2wb.reg_be[0] ),
    .S(_02049_),
    .X(_02051_));
 sky130_fd_sc_hd__clkbuf_1 _05779_ (.A(_02051_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _05780_ (.A0(\u_spi2wb.reg_be[2] ),
    .A1(\u_spi2wb.reg_be[1] ),
    .S(_02049_),
    .X(_02052_));
 sky130_fd_sc_hd__clkbuf_1 _05781_ (.A(_02052_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _05782_ (.A0(\u_spi2wb.reg_be[3] ),
    .A1(\u_spi2wb.reg_be[2] ),
    .S(_02049_),
    .X(_02053_));
 sky130_fd_sc_hd__clkbuf_1 _05783_ (.A(_02053_),
    .X(_00090_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05784_ (.A(_02048_),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _05785_ (.A0(\u_spi2wb.u_if.cmd_reg[4] ),
    .A1(\u_spi2wb.reg_be[3] ),
    .S(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__clkbuf_1 _05786_ (.A(_02055_),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _05787_ (.A0(\u_spi2wb.u_if.cmd_reg[5] ),
    .A1(\u_spi2wb.u_if.cmd_reg[4] ),
    .S(_02054_),
    .X(_02056_));
 sky130_fd_sc_hd__clkbuf_1 _05788_ (.A(_02056_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _05789_ (.A0(\u_spi2wb.u_if.cmd_reg[6] ),
    .A1(\u_spi2wb.u_if.cmd_reg[5] ),
    .S(_02054_),
    .X(_02057_));
 sky130_fd_sc_hd__clkbuf_1 _05790_ (.A(_02057_),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _05791_ (.A0(\u_spi2wb.u_if.cmd_reg[7] ),
    .A1(\u_spi2wb.u_if.cmd_reg[6] ),
    .S(_02054_),
    .X(_02058_));
 sky130_fd_sc_hd__clkbuf_1 _05792_ (.A(_02058_),
    .X(_00094_));
 sky130_fd_sc_hd__nor2_4 _05793_ (.A(_01455_),
    .B(_01113_),
    .Y(_02059_));
 sky130_fd_sc_hd__clkbuf_1 _05794_ (.A(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05795_ (.A(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _05796_ (.A0(\u_spi2wb.reg_addr[0] ),
    .A1(net308),
    .S(_02061_),
    .X(_02062_));
 sky130_fd_sc_hd__clkbuf_1 _05797_ (.A(_02062_),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _05798_ (.A0(\u_spi2wb.reg_addr[1] ),
    .A1(\u_spi2wb.reg_addr[0] ),
    .S(_02061_),
    .X(_02063_));
 sky130_fd_sc_hd__clkbuf_1 _05799_ (.A(_02063_),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _05800_ (.A0(\u_spi2wb.reg_addr[2] ),
    .A1(\u_spi2wb.reg_addr[1] ),
    .S(_02061_),
    .X(_02064_));
 sky130_fd_sc_hd__clkbuf_1 _05801_ (.A(_02064_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _05802_ (.A0(\u_spi2wb.reg_addr[3] ),
    .A1(\u_spi2wb.reg_addr[2] ),
    .S(_02061_),
    .X(_02065_));
 sky130_fd_sc_hd__clkbuf_1 _05803_ (.A(_02065_),
    .X(_00098_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05804_ (.A(_02060_),
    .X(_02066_));
 sky130_fd_sc_hd__mux2_1 _05805_ (.A0(\u_spi2wb.reg_addr[4] ),
    .A1(\u_spi2wb.reg_addr[3] ),
    .S(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__clkbuf_1 _05806_ (.A(_02067_),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _05807_ (.A0(\u_spi2wb.reg_addr[5] ),
    .A1(\u_spi2wb.reg_addr[4] ),
    .S(_02066_),
    .X(_02068_));
 sky130_fd_sc_hd__clkbuf_1 _05808_ (.A(_02068_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _05809_ (.A0(\u_spi2wb.reg_addr[6] ),
    .A1(\u_spi2wb.reg_addr[5] ),
    .S(_02066_),
    .X(_02069_));
 sky130_fd_sc_hd__clkbuf_1 _05810_ (.A(_02069_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _05811_ (.A0(\u_spi2wb.reg_addr[7] ),
    .A1(\u_spi2wb.reg_addr[6] ),
    .S(_02066_),
    .X(_02070_));
 sky130_fd_sc_hd__clkbuf_1 _05812_ (.A(_02070_),
    .X(_00102_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05813_ (.A(_02060_),
    .X(_02071_));
 sky130_fd_sc_hd__mux2_1 _05814_ (.A0(\u_spi2wb.reg_addr[8] ),
    .A1(\u_spi2wb.reg_addr[7] ),
    .S(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__clkbuf_1 _05815_ (.A(_02072_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _05816_ (.A0(\u_spi2wb.reg_addr[9] ),
    .A1(\u_spi2wb.reg_addr[8] ),
    .S(_02071_),
    .X(_02073_));
 sky130_fd_sc_hd__clkbuf_1 _05817_ (.A(_02073_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _05818_ (.A0(\u_spi2wb.reg_addr[10] ),
    .A1(\u_spi2wb.reg_addr[9] ),
    .S(_02071_),
    .X(_02074_));
 sky130_fd_sc_hd__clkbuf_1 _05819_ (.A(_02074_),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _05820_ (.A0(\u_spi2wb.reg_addr[11] ),
    .A1(\u_spi2wb.reg_addr[10] ),
    .S(_02071_),
    .X(_02075_));
 sky130_fd_sc_hd__clkbuf_1 _05821_ (.A(_02075_),
    .X(_00106_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05822_ (.A(_02060_),
    .X(_02076_));
 sky130_fd_sc_hd__mux2_1 _05823_ (.A0(\u_spi2wb.reg_addr[12] ),
    .A1(\u_spi2wb.reg_addr[11] ),
    .S(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__clkbuf_1 _05824_ (.A(_02077_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _05825_ (.A0(\u_spi2wb.reg_addr[13] ),
    .A1(\u_spi2wb.reg_addr[12] ),
    .S(_02076_),
    .X(_02078_));
 sky130_fd_sc_hd__clkbuf_1 _05826_ (.A(_02078_),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _05827_ (.A0(\u_spi2wb.reg_addr[14] ),
    .A1(\u_spi2wb.reg_addr[13] ),
    .S(_02076_),
    .X(_02079_));
 sky130_fd_sc_hd__clkbuf_1 _05828_ (.A(_02079_),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _05829_ (.A0(\u_spi2wb.reg_addr[15] ),
    .A1(\u_spi2wb.reg_addr[14] ),
    .S(_02076_),
    .X(_02080_));
 sky130_fd_sc_hd__clkbuf_1 _05830_ (.A(_02080_),
    .X(_00110_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05831_ (.A(_02059_),
    .X(_02081_));
 sky130_fd_sc_hd__mux2_1 _05832_ (.A0(\u_spi2wb.reg_addr[16] ),
    .A1(\u_spi2wb.reg_addr[15] ),
    .S(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__clkbuf_1 _05833_ (.A(_02082_),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _05834_ (.A0(\u_spi2wb.reg_addr[17] ),
    .A1(\u_spi2wb.reg_addr[16] ),
    .S(_02081_),
    .X(_02083_));
 sky130_fd_sc_hd__clkbuf_1 _05835_ (.A(_02083_),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _05836_ (.A0(\u_spi2wb.reg_addr[18] ),
    .A1(\u_spi2wb.reg_addr[17] ),
    .S(_02081_),
    .X(_02084_));
 sky130_fd_sc_hd__clkbuf_1 _05837_ (.A(_02084_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _05838_ (.A0(\u_spi2wb.reg_addr[19] ),
    .A1(\u_spi2wb.reg_addr[18] ),
    .S(_02081_),
    .X(_02085_));
 sky130_fd_sc_hd__clkbuf_1 _05839_ (.A(_02085_),
    .X(_00114_));
 sky130_fd_sc_hd__and2_2 _05840_ (.A(\u_spi2wb.u_if.wr_phase ),
    .B(_01129_),
    .X(_02086_));
 sky130_fd_sc_hd__clkbuf_1 _05841_ (.A(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05842_ (.A(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_1 _05843_ (.A0(\u_spi2wb.reg_wdata[0] ),
    .A1(net308),
    .S(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__clkbuf_1 _05844_ (.A(_02089_),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _05845_ (.A0(\u_spi2wb.reg_wdata[1] ),
    .A1(\u_spi2wb.reg_wdata[0] ),
    .S(_02088_),
    .X(_02090_));
 sky130_fd_sc_hd__clkbuf_1 _05846_ (.A(_02090_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _05847_ (.A0(\u_spi2wb.reg_wdata[2] ),
    .A1(\u_spi2wb.reg_wdata[1] ),
    .S(_02088_),
    .X(_02091_));
 sky130_fd_sc_hd__clkbuf_1 _05848_ (.A(_02091_),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _05849_ (.A0(\u_spi2wb.reg_wdata[3] ),
    .A1(\u_spi2wb.reg_wdata[2] ),
    .S(_02088_),
    .X(_02092_));
 sky130_fd_sc_hd__clkbuf_1 _05850_ (.A(_02092_),
    .X(_00118_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05851_ (.A(_02087_),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_1 _05852_ (.A0(\u_spi2wb.reg_wdata[4] ),
    .A1(\u_spi2wb.reg_wdata[3] ),
    .S(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__clkbuf_1 _05853_ (.A(_02094_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _05854_ (.A0(\u_spi2wb.reg_wdata[5] ),
    .A1(\u_spi2wb.reg_wdata[4] ),
    .S(_02093_),
    .X(_02095_));
 sky130_fd_sc_hd__clkbuf_1 _05855_ (.A(_02095_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _05856_ (.A0(\u_spi2wb.reg_wdata[6] ),
    .A1(\u_spi2wb.reg_wdata[5] ),
    .S(_02093_),
    .X(_02096_));
 sky130_fd_sc_hd__clkbuf_1 _05857_ (.A(_02096_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _05858_ (.A0(\u_spi2wb.reg_wdata[7] ),
    .A1(\u_spi2wb.reg_wdata[6] ),
    .S(_02093_),
    .X(_02097_));
 sky130_fd_sc_hd__clkbuf_1 _05859_ (.A(_02097_),
    .X(_00122_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05860_ (.A(_02087_),
    .X(_02098_));
 sky130_fd_sc_hd__mux2_1 _05861_ (.A0(\u_spi2wb.reg_wdata[8] ),
    .A1(\u_spi2wb.reg_wdata[7] ),
    .S(_02098_),
    .X(_02099_));
 sky130_fd_sc_hd__clkbuf_1 _05862_ (.A(_02099_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _05863_ (.A0(\u_spi2wb.reg_wdata[9] ),
    .A1(\u_spi2wb.reg_wdata[8] ),
    .S(_02098_),
    .X(_02100_));
 sky130_fd_sc_hd__clkbuf_1 _05864_ (.A(_02100_),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _05865_ (.A0(\u_spi2wb.reg_wdata[10] ),
    .A1(\u_spi2wb.reg_wdata[9] ),
    .S(_02098_),
    .X(_02101_));
 sky130_fd_sc_hd__clkbuf_1 _05866_ (.A(_02101_),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _05867_ (.A0(\u_spi2wb.reg_wdata[11] ),
    .A1(\u_spi2wb.reg_wdata[10] ),
    .S(_02098_),
    .X(_02102_));
 sky130_fd_sc_hd__clkbuf_1 _05868_ (.A(_02102_),
    .X(_00126_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05869_ (.A(_02087_),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_1 _05870_ (.A0(\u_spi2wb.reg_wdata[12] ),
    .A1(\u_spi2wb.reg_wdata[11] ),
    .S(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__clkbuf_1 _05871_ (.A(_02104_),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _05872_ (.A0(\u_spi2wb.reg_wdata[13] ),
    .A1(\u_spi2wb.reg_wdata[12] ),
    .S(_02103_),
    .X(_02105_));
 sky130_fd_sc_hd__clkbuf_1 _05873_ (.A(_02105_),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _05874_ (.A0(\u_spi2wb.reg_wdata[14] ),
    .A1(\u_spi2wb.reg_wdata[13] ),
    .S(_02103_),
    .X(_02106_));
 sky130_fd_sc_hd__clkbuf_1 _05875_ (.A(_02106_),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _05876_ (.A0(\u_spi2wb.reg_wdata[15] ),
    .A1(\u_spi2wb.reg_wdata[14] ),
    .S(_02103_),
    .X(_02107_));
 sky130_fd_sc_hd__clkbuf_1 _05877_ (.A(_02107_),
    .X(_00130_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05878_ (.A(_02086_),
    .X(_02108_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05879_ (.A(_02108_),
    .X(_02109_));
 sky130_fd_sc_hd__mux2_1 _05880_ (.A0(\u_spi2wb.reg_wdata[16] ),
    .A1(\u_spi2wb.reg_wdata[15] ),
    .S(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__clkbuf_1 _05881_ (.A(_02110_),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _05882_ (.A0(\u_spi2wb.reg_wdata[17] ),
    .A1(\u_spi2wb.reg_wdata[16] ),
    .S(_02109_),
    .X(_02111_));
 sky130_fd_sc_hd__clkbuf_1 _05883_ (.A(_02111_),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _05884_ (.A0(\u_spi2wb.reg_wdata[18] ),
    .A1(\u_spi2wb.reg_wdata[17] ),
    .S(_02109_),
    .X(_02112_));
 sky130_fd_sc_hd__clkbuf_1 _05885_ (.A(_02112_),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _05886_ (.A0(\u_spi2wb.reg_wdata[19] ),
    .A1(\u_spi2wb.reg_wdata[18] ),
    .S(_02109_),
    .X(_02113_));
 sky130_fd_sc_hd__clkbuf_1 _05887_ (.A(_02113_),
    .X(_00134_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05888_ (.A(_02108_),
    .X(_02114_));
 sky130_fd_sc_hd__mux2_1 _05889_ (.A0(\u_spi2wb.reg_wdata[20] ),
    .A1(\u_spi2wb.reg_wdata[19] ),
    .S(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__clkbuf_1 _05890_ (.A(_02115_),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _05891_ (.A0(\u_spi2wb.reg_wdata[21] ),
    .A1(\u_spi2wb.reg_wdata[20] ),
    .S(_02114_),
    .X(_02116_));
 sky130_fd_sc_hd__clkbuf_1 _05892_ (.A(_02116_),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _05893_ (.A0(\u_spi2wb.reg_wdata[22] ),
    .A1(\u_spi2wb.reg_wdata[21] ),
    .S(_02114_),
    .X(_02117_));
 sky130_fd_sc_hd__clkbuf_1 _05894_ (.A(_02117_),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _05895_ (.A0(\u_spi2wb.reg_wdata[23] ),
    .A1(\u_spi2wb.reg_wdata[22] ),
    .S(_02114_),
    .X(_02118_));
 sky130_fd_sc_hd__clkbuf_1 _05896_ (.A(_02118_),
    .X(_00138_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05897_ (.A(_02108_),
    .X(_02119_));
 sky130_fd_sc_hd__mux2_1 _05898_ (.A0(\u_spi2wb.reg_wdata[24] ),
    .A1(\u_spi2wb.reg_wdata[23] ),
    .S(_02119_),
    .X(_02120_));
 sky130_fd_sc_hd__clkbuf_1 _05899_ (.A(_02120_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _05900_ (.A0(\u_spi2wb.reg_wdata[25] ),
    .A1(\u_spi2wb.reg_wdata[24] ),
    .S(_02119_),
    .X(_02121_));
 sky130_fd_sc_hd__clkbuf_1 _05901_ (.A(_02121_),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _05902_ (.A0(\u_spi2wb.reg_wdata[26] ),
    .A1(\u_spi2wb.reg_wdata[25] ),
    .S(_02119_),
    .X(_02122_));
 sky130_fd_sc_hd__clkbuf_1 _05903_ (.A(_02122_),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _05904_ (.A0(\u_spi2wb.reg_wdata[27] ),
    .A1(\u_spi2wb.reg_wdata[26] ),
    .S(_02119_),
    .X(_02123_));
 sky130_fd_sc_hd__clkbuf_1 _05905_ (.A(_02123_),
    .X(_00142_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05906_ (.A(_02108_),
    .X(_02124_));
 sky130_fd_sc_hd__mux2_1 _05907_ (.A0(\u_spi2wb.reg_wdata[28] ),
    .A1(\u_spi2wb.reg_wdata[27] ),
    .S(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__clkbuf_1 _05908_ (.A(_02125_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _05909_ (.A0(\u_spi2wb.reg_wdata[29] ),
    .A1(\u_spi2wb.reg_wdata[28] ),
    .S(_02124_),
    .X(_02126_));
 sky130_fd_sc_hd__clkbuf_1 _05910_ (.A(_02126_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _05911_ (.A0(\u_spi2wb.reg_wdata[30] ),
    .A1(\u_spi2wb.reg_wdata[29] ),
    .S(_02124_),
    .X(_02127_));
 sky130_fd_sc_hd__clkbuf_1 _05912_ (.A(_02127_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _05913_ (.A0(\u_spi2wb.reg_wdata[31] ),
    .A1(\u_spi2wb.reg_wdata[30] ),
    .S(_02124_),
    .X(_02128_));
 sky130_fd_sc_hd__clkbuf_1 _05914_ (.A(_02128_),
    .X(_00146_));
 sky130_fd_sc_hd__clkbuf_1 _05915_ (.A(\u_reset_fsm.state[0] ),
    .X(_02129_));
 sky130_fd_sc_hd__or3_1 _05916_ (.A(\u_reset_fsm.state[1] ),
    .B(_02129_),
    .C(_01967_),
    .X(_02130_));
 sky130_fd_sc_hd__o22a_1 _05917_ (.A1(\u_reset_fsm.boot_req_ss ),
    .A2(_02012_),
    .B1(_01981_),
    .B2(_02007_),
    .X(_02131_));
 sky130_fd_sc_hd__o21ai_2 _05918_ (.A1(_01980_),
    .A2(_02130_),
    .B1(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__nand2_1 _05919_ (.A(_01962_),
    .B(_02129_),
    .Y(_02133_));
 sky130_fd_sc_hd__clkbuf_1 _05920_ (.A(\u_reset_fsm.state[1] ),
    .X(_02134_));
 sky130_fd_sc_hd__inv_2 _05921_ (.A(_01967_),
    .Y(_02135_));
 sky130_fd_sc_hd__clkbuf_1 _05922_ (.A(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__a21oi_1 _05923_ (.A1(_02134_),
    .A2(_02136_),
    .B1(_02132_),
    .Y(_02137_));
 sky130_fd_sc_hd__clkbuf_1 _05924_ (.A(_02129_),
    .X(_02138_));
 sky130_fd_sc_hd__o22a_1 _05925_ (.A1(_02132_),
    .A2(_02133_),
    .B1(_02137_),
    .B2(_02138_),
    .X(_00147_));
 sky130_fd_sc_hd__o211ai_1 _05926_ (.A1(_02135_),
    .A2(_02133_),
    .B1(_02130_),
    .C1(_02012_),
    .Y(_02139_));
 sky130_fd_sc_hd__mux2_1 _05927_ (.A0(_02139_),
    .A1(_02134_),
    .S(_02132_),
    .X(_02140_));
 sky130_fd_sc_hd__clkbuf_1 _05928_ (.A(_02140_),
    .X(_00148_));
 sky130_fd_sc_hd__o21ai_1 _05929_ (.A1(_02132_),
    .A2(_02133_),
    .B1(_02136_),
    .Y(_00149_));
 sky130_fd_sc_hd__or4_1 _05930_ (.A(_02134_),
    .B(_02138_),
    .C(_02136_),
    .D(_02009_),
    .X(_02141_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05931_ (.A(_01965_),
    .X(_02142_));
 sky130_fd_sc_hd__a21o_1 _05932_ (.A1(\u_reg.force_refclk ),
    .A2(_02141_),
    .B1(_02142_),
    .X(_00150_));
 sky130_fd_sc_hd__inv_2 _05933_ (.A(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__a31o_1 _05934_ (.A1(_02134_),
    .A2(_02012_),
    .A3(_02008_),
    .B1(_02142_),
    .X(_02144_));
 sky130_fd_sc_hd__a22o_1 _05935_ (.A1(\u_reg.clk_enb ),
    .A2(_02143_),
    .B1(_02144_),
    .B2(_02138_),
    .X(_00151_));
 sky130_fd_sc_hd__or2_1 _05936_ (.A(\u_reg.soft_reboot ),
    .B(_02142_),
    .X(_02145_));
 sky130_fd_sc_hd__clkbuf_1 _05937_ (.A(_02145_),
    .X(_00152_));
 sky130_fd_sc_hd__and3_1 _05938_ (.A(_02129_),
    .B(_01967_),
    .C(_02008_),
    .X(_02146_));
 sky130_fd_sc_hd__mux2_1 _05939_ (.A0(_01794_),
    .A1(_01962_),
    .S(_02146_),
    .X(_02147_));
 sky130_fd_sc_hd__clkbuf_1 _05940_ (.A(_02147_),
    .X(_00153_));
 sky130_fd_sc_hd__a41o_1 _05941_ (.A1(_01962_),
    .A2(_02138_),
    .A3(_02136_),
    .A4(_02008_),
    .B1(_01799_),
    .X(_00154_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05942_ (.A(_01737_),
    .X(_02148_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05943_ (.A(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__clkbuf_1 _05944_ (.A(_01481_),
    .X(_02150_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05945_ (.A(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__and2_1 _05946_ (.A(_02151_),
    .B(\u_spi2wb.reg_wdata[8] ),
    .X(_02152_));
 sky130_fd_sc_hd__a221o_1 _05947_ (.A1(wbm_dat_i[8]),
    .A2(_01775_),
    .B1(_02149_),
    .B2(\u_uart2wb.reg_wdata[8] ),
    .C1(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05948_ (.A(net224),
    .X(_02154_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05949_ (.A(_01481_),
    .X(_02155_));
 sky130_fd_sc_hd__inv_2 _05950_ (.A(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__or2_1 _05951_ (.A(\u_arb.gnt[0] ),
    .B(_02155_),
    .X(_02157_));
 sky130_fd_sc_hd__o22a_1 _05952_ (.A1(_02156_),
    .A2(\u_spi2wb.reg_be[1] ),
    .B1(_02157_),
    .B2(wbm_sel_i[1]),
    .X(_02158_));
 sky130_fd_sc_hd__inv_2 _05953_ (.A(_01484_),
    .Y(_02159_));
 sky130_fd_sc_hd__a22o_1 _05954_ (.A1(_01471_),
    .A2(\u_spi2wb.reg_addr[2] ),
    .B1(wbm_adr_i[2]),
    .B2(_01474_),
    .X(_02160_));
 sky130_fd_sc_hd__a21o_2 _05955_ (.A1(\u_uart2wb.reg_addr[2] ),
    .A2(_01480_),
    .B1(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__clkbuf_2 _05956_ (.A(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__and2_1 _05957_ (.A(_01471_),
    .B(\u_spi2wb.reg_addr[3] ),
    .X(_02163_));
 sky130_fd_sc_hd__a221o_2 _05958_ (.A1(wbm_adr_i[3]),
    .A2(_01482_),
    .B1(_01473_),
    .B2(\u_uart2wb.reg_addr[3] ),
    .C1(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__clkbuf_2 _05959_ (.A(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__a22o_1 _05960_ (.A1(_01471_),
    .A2(\u_spi2wb.reg_addr[4] ),
    .B1(wbm_adr_i[4]),
    .B2(_01474_),
    .X(_02166_));
 sky130_fd_sc_hd__a21o_2 _05961_ (.A1(\u_uart2wb.reg_addr[4] ),
    .A2(_01480_),
    .B1(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__clkbuf_2 _05962_ (.A(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__nor3_4 _05963_ (.A(_02162_),
    .B(_02165_),
    .C(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__or3b_1 _05964_ (.A(_01477_),
    .B(_02159_),
    .C_N(_02169_),
    .X(_02170_));
 sky130_fd_sc_hd__clkinv_2 _05965_ (.A(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__and2_1 _05966_ (.A(_02158_),
    .B(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__clkbuf_2 _05967_ (.A(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__mux2_1 _05968_ (.A0(\u_reg.cfg_glb_ctrl[8] ),
    .A1(_02154_),
    .S(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__clkbuf_1 _05969_ (.A(_02174_),
    .X(_00155_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05970_ (.A(_01738_),
    .X(_02175_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05971_ (.A(_02155_),
    .X(_02176_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05972_ (.A(_01734_),
    .X(_02177_));
 sky130_fd_sc_hd__a22o_1 _05973_ (.A1(_02176_),
    .A2(\u_spi2wb.reg_wdata[9] ),
    .B1(wbm_dat_i[9]),
    .B2(_02177_),
    .X(_02178_));
 sky130_fd_sc_hd__a21o_1 _05974_ (.A1(\u_uart2wb.reg_wdata[9] ),
    .A2(_02175_),
    .B1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__clkbuf_1 _05975_ (.A(net223),
    .X(_02180_));
 sky130_fd_sc_hd__clkbuf_2 _05976_ (.A(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__mux2_1 _05977_ (.A0(\u_reg.cfg_glb_ctrl[9] ),
    .A1(_02181_),
    .S(_02173_),
    .X(_02182_));
 sky130_fd_sc_hd__clkbuf_1 _05978_ (.A(_02182_),
    .X(_00156_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05979_ (.A(_02155_),
    .X(_02183_));
 sky130_fd_sc_hd__a22o_1 _05980_ (.A1(_02183_),
    .A2(\u_spi2wb.reg_wdata[10] ),
    .B1(wbm_dat_i[10]),
    .B2(_02177_),
    .X(_02184_));
 sky130_fd_sc_hd__a21o_1 _05981_ (.A1(\u_uart2wb.reg_wdata[10] ),
    .A2(_02175_),
    .B1(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__clkbuf_1 _05982_ (.A(net222),
    .X(_02186_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05983_ (.A(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _05984_ (.A0(\u_reg.cfg_glb_ctrl[10] ),
    .A1(_02187_),
    .S(_02173_),
    .X(_02188_));
 sky130_fd_sc_hd__clkbuf_1 _05985_ (.A(_02188_),
    .X(_00157_));
 sky130_fd_sc_hd__and2_1 _05986_ (.A(_02151_),
    .B(\u_spi2wb.reg_wdata[11] ),
    .X(_02189_));
 sky130_fd_sc_hd__a221o_1 _05987_ (.A1(wbm_dat_i[11]),
    .A2(_01775_),
    .B1(_02149_),
    .B2(\u_uart2wb.reg_wdata[11] ),
    .C1(_02189_),
    .X(_02190_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05988_ (.A(net221),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _05989_ (.A0(\u_reg.cfg_glb_ctrl[11] ),
    .A1(_02191_),
    .S(_02173_),
    .X(_02192_));
 sky130_fd_sc_hd__clkbuf_1 _05990_ (.A(_02192_),
    .X(_00158_));
 sky130_fd_sc_hd__clkbuf_1 _05991_ (.A(_01482_),
    .X(_02193_));
 sky130_fd_sc_hd__clkbuf_2 _05992_ (.A(_02193_),
    .X(_02194_));
 sky130_fd_sc_hd__clkbuf_2 _05993_ (.A(_01738_),
    .X(_02195_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05994_ (.A(_01728_),
    .X(_02196_));
 sky130_fd_sc_hd__and2_1 _05995_ (.A(_02196_),
    .B(\u_spi2wb.reg_wdata[12] ),
    .X(_02197_));
 sky130_fd_sc_hd__a221o_1 _05996_ (.A1(wbm_dat_i[12]),
    .A2(_02194_),
    .B1(_02195_),
    .B2(\u_uart2wb.reg_wdata[12] ),
    .C1(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__clkbuf_1 _05997_ (.A(net220),
    .X(_02199_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _05998_ (.A(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__clkbuf_2 _05999_ (.A(_02172_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _06000_ (.A0(\u_reg.cfg_glb_ctrl[12] ),
    .A1(_02200_),
    .S(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__clkbuf_1 _06001_ (.A(_02202_),
    .X(_00159_));
 sky130_fd_sc_hd__and2_1 _06002_ (.A(_02150_),
    .B(\u_spi2wb.reg_wdata[13] ),
    .X(_02203_));
 sky130_fd_sc_hd__a221o_1 _06003_ (.A1(wbm_dat_i[13]),
    .A2(_01774_),
    .B1(_02148_),
    .B2(\u_uart2wb.reg_wdata[13] ),
    .C1(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__clkbuf_1 _06004_ (.A(net229),
    .X(_02205_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06005_ (.A(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _06006_ (.A0(\u_reg.cfg_glb_ctrl[13] ),
    .A1(_02206_),
    .S(_02201_),
    .X(_02207_));
 sky130_fd_sc_hd__clkbuf_1 _06007_ (.A(_02207_),
    .X(_00160_));
 sky130_fd_sc_hd__a22o_1 _06008_ (.A1(_02183_),
    .A2(\u_spi2wb.reg_wdata[14] ),
    .B1(wbm_dat_i[14]),
    .B2(_02177_),
    .X(_02208_));
 sky130_fd_sc_hd__a21o_1 _06009_ (.A1(\u_uart2wb.reg_wdata[14] ),
    .A2(_02175_),
    .B1(_02208_),
    .X(_02209_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06010_ (.A(net219),
    .X(_02210_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06011_ (.A(_02210_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _06012_ (.A0(\u_reg.cfg_glb_ctrl[14] ),
    .A1(_02211_),
    .S(_02201_),
    .X(_02212_));
 sky130_fd_sc_hd__clkbuf_1 _06013_ (.A(_02212_),
    .X(_00161_));
 sky130_fd_sc_hd__clkbuf_2 _06014_ (.A(_01774_),
    .X(_02213_));
 sky130_fd_sc_hd__and2_1 _06015_ (.A(_02151_),
    .B(\u_spi2wb.reg_wdata[15] ),
    .X(_02214_));
 sky130_fd_sc_hd__a221o_4 _06016_ (.A1(wbm_dat_i[15]),
    .A2(_02213_),
    .B1(_02149_),
    .B2(\u_uart2wb.reg_wdata[15] ),
    .C1(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__clkbuf_1 _06017_ (.A(_02215_),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _06018_ (.A0(\u_reg.cfg_glb_ctrl[15] ),
    .A1(_02216_),
    .S(_02201_),
    .X(_02217_));
 sky130_fd_sc_hd__clkbuf_1 _06019_ (.A(_02217_),
    .X(_00162_));
 sky130_fd_sc_hd__clkbuf_1 _06020_ (.A(\u_async_wb.m_cmd_wr_data[61] ),
    .X(_02218_));
 sky130_fd_sc_hd__and2_1 _06021_ (.A(wb_req),
    .B(_01476_),
    .X(_02219_));
 sky130_fd_sc_hd__nor3b_2 _06022_ (.A(_02165_),
    .B(_02168_),
    .C_N(_02162_),
    .Y(_02220_));
 sky130_fd_sc_hd__and3_2 _06023_ (.A(_02219_),
    .B(_01485_),
    .C(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__clkbuf_2 _06024_ (.A(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _06025_ (.A0(_02218_),
    .A1(_02154_),
    .S(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__clkbuf_1 _06026_ (.A(_02223_),
    .X(_00163_));
 sky130_fd_sc_hd__clkbuf_1 _06027_ (.A(\u_async_wb.m_cmd_wr_data[60] ),
    .X(_02224_));
 sky130_fd_sc_hd__and2_1 _06028_ (.A(_02196_),
    .B(\u_spi2wb.reg_wdata[7] ),
    .X(_02225_));
 sky130_fd_sc_hd__a221o_1 _06029_ (.A1(wbm_dat_i[7]),
    .A2(_02194_),
    .B1(_02195_),
    .B2(\u_uart2wb.reg_wdata[7] ),
    .C1(_02225_),
    .X(_02226_));
 sky130_fd_sc_hd__clkbuf_1 _06030_ (.A(net218),
    .X(_02227_));
 sky130_fd_sc_hd__clkbuf_2 _06031_ (.A(_02227_),
    .X(_02228_));
 sky130_fd_sc_hd__mux2_1 _06032_ (.A0(_02224_),
    .A1(_02228_),
    .S(_02222_),
    .X(_02229_));
 sky130_fd_sc_hd__clkbuf_1 _06033_ (.A(_02229_),
    .X(_00164_));
 sky130_fd_sc_hd__clkbuf_1 _06034_ (.A(\u_async_wb.m_cmd_wr_data[59] ),
    .X(_02230_));
 sky130_fd_sc_hd__and2_1 _06035_ (.A(_02176_),
    .B(\u_spi2wb.reg_wdata[6] ),
    .X(_02231_));
 sky130_fd_sc_hd__a221o_1 _06036_ (.A1(wbm_dat_i[6]),
    .A2(_02213_),
    .B1(_02149_),
    .B2(\u_uart2wb.reg_wdata[6] ),
    .C1(_02231_),
    .X(_02232_));
 sky130_fd_sc_hd__clkbuf_2 _06037_ (.A(net217),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _06038_ (.A0(_02230_),
    .A1(_02233_),
    .S(_02222_),
    .X(_02234_));
 sky130_fd_sc_hd__clkbuf_1 _06039_ (.A(_02234_),
    .X(_00165_));
 sky130_fd_sc_hd__clkbuf_1 _06040_ (.A(\u_async_wb.m_cmd_wr_data[58] ),
    .X(_02235_));
 sky130_fd_sc_hd__and2_1 _06041_ (.A(_02150_),
    .B(\u_spi2wb.reg_wdata[5] ),
    .X(_02236_));
 sky130_fd_sc_hd__a221o_1 _06042_ (.A1(wbm_dat_i[5]),
    .A2(_01774_),
    .B1(_02148_),
    .B2(\u_uart2wb.reg_wdata[5] ),
    .C1(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06043_ (.A(net228),
    .X(_02238_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06044_ (.A(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _06045_ (.A0(_02235_),
    .A1(_02239_),
    .S(_02222_),
    .X(_02240_));
 sky130_fd_sc_hd__clkbuf_1 _06046_ (.A(_02240_),
    .X(_00166_));
 sky130_fd_sc_hd__clkbuf_1 _06047_ (.A(\u_async_wb.m_cmd_wr_data[57] ),
    .X(_02241_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06048_ (.A(_01737_),
    .X(_02242_));
 sky130_fd_sc_hd__and2_1 _06049_ (.A(_02196_),
    .B(\u_spi2wb.reg_wdata[4] ),
    .X(_02243_));
 sky130_fd_sc_hd__a221o_1 _06050_ (.A1(wbm_dat_i[4]),
    .A2(_02194_),
    .B1(_02242_),
    .B2(\u_uart2wb.reg_wdata[4] ),
    .C1(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__clkbuf_1 _06051_ (.A(net227),
    .X(_02245_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06052_ (.A(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__clkbuf_2 _06053_ (.A(_02221_),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _06054_ (.A0(_02241_),
    .A1(_02246_),
    .S(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__clkbuf_1 _06055_ (.A(_02248_),
    .X(_00167_));
 sky130_fd_sc_hd__clkbuf_1 _06056_ (.A(\u_async_wb.m_cmd_wr_data[56] ),
    .X(_02249_));
 sky130_fd_sc_hd__clkbuf_2 _06057_ (.A(_01738_),
    .X(_02250_));
 sky130_fd_sc_hd__a22o_1 _06058_ (.A1(_02183_),
    .A2(\u_spi2wb.reg_wdata[3] ),
    .B1(wbm_dat_i[3]),
    .B2(_01735_),
    .X(_02251_));
 sky130_fd_sc_hd__a21o_1 _06059_ (.A1(\u_uart2wb.reg_wdata[3] ),
    .A2(_02250_),
    .B1(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__clkbuf_1 _06060_ (.A(net216),
    .X(_02253_));
 sky130_fd_sc_hd__clkbuf_2 _06061_ (.A(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _06062_ (.A0(_02249_),
    .A1(_02254_),
    .S(_02247_),
    .X(_02255_));
 sky130_fd_sc_hd__clkbuf_1 _06063_ (.A(_02255_),
    .X(_00168_));
 sky130_fd_sc_hd__a22o_1 _06064_ (.A1(_02183_),
    .A2(\u_spi2wb.reg_wdata[2] ),
    .B1(wbm_dat_i[2]),
    .B2(_02177_),
    .X(_02256_));
 sky130_fd_sc_hd__a21o_1 _06065_ (.A1(\u_uart2wb.reg_wdata[2] ),
    .A2(_02175_),
    .B1(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__clkbuf_1 _06066_ (.A(net215),
    .X(_02258_));
 sky130_fd_sc_hd__clkbuf_2 _06067_ (.A(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _06068_ (.A0(\u_reg.u_bank_sel.gen_bit_reg[2].u_bit_reg.data_out ),
    .A1(_02259_),
    .S(_02247_),
    .X(_02260_));
 sky130_fd_sc_hd__clkbuf_1 _06069_ (.A(_02260_),
    .X(_00169_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06070_ (.A(_02193_),
    .X(_02261_));
 sky130_fd_sc_hd__clkbuf_1 _06071_ (.A(_01728_),
    .X(_02262_));
 sky130_fd_sc_hd__and2_1 _06072_ (.A(_02262_),
    .B(\u_spi2wb.reg_wdata[1] ),
    .X(_02263_));
 sky130_fd_sc_hd__a221o_1 _06073_ (.A1(wbm_dat_i[1]),
    .A2(_02261_),
    .B1(_02242_),
    .B2(\u_uart2wb.reg_wdata[1] ),
    .C1(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__clkbuf_1 _06074_ (.A(net226),
    .X(_02265_));
 sky130_fd_sc_hd__clkbuf_2 _06075_ (.A(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _06076_ (.A0(\u_reg.u_bank_sel.gen_bit_reg[1].u_bit_reg.data_out ),
    .A1(_02266_),
    .S(_02247_),
    .X(_02267_));
 sky130_fd_sc_hd__clkbuf_1 _06077_ (.A(_02267_),
    .X(_00170_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06078_ (.A(\u_async_wb.m_cmd_wr_data[68] ),
    .X(_02268_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06079_ (.A(_02221_),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _06080_ (.A0(_02268_),
    .A1(_02216_),
    .S(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__clkbuf_1 _06081_ (.A(_02270_),
    .X(_00171_));
 sky130_fd_sc_hd__clkbuf_1 _06082_ (.A(\u_async_wb.m_cmd_wr_data[67] ),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _06083_ (.A0(_02271_),
    .A1(_02210_),
    .S(_02269_),
    .X(_02272_));
 sky130_fd_sc_hd__clkbuf_1 _06084_ (.A(_02272_),
    .X(_00172_));
 sky130_fd_sc_hd__clkbuf_1 _06085_ (.A(\u_async_wb.m_cmd_wr_data[66] ),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _06086_ (.A0(_02273_),
    .A1(_02206_),
    .S(_02269_),
    .X(_02274_));
 sky130_fd_sc_hd__clkbuf_1 _06087_ (.A(_02274_),
    .X(_00173_));
 sky130_fd_sc_hd__clkbuf_1 _06088_ (.A(\u_async_wb.m_cmd_wr_data[65] ),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _06089_ (.A0(_02275_),
    .A1(_02199_),
    .S(_02269_),
    .X(_02276_));
 sky130_fd_sc_hd__clkbuf_1 _06090_ (.A(_02276_),
    .X(_00174_));
 sky130_fd_sc_hd__clkbuf_1 _06091_ (.A(\u_async_wb.m_cmd_wr_data[64] ),
    .X(_02277_));
 sky130_fd_sc_hd__clkbuf_2 _06092_ (.A(_02221_),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _06093_ (.A0(_02277_),
    .A1(_02191_),
    .S(_02278_),
    .X(_02279_));
 sky130_fd_sc_hd__clkbuf_1 _06094_ (.A(_02279_),
    .X(_00175_));
 sky130_fd_sc_hd__clkbuf_1 _06095_ (.A(\u_async_wb.m_cmd_wr_data[63] ),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _06096_ (.A0(_02280_),
    .A1(_02186_),
    .S(_02278_),
    .X(_02281_));
 sky130_fd_sc_hd__clkbuf_1 _06097_ (.A(_02281_),
    .X(_00176_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06098_ (.A(_02193_),
    .X(_02282_));
 sky130_fd_sc_hd__and2_1 _06099_ (.A(_02262_),
    .B(\u_spi2wb.reg_wdata[0] ),
    .X(_02283_));
 sky130_fd_sc_hd__a221o_1 _06100_ (.A1(wbm_dat_i[0]),
    .A2(_02282_),
    .B1(_02242_),
    .B2(\u_uart2wb.reg_wdata[0] ),
    .C1(_02283_),
    .X(_02284_));
 sky130_fd_sc_hd__clkbuf_1 _06101_ (.A(net225),
    .X(_02285_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06102_ (.A(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _06103_ (.A0(\u_reg.u_bank_sel.gen_bit_reg[0].u_bit_reg.data_out ),
    .A1(_02286_),
    .S(_02278_),
    .X(_02287_));
 sky130_fd_sc_hd__clkbuf_1 _06104_ (.A(_02287_),
    .X(_00177_));
 sky130_fd_sc_hd__and3b_2 _06105_ (.A_N(_02164_),
    .B(_02167_),
    .C(_02161_),
    .X(_02288_));
 sky130_fd_sc_hd__and3_2 _06106_ (.A(_02219_),
    .B(_01484_),
    .C(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06107_ (.A(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06108_ (.A(_02290_),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _06109_ (.A0(net73),
    .A1(net225),
    .S(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _06110_ (.A0(strap_sticky[0]),
    .A1(_02292_),
    .S(_01794_),
    .X(_02293_));
 sky130_fd_sc_hd__clkbuf_1 _06111_ (.A(_02293_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _06112_ (.A0(net84),
    .A1(net226),
    .S(_02291_),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _06113_ (.A0(strap_sticky[1]),
    .A1(_02294_),
    .S(_01794_),
    .X(_02295_));
 sky130_fd_sc_hd__clkbuf_1 _06114_ (.A(_02295_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _06115_ (.A0(net95),
    .A1(net215),
    .S(_02291_),
    .X(_02296_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06116_ (.A(_01793_),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _06117_ (.A0(strap_sticky[2]),
    .A1(_02296_),
    .S(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__clkbuf_1 _06118_ (.A(_02298_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _06119_ (.A0(net98),
    .A1(net216),
    .S(_02291_),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _06120_ (.A0(strap_sticky[3]),
    .A1(_02299_),
    .S(_02297_),
    .X(_02300_));
 sky130_fd_sc_hd__clkbuf_1 _06121_ (.A(_02300_),
    .X(_00181_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06122_ (.A(_02290_),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _06123_ (.A0(net99),
    .A1(net227),
    .S(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__mux2_1 _06124_ (.A0(strap_sticky[4]),
    .A1(_02302_),
    .S(_02297_),
    .X(_02303_));
 sky130_fd_sc_hd__clkbuf_1 _06125_ (.A(_02303_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _06126_ (.A0(net100),
    .A1(net228),
    .S(_02301_),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _06127_ (.A0(strap_sticky[5]),
    .A1(_02304_),
    .S(_02297_),
    .X(_02305_));
 sky130_fd_sc_hd__clkbuf_1 _06128_ (.A(_02305_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _06129_ (.A0(net101),
    .A1(net217),
    .S(_02301_),
    .X(_02306_));
 sky130_fd_sc_hd__clkbuf_1 _06130_ (.A(net304),
    .X(_02307_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06131_ (.A(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__mux2_1 _06132_ (.A0(strap_sticky[6]),
    .A1(_02306_),
    .S(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__clkbuf_1 _06133_ (.A(_02309_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _06134_ (.A0(net102),
    .A1(net218),
    .S(_02301_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _06135_ (.A0(strap_sticky[7]),
    .A1(_02310_),
    .S(_02308_),
    .X(_02311_));
 sky130_fd_sc_hd__clkbuf_1 _06136_ (.A(_02311_),
    .X(_00185_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06137_ (.A(_02290_),
    .X(_02312_));
 sky130_fd_sc_hd__mux2_1 _06138_ (.A0(net103),
    .A1(net224),
    .S(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _06139_ (.A0(strap_sticky[8]),
    .A1(_02313_),
    .S(_02308_),
    .X(_02314_));
 sky130_fd_sc_hd__clkbuf_1 _06140_ (.A(_02314_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _06141_ (.A0(net104),
    .A1(net223),
    .S(_02312_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _06142_ (.A0(strap_sticky[9]),
    .A1(_02315_),
    .S(_02308_),
    .X(_02316_));
 sky130_fd_sc_hd__clkbuf_1 _06143_ (.A(_02316_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _06144_ (.A0(net74),
    .A1(net222),
    .S(_02312_),
    .X(_02317_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06145_ (.A(_02307_),
    .X(_02318_));
 sky130_fd_sc_hd__mux2_1 _06146_ (.A0(strap_sticky[10]),
    .A1(_02317_),
    .S(_02318_),
    .X(_02319_));
 sky130_fd_sc_hd__clkbuf_1 _06147_ (.A(_02319_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _06148_ (.A0(net75),
    .A1(net221),
    .S(_02312_),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _06149_ (.A0(strap_sticky[11]),
    .A1(_02320_),
    .S(_02318_),
    .X(_02321_));
 sky130_fd_sc_hd__clkbuf_1 _06150_ (.A(_02321_),
    .X(_00189_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06151_ (.A(_02290_),
    .X(_02322_));
 sky130_fd_sc_hd__mux2_1 _06152_ (.A0(net76),
    .A1(net220),
    .S(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _06153_ (.A0(strap_sticky[12]),
    .A1(_02323_),
    .S(_02318_),
    .X(_02324_));
 sky130_fd_sc_hd__clkbuf_1 _06154_ (.A(_02324_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _06155_ (.A0(net77),
    .A1(net229),
    .S(_02322_),
    .X(_02325_));
 sky130_fd_sc_hd__mux2_1 _06156_ (.A0(strap_sticky[13]),
    .A1(_02325_),
    .S(_02318_),
    .X(_02326_));
 sky130_fd_sc_hd__clkbuf_1 _06157_ (.A(_02326_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _06158_ (.A0(net78),
    .A1(net219),
    .S(_02322_),
    .X(_02327_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06159_ (.A(_02307_),
    .X(_02328_));
 sky130_fd_sc_hd__mux2_1 _06160_ (.A0(strap_sticky[14]),
    .A1(_02327_),
    .S(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__clkbuf_1 _06161_ (.A(_02329_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _06162_ (.A0(net79),
    .A1(_02215_),
    .S(_02322_),
    .X(_02330_));
 sky130_fd_sc_hd__mux2_1 _06163_ (.A0(strap_sticky[15]),
    .A1(_02330_),
    .S(_02328_),
    .X(_02331_));
 sky130_fd_sc_hd__clkbuf_1 _06164_ (.A(_02331_),
    .X(_00193_));
 sky130_fd_sc_hd__and2_1 _06165_ (.A(_02196_),
    .B(\u_spi2wb.reg_wdata[16] ),
    .X(_02332_));
 sky130_fd_sc_hd__a221o_4 _06166_ (.A1(wbm_dat_i[16]),
    .A2(_02194_),
    .B1(_02195_),
    .B2(\u_uart2wb.reg_wdata[16] ),
    .C1(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__clkbuf_1 _06167_ (.A(_02289_),
    .X(_02334_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06168_ (.A(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _06169_ (.A0(net80),
    .A1(_02333_),
    .S(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__mux2_1 _06170_ (.A0(strap_sticky[16]),
    .A1(_02336_),
    .S(_02328_),
    .X(_02337_));
 sky130_fd_sc_hd__clkbuf_1 _06171_ (.A(_02337_),
    .X(_00194_));
 sky130_fd_sc_hd__clkbuf_2 _06172_ (.A(_01734_),
    .X(_02338_));
 sky130_fd_sc_hd__and2_1 _06173_ (.A(_02262_),
    .B(\u_spi2wb.reg_wdata[17] ),
    .X(_02339_));
 sky130_fd_sc_hd__a221o_4 _06174_ (.A1(wbm_dat_i[17]),
    .A2(_02338_),
    .B1(_02242_),
    .B2(\u_uart2wb.reg_wdata[17] ),
    .C1(_02339_),
    .X(_02340_));
 sky130_fd_sc_hd__mux2_1 _06175_ (.A0(net81),
    .A1(_02340_),
    .S(_02335_),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _06176_ (.A0(strap_sticky[17]),
    .A1(_02341_),
    .S(_02328_),
    .X(_02342_));
 sky130_fd_sc_hd__clkbuf_1 _06177_ (.A(_02342_),
    .X(_00195_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06178_ (.A(_01737_),
    .X(_02343_));
 sky130_fd_sc_hd__and2_1 _06179_ (.A(_02262_),
    .B(\u_spi2wb.reg_wdata[18] ),
    .X(_02344_));
 sky130_fd_sc_hd__a221o_4 _06180_ (.A1(wbm_dat_i[18]),
    .A2(_02338_),
    .B1(_02343_),
    .B2(\u_uart2wb.reg_wdata[18] ),
    .C1(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__mux2_1 _06181_ (.A0(net82),
    .A1(_02345_),
    .S(_02335_),
    .X(_02346_));
 sky130_fd_sc_hd__clkbuf_2 _06182_ (.A(_02307_),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _06183_ (.A0(strap_sticky[18]),
    .A1(_02346_),
    .S(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__clkbuf_1 _06184_ (.A(_02348_),
    .X(_00196_));
 sky130_fd_sc_hd__clkbuf_1 _06185_ (.A(_01728_),
    .X(_02349_));
 sky130_fd_sc_hd__a22o_1 _06186_ (.A1(_02349_),
    .A2(\u_spi2wb.reg_wdata[19] ),
    .B1(wbm_dat_i[19]),
    .B2(_02193_),
    .X(_02350_));
 sky130_fd_sc_hd__a21o_4 _06187_ (.A1(\u_uart2wb.reg_wdata[19] ),
    .A2(_02195_),
    .B1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__mux2_1 _06188_ (.A0(net83),
    .A1(_02351_),
    .S(_02335_),
    .X(_02352_));
 sky130_fd_sc_hd__mux2_1 _06189_ (.A0(strap_sticky[19]),
    .A1(_02352_),
    .S(_02347_),
    .X(_02353_));
 sky130_fd_sc_hd__clkbuf_1 _06190_ (.A(_02353_),
    .X(_00197_));
 sky130_fd_sc_hd__a22o_1 _06191_ (.A1(_02349_),
    .A2(\u_spi2wb.reg_wdata[20] ),
    .B1(wbm_dat_i[20]),
    .B2(_01735_),
    .X(_02354_));
 sky130_fd_sc_hd__a21o_2 _06192_ (.A1(\u_uart2wb.reg_wdata[20] ),
    .A2(_02250_),
    .B1(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06193_ (.A(_02334_),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _06194_ (.A0(net85),
    .A1(_02355_),
    .S(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__mux2_1 _06195_ (.A0(strap_sticky[20]),
    .A1(_02357_),
    .S(_02347_),
    .X(_02358_));
 sky130_fd_sc_hd__clkbuf_1 _06196_ (.A(_02358_),
    .X(_00198_));
 sky130_fd_sc_hd__and2_1 _06197_ (.A(_01729_),
    .B(\u_spi2wb.reg_wdata[21] ),
    .X(_02359_));
 sky130_fd_sc_hd__a221o_4 _06198_ (.A1(wbm_dat_i[21]),
    .A2(_02338_),
    .B1(_02343_),
    .B2(\u_uart2wb.reg_wdata[21] ),
    .C1(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__mux2_1 _06199_ (.A0(net86),
    .A1(_02360_),
    .S(_02356_),
    .X(_02361_));
 sky130_fd_sc_hd__mux2_1 _06200_ (.A0(strap_sticky[21]),
    .A1(_02361_),
    .S(_02347_),
    .X(_02362_));
 sky130_fd_sc_hd__clkbuf_1 _06201_ (.A(_02362_),
    .X(_00199_));
 sky130_fd_sc_hd__a22o_1 _06202_ (.A1(_02349_),
    .A2(\u_spi2wb.reg_wdata[22] ),
    .B1(wbm_dat_i[22]),
    .B2(_01735_),
    .X(_02363_));
 sky130_fd_sc_hd__a21o_4 _06203_ (.A1(\u_uart2wb.reg_wdata[22] ),
    .A2(_02250_),
    .B1(_02363_),
    .X(_02364_));
 sky130_fd_sc_hd__mux2_1 _06204_ (.A0(net87),
    .A1(_02364_),
    .S(_02356_),
    .X(_02365_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06205_ (.A(net304),
    .X(_02366_));
 sky130_fd_sc_hd__mux2_1 _06206_ (.A0(strap_sticky[22]),
    .A1(_02365_),
    .S(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__clkbuf_1 _06207_ (.A(_02367_),
    .X(_00200_));
 sky130_fd_sc_hd__and2_1 _06208_ (.A(_02150_),
    .B(\u_spi2wb.reg_wdata[23] ),
    .X(_02368_));
 sky130_fd_sc_hd__a221o_4 _06209_ (.A1(wbm_dat_i[23]),
    .A2(_02338_),
    .B1(_02148_),
    .B2(\u_uart2wb.reg_wdata[23] ),
    .C1(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__mux2_1 _06210_ (.A0(net88),
    .A1(_02369_),
    .S(_02356_),
    .X(_02370_));
 sky130_fd_sc_hd__mux2_1 _06211_ (.A0(strap_sticky[23]),
    .A1(_02370_),
    .S(_02366_),
    .X(_02371_));
 sky130_fd_sc_hd__clkbuf_1 _06212_ (.A(_02371_),
    .X(_00201_));
 sky130_fd_sc_hd__clkbuf_2 _06213_ (.A(_02343_),
    .X(_02372_));
 sky130_fd_sc_hd__a22o_1 _06214_ (.A1(_01730_),
    .A2(\u_spi2wb.reg_wdata[24] ),
    .B1(wbm_dat_i[24]),
    .B2(_02282_),
    .X(_02373_));
 sky130_fd_sc_hd__a21o_4 _06215_ (.A1(\u_uart2wb.reg_wdata[24] ),
    .A2(_02372_),
    .B1(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06216_ (.A(_02334_),
    .X(_02375_));
 sky130_fd_sc_hd__mux2_1 _06217_ (.A0(net89),
    .A1(_02374_),
    .S(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _06218_ (.A0(strap_sticky[24]),
    .A1(_02376_),
    .S(_02366_),
    .X(_02377_));
 sky130_fd_sc_hd__clkbuf_1 _06219_ (.A(_02377_),
    .X(_00202_));
 sky130_fd_sc_hd__clkbuf_1 _06220_ (.A(_01729_),
    .X(_02378_));
 sky130_fd_sc_hd__a22o_1 _06221_ (.A1(_02378_),
    .A2(\u_spi2wb.reg_wdata[25] ),
    .B1(wbm_dat_i[25]),
    .B2(_02282_),
    .X(_02379_));
 sky130_fd_sc_hd__a21o_4 _06222_ (.A1(\u_uart2wb.reg_wdata[25] ),
    .A2(_02372_),
    .B1(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _06223_ (.A0(net90),
    .A1(_02380_),
    .S(_02375_),
    .X(_02381_));
 sky130_fd_sc_hd__mux2_1 _06224_ (.A0(strap_sticky[25]),
    .A1(_02381_),
    .S(_02366_),
    .X(_02382_));
 sky130_fd_sc_hd__clkbuf_1 _06225_ (.A(_02382_),
    .X(_00203_));
 sky130_fd_sc_hd__clkbuf_2 _06226_ (.A(_02343_),
    .X(_02383_));
 sky130_fd_sc_hd__a22o_1 _06227_ (.A1(_02378_),
    .A2(\u_spi2wb.reg_wdata[26] ),
    .B1(wbm_dat_i[26]),
    .B2(_02282_),
    .X(_02384_));
 sky130_fd_sc_hd__a21o_4 _06228_ (.A1(\u_uart2wb.reg_wdata[26] ),
    .A2(_02383_),
    .B1(_02384_),
    .X(_02385_));
 sky130_fd_sc_hd__mux2_1 _06229_ (.A0(net91),
    .A1(_02385_),
    .S(_02375_),
    .X(_02386_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06230_ (.A(net304),
    .X(_02387_));
 sky130_fd_sc_hd__mux2_1 _06231_ (.A0(strap_sticky[26]),
    .A1(_02386_),
    .S(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__clkbuf_1 _06232_ (.A(_02388_),
    .X(_00204_));
 sky130_fd_sc_hd__and2_1 _06233_ (.A(_02176_),
    .B(\u_spi2wb.reg_wdata[27] ),
    .X(_02389_));
 sky130_fd_sc_hd__a221o_4 _06234_ (.A1(wbm_dat_i[27]),
    .A2(_02213_),
    .B1(_01739_),
    .B2(\u_uart2wb.reg_wdata[27] ),
    .C1(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__mux2_1 _06235_ (.A0(net92),
    .A1(_02390_),
    .S(_02375_),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_1 _06236_ (.A0(strap_sticky[27]),
    .A1(_02391_),
    .S(_02387_),
    .X(_02392_));
 sky130_fd_sc_hd__clkbuf_1 _06237_ (.A(_02392_),
    .X(_00205_));
 sky130_fd_sc_hd__a22o_1 _06238_ (.A1(_02378_),
    .A2(\u_spi2wb.reg_wdata[28] ),
    .B1(wbm_dat_i[28]),
    .B2(_02261_),
    .X(_02393_));
 sky130_fd_sc_hd__a21o_4 _06239_ (.A1(\u_uart2wb.reg_wdata[28] ),
    .A2(_02383_),
    .B1(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06240_ (.A(_02334_),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _06241_ (.A0(net93),
    .A1(_02394_),
    .S(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__mux2_1 _06242_ (.A0(strap_sticky[28]),
    .A1(_02396_),
    .S(_02387_),
    .X(_02397_));
 sky130_fd_sc_hd__clkbuf_1 _06243_ (.A(_02397_),
    .X(_00206_));
 sky130_fd_sc_hd__and2_1 _06244_ (.A(_02176_),
    .B(\u_spi2wb.reg_wdata[29] ),
    .X(_02398_));
 sky130_fd_sc_hd__a221o_4 _06245_ (.A1(wbm_dat_i[29]),
    .A2(_02213_),
    .B1(_01739_),
    .B2(\u_uart2wb.reg_wdata[29] ),
    .C1(_02398_),
    .X(_02399_));
 sky130_fd_sc_hd__mux2_1 _06246_ (.A0(net94),
    .A1(_02399_),
    .S(_02395_),
    .X(_02400_));
 sky130_fd_sc_hd__mux2_1 _06247_ (.A0(strap_sticky[29]),
    .A1(_02400_),
    .S(_02387_),
    .X(_02401_));
 sky130_fd_sc_hd__clkbuf_1 _06248_ (.A(_02401_),
    .X(_00207_));
 sky130_fd_sc_hd__a22o_1 _06249_ (.A1(_02378_),
    .A2(\u_spi2wb.reg_wdata[30] ),
    .B1(wbm_dat_i[30]),
    .B2(_02261_),
    .X(_02402_));
 sky130_fd_sc_hd__a21o_4 _06250_ (.A1(\u_uart2wb.reg_wdata[30] ),
    .A2(_02383_),
    .B1(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__mux2_1 _06251_ (.A0(net96),
    .A1(_02403_),
    .S(_02395_),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _06252_ (.A0(strap_sticky[30]),
    .A1(_02404_),
    .S(_01793_),
    .X(_02405_));
 sky130_fd_sc_hd__clkbuf_1 _06253_ (.A(_02405_),
    .X(_00208_));
 sky130_fd_sc_hd__a22o_1 _06254_ (.A1(_02151_),
    .A2(\u_spi2wb.reg_wdata[31] ),
    .B1(wbm_dat_i[31]),
    .B2(_02261_),
    .X(_02406_));
 sky130_fd_sc_hd__a21o_4 _06255_ (.A1(\u_uart2wb.reg_wdata[31] ),
    .A2(_02383_),
    .B1(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _06256_ (.A0(net97),
    .A1(_02407_),
    .S(_02395_),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _06257_ (.A0(\u_reg.soft_reboot ),
    .A1(_02408_),
    .S(_01793_),
    .X(_02409_));
 sky130_fd_sc_hd__clkbuf_1 _06258_ (.A(_02409_),
    .X(_00209_));
 sky130_fd_sc_hd__clkbuf_1 _06259_ (.A(\u_async_wb.m_cmd_wr_data[62] ),
    .X(_02410_));
 sky130_fd_sc_hd__mux2_1 _06260_ (.A0(_02410_),
    .A1(_02180_),
    .S(_02278_),
    .X(_02411_));
 sky130_fd_sc_hd__clkbuf_1 _06261_ (.A(_02411_),
    .X(_00210_));
 sky130_fd_sc_hd__clkbuf_1 _06262_ (.A(_02333_),
    .X(_02412_));
 sky130_fd_sc_hd__buf_2 _06263_ (.A(_02412_),
    .X(_02413_));
 sky130_fd_sc_hd__clkbuf_1 _06264_ (.A(_01796_),
    .X(_02414_));
 sky130_fd_sc_hd__o22a_4 _06265_ (.A1(_02156_),
    .A2(\u_spi2wb.reg_be[2] ),
    .B1(_02157_),
    .B2(wbm_sel_i[2]),
    .X(_02415_));
 sky130_fd_sc_hd__and3_1 _06266_ (.A(_02414_),
    .B(_02171_),
    .C(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__clkbuf_1 _06267_ (.A(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__a21oi_2 _06268_ (.A1(_02171_),
    .A2(_02415_),
    .B1(_01107_),
    .Y(_02418_));
 sky130_fd_sc_hd__clkbuf_1 _06269_ (.A(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__clkbuf_2 _06270_ (.A(_01106_),
    .X(_02420_));
 sky130_fd_sc_hd__clkbuf_1 _06271_ (.A(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__and2_1 _06272_ (.A(_02421_),
    .B(strap_sticky[0]),
    .X(_02422_));
 sky130_fd_sc_hd__a221o_1 _06273_ (.A1(_02413_),
    .A2(_02417_),
    .B1(_02419_),
    .B2(\u_reg.cfg_clk_ctrl[0] ),
    .C1(_02422_),
    .X(_00211_));
 sky130_fd_sc_hd__clkbuf_1 _06274_ (.A(_02340_),
    .X(_02423_));
 sky130_fd_sc_hd__buf_2 _06275_ (.A(_02423_),
    .X(_02424_));
 sky130_fd_sc_hd__and2_1 _06276_ (.A(_02421_),
    .B(strap_sticky[1]),
    .X(_02425_));
 sky130_fd_sc_hd__a221o_1 _06277_ (.A1(_02424_),
    .A2(_02417_),
    .B1(_02419_),
    .B2(\u_reg.cfg_clk_ctrl[1] ),
    .C1(_02425_),
    .X(_00212_));
 sky130_fd_sc_hd__clkbuf_1 _06278_ (.A(_02345_),
    .X(_02426_));
 sky130_fd_sc_hd__buf_2 _06279_ (.A(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__and2_1 _06280_ (.A(_02421_),
    .B(strap_sticky[2]),
    .X(_02428_));
 sky130_fd_sc_hd__a221o_1 _06281_ (.A1(_02427_),
    .A2(_02417_),
    .B1(_02419_),
    .B2(_01516_),
    .C1(_02428_),
    .X(_00213_));
 sky130_fd_sc_hd__clkbuf_1 _06282_ (.A(_02351_),
    .X(_02429_));
 sky130_fd_sc_hd__clkbuf_2 _06283_ (.A(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__and2_1 _06284_ (.A(_02421_),
    .B(strap_sticky[3]),
    .X(_02431_));
 sky130_fd_sc_hd__a221o_1 _06285_ (.A1(_02430_),
    .A2(_02417_),
    .B1(_02419_),
    .B2(_01513_),
    .C1(_02431_),
    .X(_00214_));
 sky130_fd_sc_hd__clkbuf_1 _06286_ (.A(_02355_),
    .X(_02432_));
 sky130_fd_sc_hd__clkbuf_2 _06287_ (.A(_02432_),
    .X(_02433_));
 sky130_fd_sc_hd__clkbuf_1 _06288_ (.A(_02416_),
    .X(_02434_));
 sky130_fd_sc_hd__clkbuf_1 _06289_ (.A(_02418_),
    .X(_02435_));
 sky130_fd_sc_hd__clkbuf_1 _06290_ (.A(_02420_),
    .X(_02436_));
 sky130_fd_sc_hd__and2_1 _06291_ (.A(_02436_),
    .B(strap_sticky[4]),
    .X(_02437_));
 sky130_fd_sc_hd__a221o_1 _06292_ (.A1(_02433_),
    .A2(_02434_),
    .B1(_02435_),
    .B2(\u_reg.cfg_clk_ctrl[4] ),
    .C1(_02437_),
    .X(_00215_));
 sky130_fd_sc_hd__clkbuf_1 _06293_ (.A(_02360_),
    .X(_02438_));
 sky130_fd_sc_hd__clkbuf_2 _06294_ (.A(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__and2_1 _06295_ (.A(_02436_),
    .B(strap_sticky[5]),
    .X(_02440_));
 sky130_fd_sc_hd__a221o_1 _06296_ (.A1(_02439_),
    .A2(_02434_),
    .B1(_02435_),
    .B2(\u_reg.cfg_clk_ctrl[5] ),
    .C1(_02440_),
    .X(_00216_));
 sky130_fd_sc_hd__clkbuf_1 _06297_ (.A(_02364_),
    .X(_02441_));
 sky130_fd_sc_hd__clkbuf_2 _06298_ (.A(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__and2_1 _06299_ (.A(_02436_),
    .B(strap_sticky[6]),
    .X(_02443_));
 sky130_fd_sc_hd__a221o_1 _06300_ (.A1(_02442_),
    .A2(_02434_),
    .B1(_02435_),
    .B2(\u_reg.cfg_clk_ctrl[6] ),
    .C1(_02443_),
    .X(_00217_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06301_ (.A(_02369_),
    .X(_02444_));
 sky130_fd_sc_hd__clkbuf_2 _06302_ (.A(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__and2_1 _06303_ (.A(_02436_),
    .B(strap_sticky[7]),
    .X(_02446_));
 sky130_fd_sc_hd__a221o_1 _06304_ (.A1(_02445_),
    .A2(_02434_),
    .B1(_02435_),
    .B2(\u_reg.cfg_clk_ctrl[7] ),
    .C1(_02446_),
    .X(_00218_));
 sky130_fd_sc_hd__and3b_2 _06305_ (.A_N(_02167_),
    .B(_02164_),
    .C(_02161_),
    .X(_02447_));
 sky130_fd_sc_hd__and3_1 _06306_ (.A(_02219_),
    .B(_01485_),
    .C(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06307_ (.A(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__clkbuf_2 _06308_ (.A(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _06309_ (.A0(net33),
    .A1(net225),
    .S(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__or2_1 _06310_ (.A(net66),
    .B(_02451_),
    .X(_02452_));
 sky130_fd_sc_hd__clkbuf_1 _06311_ (.A(_02452_),
    .X(_00219_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06312_ (.A(_02159_),
    .X(_02453_));
 sky130_fd_sc_hd__or3b_1 _06313_ (.A(_01479_),
    .B(_02453_),
    .C_N(_02447_),
    .X(_02454_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06314_ (.A(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__clkbuf_1 _06315_ (.A(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06316_ (.A(_02449_),
    .X(_02457_));
 sky130_fd_sc_hd__clkbuf_1 _06317_ (.A(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__or2_1 _06318_ (.A(net44),
    .B(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06319_ (.A(_01798_),
    .X(_02460_));
 sky130_fd_sc_hd__clkbuf_1 _06320_ (.A(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__o211a_1 _06321_ (.A1(_02266_),
    .A2(_02456_),
    .B1(_02459_),
    .C1(_02461_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _06322_ (.A0(net55),
    .A1(net215),
    .S(_02450_),
    .X(_02462_));
 sky130_fd_sc_hd__or2_1 _06323_ (.A(net66),
    .B(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__clkbuf_1 _06324_ (.A(_02463_),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _06325_ (.A0(net58),
    .A1(net216),
    .S(_02450_),
    .X(_02464_));
 sky130_fd_sc_hd__or2_1 _06326_ (.A(net66),
    .B(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__clkbuf_1 _06327_ (.A(_02465_),
    .X(_00222_));
 sky130_fd_sc_hd__clkbuf_2 _06328_ (.A(_02420_),
    .X(_02466_));
 sky130_fd_sc_hd__clkbuf_1 _06329_ (.A(_02466_),
    .X(_02467_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06330_ (.A(_02449_),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _06331_ (.A0(net59),
    .A1(net227),
    .S(_02468_),
    .X(_02469_));
 sky130_fd_sc_hd__or2_1 _06332_ (.A(_02467_),
    .B(_02469_),
    .X(_02470_));
 sky130_fd_sc_hd__clkbuf_1 _06333_ (.A(_02470_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _06334_ (.A0(net60),
    .A1(_02238_),
    .S(_02468_),
    .X(_02471_));
 sky130_fd_sc_hd__or2_1 _06335_ (.A(_02467_),
    .B(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__clkbuf_1 _06336_ (.A(_02472_),
    .X(_00224_));
 sky130_fd_sc_hd__clkbuf_2 _06337_ (.A(net217),
    .X(_02473_));
 sky130_fd_sc_hd__or2_1 _06338_ (.A(net61),
    .B(_02458_),
    .X(_02474_));
 sky130_fd_sc_hd__o211a_1 _06339_ (.A1(_02473_),
    .A2(_02456_),
    .B1(_02474_),
    .C1(_02461_),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _06340_ (.A0(net62),
    .A1(net218),
    .S(_02468_),
    .X(_02475_));
 sky130_fd_sc_hd__or2_1 _06341_ (.A(_02467_),
    .B(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__clkbuf_1 _06342_ (.A(_02476_),
    .X(_00226_));
 sky130_fd_sc_hd__clkbuf_2 _06343_ (.A(net224),
    .X(_02477_));
 sky130_fd_sc_hd__or2_1 _06344_ (.A(net63),
    .B(_02458_),
    .X(_02478_));
 sky130_fd_sc_hd__o211a_1 _06345_ (.A1(_02477_),
    .A2(_02456_),
    .B1(_02478_),
    .C1(_02461_),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _06346_ (.A0(net64),
    .A1(net223),
    .S(_02468_),
    .X(_02479_));
 sky130_fd_sc_hd__or2_1 _06347_ (.A(_02467_),
    .B(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__clkbuf_1 _06348_ (.A(_02480_),
    .X(_00228_));
 sky130_fd_sc_hd__clkbuf_1 _06349_ (.A(_01107_),
    .X(_02481_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06350_ (.A(_02449_),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _06351_ (.A0(net34),
    .A1(net222),
    .S(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__or2_1 _06352_ (.A(_02481_),
    .B(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__clkbuf_1 _06353_ (.A(_02484_),
    .X(_00229_));
 sky130_fd_sc_hd__clkbuf_2 _06354_ (.A(net221),
    .X(_02485_));
 sky130_fd_sc_hd__or2_1 _06355_ (.A(net35),
    .B(_02458_),
    .X(_02486_));
 sky130_fd_sc_hd__o211a_1 _06356_ (.A1(_02485_),
    .A2(_02456_),
    .B1(_02486_),
    .C1(_02461_),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _06357_ (.A0(net36),
    .A1(net220),
    .S(_02482_),
    .X(_02487_));
 sky130_fd_sc_hd__or2_1 _06358_ (.A(_02481_),
    .B(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__clkbuf_1 _06359_ (.A(_02488_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _06360_ (.A0(net37),
    .A1(_02205_),
    .S(_02482_),
    .X(_02489_));
 sky130_fd_sc_hd__or2_1 _06361_ (.A(_02481_),
    .B(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__clkbuf_1 _06362_ (.A(_02490_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _06363_ (.A0(net38),
    .A1(net219),
    .S(_02482_),
    .X(_02491_));
 sky130_fd_sc_hd__or2_1 _06364_ (.A(_02481_),
    .B(_02491_),
    .X(_02492_));
 sky130_fd_sc_hd__clkbuf_1 _06365_ (.A(_02492_),
    .X(_00233_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06366_ (.A(_02215_),
    .X(_02493_));
 sky130_fd_sc_hd__clkbuf_1 _06367_ (.A(_02455_),
    .X(_02494_));
 sky130_fd_sc_hd__clkbuf_1 _06368_ (.A(_02457_),
    .X(_02495_));
 sky130_fd_sc_hd__or2_1 _06369_ (.A(net39),
    .B(_02495_),
    .X(_02496_));
 sky130_fd_sc_hd__clkbuf_1 _06370_ (.A(_02460_),
    .X(_02497_));
 sky130_fd_sc_hd__o211a_1 _06371_ (.A1(_02493_),
    .A2(_02494_),
    .B1(_02496_),
    .C1(_02497_),
    .X(_00234_));
 sky130_fd_sc_hd__or2_1 _06372_ (.A(net40),
    .B(_02495_),
    .X(_02498_));
 sky130_fd_sc_hd__o211a_1 _06373_ (.A1(_02413_),
    .A2(_02494_),
    .B1(_02498_),
    .C1(_02497_),
    .X(_00235_));
 sky130_fd_sc_hd__or2_1 _06374_ (.A(net41),
    .B(_02495_),
    .X(_02499_));
 sky130_fd_sc_hd__o211a_1 _06375_ (.A1(_02424_),
    .A2(_02494_),
    .B1(_02499_),
    .C1(_02497_),
    .X(_00236_));
 sky130_fd_sc_hd__or2_1 _06376_ (.A(net42),
    .B(_02495_),
    .X(_02500_));
 sky130_fd_sc_hd__o211a_1 _06377_ (.A1(_02427_),
    .A2(_02494_),
    .B1(_02500_),
    .C1(_02497_),
    .X(_00237_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06378_ (.A(_01107_),
    .X(_02501_));
 sky130_fd_sc_hd__clkbuf_2 _06379_ (.A(_02448_),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _06380_ (.A0(net43),
    .A1(_02429_),
    .S(_02502_),
    .X(_02503_));
 sky130_fd_sc_hd__or2_1 _06381_ (.A(_02501_),
    .B(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__clkbuf_1 _06382_ (.A(_02504_),
    .X(_00238_));
 sky130_fd_sc_hd__clkbuf_1 _06383_ (.A(_02455_),
    .X(_02505_));
 sky130_fd_sc_hd__clkbuf_1 _06384_ (.A(_02457_),
    .X(_02506_));
 sky130_fd_sc_hd__or2_1 _06385_ (.A(net45),
    .B(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__clkbuf_1 _06386_ (.A(_02460_),
    .X(_02508_));
 sky130_fd_sc_hd__o211a_1 _06387_ (.A1(_02433_),
    .A2(_02505_),
    .B1(_02507_),
    .C1(_02508_),
    .X(_00239_));
 sky130_fd_sc_hd__or2_1 _06388_ (.A(net46),
    .B(_02506_),
    .X(_02509_));
 sky130_fd_sc_hd__o211a_1 _06389_ (.A1(_02439_),
    .A2(_02505_),
    .B1(_02509_),
    .C1(_02508_),
    .X(_00240_));
 sky130_fd_sc_hd__or2_1 _06390_ (.A(net47),
    .B(_02506_),
    .X(_02510_));
 sky130_fd_sc_hd__o211a_1 _06391_ (.A1(_02442_),
    .A2(_02505_),
    .B1(_02510_),
    .C1(_02508_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _06392_ (.A0(net48),
    .A1(_02444_),
    .S(_02502_),
    .X(_02511_));
 sky130_fd_sc_hd__or2_1 _06393_ (.A(_02501_),
    .B(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__clkbuf_1 _06394_ (.A(_02512_),
    .X(_00242_));
 sky130_fd_sc_hd__clkbuf_2 _06395_ (.A(_02374_),
    .X(_02513_));
 sky130_fd_sc_hd__or2_1 _06396_ (.A(net49),
    .B(_02506_),
    .X(_02514_));
 sky130_fd_sc_hd__o211a_1 _06397_ (.A1(_02513_),
    .A2(_02505_),
    .B1(_02514_),
    .C1(_02508_),
    .X(_00243_));
 sky130_fd_sc_hd__clkbuf_2 _06398_ (.A(_02380_),
    .X(_02515_));
 sky130_fd_sc_hd__clkbuf_1 _06399_ (.A(_02454_),
    .X(_02516_));
 sky130_fd_sc_hd__clkbuf_1 _06400_ (.A(_02450_),
    .X(_02517_));
 sky130_fd_sc_hd__or2_1 _06401_ (.A(net50),
    .B(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06402_ (.A(_02414_),
    .X(_02519_));
 sky130_fd_sc_hd__clkbuf_1 _06403_ (.A(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__o211a_1 _06404_ (.A1(_02515_),
    .A2(_02516_),
    .B1(_02518_),
    .C1(_02520_),
    .X(_00244_));
 sky130_fd_sc_hd__clkbuf_2 _06405_ (.A(_02385_),
    .X(_02521_));
 sky130_fd_sc_hd__or2_1 _06406_ (.A(net51),
    .B(_02517_),
    .X(_02522_));
 sky130_fd_sc_hd__o211a_1 _06407_ (.A1(_02521_),
    .A2(_02516_),
    .B1(_02522_),
    .C1(_02520_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _06408_ (.A0(net52),
    .A1(_02390_),
    .S(_02502_),
    .X(_02523_));
 sky130_fd_sc_hd__or2_1 _06409_ (.A(_02501_),
    .B(_02523_),
    .X(_02524_));
 sky130_fd_sc_hd__clkbuf_1 _06410_ (.A(_02524_),
    .X(_00246_));
 sky130_fd_sc_hd__clkbuf_2 _06411_ (.A(_02394_),
    .X(_02525_));
 sky130_fd_sc_hd__or2_1 _06412_ (.A(net53),
    .B(_02517_),
    .X(_02526_));
 sky130_fd_sc_hd__o211a_1 _06413_ (.A1(_02525_),
    .A2(_02516_),
    .B1(_02526_),
    .C1(_02520_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _06414_ (.A0(net54),
    .A1(_02399_),
    .S(_02502_),
    .X(_02527_));
 sky130_fd_sc_hd__or2_1 _06415_ (.A(_02501_),
    .B(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__clkbuf_1 _06416_ (.A(_02528_),
    .X(_00248_));
 sky130_fd_sc_hd__buf_2 _06417_ (.A(_02403_),
    .X(_02529_));
 sky130_fd_sc_hd__or2_1 _06418_ (.A(net56),
    .B(_02517_),
    .X(_02530_));
 sky130_fd_sc_hd__o211a_1 _06419_ (.A1(_02529_),
    .A2(_02516_),
    .B1(_02530_),
    .C1(_02520_),
    .X(_00249_));
 sky130_fd_sc_hd__clkbuf_2 _06420_ (.A(_02407_),
    .X(_02531_));
 sky130_fd_sc_hd__or2_1 _06421_ (.A(net57),
    .B(_02457_),
    .X(_02532_));
 sky130_fd_sc_hd__o211a_1 _06422_ (.A1(_02531_),
    .A2(_02455_),
    .B1(_02532_),
    .C1(_01799_),
    .X(_00250_));
 sky130_fd_sc_hd__and2_1 _06423_ (.A(_00020_),
    .B(_02453_),
    .X(_02533_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06424_ (.A(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06425_ (.A(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__clkbuf_1 _06426_ (.A(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06427_ (.A(_02288_),
    .X(_02537_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06428_ (.A(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__clkbuf_1 _06429_ (.A(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__nand2_1 _06430_ (.A(_00020_),
    .B(_02453_),
    .Y(_02540_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06431_ (.A(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06432_ (.A(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__clkbuf_2 _06433_ (.A(_02169_),
    .X(_02543_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06434_ (.A(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__nor3b_4 _06435_ (.A(_02162_),
    .B(_02168_),
    .C_N(_02165_),
    .Y(_02545_));
 sky130_fd_sc_hd__clkbuf_1 _06436_ (.A(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__clkbuf_2 _06437_ (.A(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06438_ (.A(_02220_),
    .X(_02548_));
 sky130_fd_sc_hd__clkbuf_2 _06439_ (.A(_02447_),
    .X(_02549_));
 sky130_fd_sc_hd__a22o_1 _06440_ (.A1(\u_reg.u_bank_sel.gen_bit_reg[0].u_bit_reg.data_out ),
    .A2(_02548_),
    .B1(_02549_),
    .B2(net33),
    .X(_02550_));
 sky130_fd_sc_hd__a221o_2 _06441_ (.A1(\u_reg.cfg_glb_ctrl[0] ),
    .A2(_02544_),
    .B1(_02547_),
    .B2(net1),
    .C1(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__a211o_1 _06442_ (.A1(net73),
    .A2(_02539_),
    .B1(_02542_),
    .C1(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__o21a_1 _06443_ (.A1(\u_reg.reg_rdata[0] ),
    .A2(_02536_),
    .B1(_02552_),
    .X(_00251_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06444_ (.A(_02537_),
    .X(_02553_));
 sky130_fd_sc_hd__clkbuf_1 _06445_ (.A(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__clkbuf_1 _06446_ (.A(_02540_),
    .X(_02555_));
 sky130_fd_sc_hd__a21o_1 _06447_ (.A1(net84),
    .A2(_02554_),
    .B1(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__clkbuf_2 _06448_ (.A(_02169_),
    .X(_02557_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06449_ (.A(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_1 _06450_ (.A(_02447_),
    .X(_02559_));
 sky130_fd_sc_hd__clkbuf_1 _06451_ (.A(_02559_),
    .X(_02560_));
 sky130_fd_sc_hd__a22o_1 _06452_ (.A1(\u_reg.cfg_glb_ctrl[1] ),
    .A2(_02558_),
    .B1(_02560_),
    .B2(net44),
    .X(_02561_));
 sky130_fd_sc_hd__clkbuf_1 _06453_ (.A(_02548_),
    .X(_02562_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06454_ (.A(_02547_),
    .X(_02563_));
 sky130_fd_sc_hd__a22o_1 _06455_ (.A1(\u_reg.u_bank_sel.gen_bit_reg[1].u_bit_reg.data_out ),
    .A2(_02562_),
    .B1(_02563_),
    .B2(net12),
    .X(_02564_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06456_ (.A(_02534_),
    .X(_02565_));
 sky130_fd_sc_hd__clkbuf_1 _06457_ (.A(_02565_),
    .X(_02566_));
 sky130_fd_sc_hd__o32a_1 _06458_ (.A1(_02556_),
    .A2(_02561_),
    .A3(_02564_),
    .B1(_02566_),
    .B2(\u_reg.reg_rdata[1] ),
    .X(_00252_));
 sky130_fd_sc_hd__clkbuf_1 _06459_ (.A(_02544_),
    .X(_02567_));
 sky130_fd_sc_hd__clkbuf_1 _06460_ (.A(_02548_),
    .X(_02568_));
 sky130_fd_sc_hd__clkbuf_2 _06461_ (.A(_02549_),
    .X(_02569_));
 sky130_fd_sc_hd__a22o_1 _06462_ (.A1(\u_reg.u_bank_sel.gen_bit_reg[2].u_bit_reg.data_out ),
    .A2(_02568_),
    .B1(_02569_),
    .B2(net55),
    .X(_02570_));
 sky130_fd_sc_hd__a221o_2 _06463_ (.A1(\u_reg.cfg_glb_ctrl[2] ),
    .A2(_02567_),
    .B1(_02563_),
    .B2(net23),
    .C1(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__clkbuf_1 _06464_ (.A(_02538_),
    .X(_02572_));
 sky130_fd_sc_hd__clkbuf_1 _06465_ (.A(_02541_),
    .X(_02573_));
 sky130_fd_sc_hd__a21o_1 _06466_ (.A1(net95),
    .A2(_02572_),
    .B1(_02573_),
    .X(_02574_));
 sky130_fd_sc_hd__o22a_1 _06467_ (.A1(\u_reg.reg_rdata[2] ),
    .A2(_02536_),
    .B1(_02571_),
    .B2(_02574_),
    .X(_00253_));
 sky130_fd_sc_hd__a21o_1 _06468_ (.A1(net98),
    .A2(_02554_),
    .B1(_02555_),
    .X(_02575_));
 sky130_fd_sc_hd__a22o_1 _06469_ (.A1(\u_reg.cfg_glb_ctrl[3] ),
    .A2(_02558_),
    .B1(_02560_),
    .B2(net58),
    .X(_02576_));
 sky130_fd_sc_hd__a22o_1 _06470_ (.A1(\u_async_wb.m_cmd_wr_data[56] ),
    .A2(_02562_),
    .B1(_02563_),
    .B2(net26),
    .X(_02577_));
 sky130_fd_sc_hd__o32a_1 _06471_ (.A1(_02575_),
    .A2(_02576_),
    .A3(_02577_),
    .B1(_02566_),
    .B2(\u_reg.reg_rdata[3] ),
    .X(_00254_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06472_ (.A(_02547_),
    .X(_02578_));
 sky130_fd_sc_hd__a22o_1 _06473_ (.A1(\u_async_wb.m_cmd_wr_data[57] ),
    .A2(_02568_),
    .B1(_02569_),
    .B2(net59),
    .X(_02579_));
 sky130_fd_sc_hd__a221o_2 _06474_ (.A1(\u_reg.cfg_glb_ctrl[4] ),
    .A2(_02567_),
    .B1(_02578_),
    .B2(net27),
    .C1(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__a21o_1 _06475_ (.A1(net99),
    .A2(_02572_),
    .B1(_02573_),
    .X(_02581_));
 sky130_fd_sc_hd__o22a_1 _06476_ (.A1(\u_reg.reg_rdata[4] ),
    .A2(_02536_),
    .B1(_02580_),
    .B2(_02581_),
    .X(_00255_));
 sky130_fd_sc_hd__a22o_1 _06477_ (.A1(\u_async_wb.m_cmd_wr_data[58] ),
    .A2(_02568_),
    .B1(_02569_),
    .B2(net60),
    .X(_02582_));
 sky130_fd_sc_hd__a221o_2 _06478_ (.A1(\u_reg.cfg_glb_ctrl[5] ),
    .A2(_02567_),
    .B1(_02578_),
    .B2(net28),
    .C1(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__a21o_1 _06479_ (.A1(net100),
    .A2(_02572_),
    .B1(_02573_),
    .X(_02584_));
 sky130_fd_sc_hd__o22a_1 _06480_ (.A1(\u_reg.reg_rdata[5] ),
    .A2(_02536_),
    .B1(_02583_),
    .B2(_02584_),
    .X(_00256_));
 sky130_fd_sc_hd__a21o_1 _06481_ (.A1(net101),
    .A2(_02554_),
    .B1(_02555_),
    .X(_02585_));
 sky130_fd_sc_hd__clkbuf_2 _06482_ (.A(_02546_),
    .X(_02586_));
 sky130_fd_sc_hd__clkbuf_1 _06483_ (.A(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__a22o_1 _06484_ (.A1(\u_reg.cfg_glb_ctrl[6] ),
    .A2(_02558_),
    .B1(_02587_),
    .B2(net29),
    .X(_02588_));
 sky130_fd_sc_hd__a22o_1 _06485_ (.A1(\u_async_wb.m_cmd_wr_data[59] ),
    .A2(_02562_),
    .B1(_02560_),
    .B2(net61),
    .X(_02589_));
 sky130_fd_sc_hd__o32a_1 _06486_ (.A1(_02585_),
    .A2(_02588_),
    .A3(_02589_),
    .B1(_02566_),
    .B2(\u_reg.reg_rdata[6] ),
    .X(_00257_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06487_ (.A(_02535_),
    .X(_02590_));
 sky130_fd_sc_hd__a22o_1 _06488_ (.A1(\u_async_wb.m_cmd_wr_data[60] ),
    .A2(_02568_),
    .B1(_02559_),
    .B2(net62),
    .X(_02591_));
 sky130_fd_sc_hd__a221o_2 _06489_ (.A1(\u_reg.cfg_glb_ctrl[7] ),
    .A2(_02558_),
    .B1(_02578_),
    .B2(net30),
    .C1(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__a21o_1 _06490_ (.A1(net102),
    .A2(_02572_),
    .B1(_02573_),
    .X(_02593_));
 sky130_fd_sc_hd__o22a_1 _06491_ (.A1(\u_reg.reg_rdata[7] ),
    .A2(_02590_),
    .B1(_02592_),
    .B2(_02593_),
    .X(_00258_));
 sky130_fd_sc_hd__a21o_1 _06492_ (.A1(net103),
    .A2(_02554_),
    .B1(_02555_),
    .X(_02594_));
 sky130_fd_sc_hd__clkbuf_1 _06493_ (.A(_02559_),
    .X(_02595_));
 sky130_fd_sc_hd__a22o_1 _06494_ (.A1(net63),
    .A2(_02595_),
    .B1(_02587_),
    .B2(net31),
    .X(_02596_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06495_ (.A(_02544_),
    .X(_02597_));
 sky130_fd_sc_hd__clkbuf_1 _06496_ (.A(_02548_),
    .X(_02598_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06497_ (.A(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__a22o_1 _06498_ (.A1(\u_reg.cfg_glb_ctrl[8] ),
    .A2(_02597_),
    .B1(_02599_),
    .B2(\u_async_wb.m_cmd_wr_data[61] ),
    .X(_02600_));
 sky130_fd_sc_hd__o32a_1 _06499_ (.A1(_02594_),
    .A2(_02596_),
    .A3(_02600_),
    .B1(_02566_),
    .B2(\u_reg.reg_rdata[8] ),
    .X(_00259_));
 sky130_fd_sc_hd__a22o_1 _06500_ (.A1(\u_reg.cfg_glb_ctrl[9] ),
    .A2(_02544_),
    .B1(_02598_),
    .B2(\u_async_wb.m_cmd_wr_data[62] ),
    .X(_02601_));
 sky130_fd_sc_hd__a221o_2 _06501_ (.A1(net64),
    .A2(_02595_),
    .B1(_02578_),
    .B2(net32),
    .C1(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06502_ (.A(_02541_),
    .X(_02603_));
 sky130_fd_sc_hd__a21o_1 _06503_ (.A1(net104),
    .A2(_02539_),
    .B1(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__o22a_1 _06504_ (.A1(\u_reg.reg_rdata[9] ),
    .A2(_02590_),
    .B1(_02602_),
    .B2(_02604_),
    .X(_00260_));
 sky130_fd_sc_hd__a22o_1 _06505_ (.A1(\u_reg.cfg_glb_ctrl[10] ),
    .A2(_02557_),
    .B1(_02598_),
    .B2(\u_async_wb.m_cmd_wr_data[63] ),
    .X(_02605_));
 sky130_fd_sc_hd__a221o_2 _06506_ (.A1(net34),
    .A2(_02595_),
    .B1(_02587_),
    .B2(net2),
    .C1(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__a21o_1 _06507_ (.A1(net74),
    .A2(_02539_),
    .B1(_02603_),
    .X(_02607_));
 sky130_fd_sc_hd__o22a_1 _06508_ (.A1(\u_reg.reg_rdata[10] ),
    .A2(_02590_),
    .B1(_02606_),
    .B2(_02607_),
    .X(_00261_));
 sky130_fd_sc_hd__clkbuf_1 _06509_ (.A(_02553_),
    .X(_02608_));
 sky130_fd_sc_hd__clkbuf_1 _06510_ (.A(_02540_),
    .X(_02609_));
 sky130_fd_sc_hd__a21o_1 _06511_ (.A1(net75),
    .A2(_02608_),
    .B1(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__clkbuf_2 _06512_ (.A(_02559_),
    .X(_02611_));
 sky130_fd_sc_hd__clkbuf_2 _06513_ (.A(_02586_),
    .X(_02612_));
 sky130_fd_sc_hd__a22o_1 _06514_ (.A1(net35),
    .A2(_02611_),
    .B1(_02612_),
    .B2(net3),
    .X(_02613_));
 sky130_fd_sc_hd__a22o_1 _06515_ (.A1(\u_reg.cfg_glb_ctrl[11] ),
    .A2(_02597_),
    .B1(_02599_),
    .B2(\u_async_wb.m_cmd_wr_data[64] ),
    .X(_02614_));
 sky130_fd_sc_hd__clkbuf_1 _06516_ (.A(_02565_),
    .X(_02615_));
 sky130_fd_sc_hd__o32a_1 _06517_ (.A1(_02610_),
    .A2(_02613_),
    .A3(_02614_),
    .B1(_02615_),
    .B2(\u_reg.reg_rdata[11] ),
    .X(_00262_));
 sky130_fd_sc_hd__a21o_1 _06518_ (.A1(net76),
    .A2(_02608_),
    .B1(_02609_),
    .X(_02616_));
 sky130_fd_sc_hd__a22o_1 _06519_ (.A1(\u_async_wb.m_cmd_wr_data[65] ),
    .A2(_02562_),
    .B1(_02560_),
    .B2(net36),
    .X(_02617_));
 sky130_fd_sc_hd__a22o_1 _06520_ (.A1(\u_reg.cfg_glb_ctrl[12] ),
    .A2(_02597_),
    .B1(_02563_),
    .B2(net4),
    .X(_02618_));
 sky130_fd_sc_hd__o32a_1 _06521_ (.A1(_02616_),
    .A2(_02617_),
    .A3(_02618_),
    .B1(_02615_),
    .B2(\u_reg.reg_rdata[12] ),
    .X(_00263_));
 sky130_fd_sc_hd__a21o_1 _06522_ (.A1(net77),
    .A2(_02608_),
    .B1(_02609_),
    .X(_02619_));
 sky130_fd_sc_hd__a22o_1 _06523_ (.A1(net37),
    .A2(_02611_),
    .B1(_02612_),
    .B2(net5),
    .X(_02620_));
 sky130_fd_sc_hd__a22o_1 _06524_ (.A1(\u_reg.cfg_glb_ctrl[13] ),
    .A2(_02597_),
    .B1(_02599_),
    .B2(\u_async_wb.m_cmd_wr_data[66] ),
    .X(_02621_));
 sky130_fd_sc_hd__o32a_1 _06525_ (.A1(_02619_),
    .A2(_02620_),
    .A3(_02621_),
    .B1(_02615_),
    .B2(\u_reg.reg_rdata[13] ),
    .X(_00264_));
 sky130_fd_sc_hd__a22o_1 _06526_ (.A1(\u_reg.cfg_glb_ctrl[14] ),
    .A2(_02557_),
    .B1(_02598_),
    .B2(\u_async_wb.m_cmd_wr_data[67] ),
    .X(_02622_));
 sky130_fd_sc_hd__a221o_2 _06527_ (.A1(net38),
    .A2(_02595_),
    .B1(_02587_),
    .B2(net6),
    .C1(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__a21o_1 _06528_ (.A1(net78),
    .A2(_02539_),
    .B1(_02603_),
    .X(_02624_));
 sky130_fd_sc_hd__o22a_1 _06529_ (.A1(\u_reg.reg_rdata[14] ),
    .A2(_02590_),
    .B1(_02623_),
    .B2(_02624_),
    .X(_00265_));
 sky130_fd_sc_hd__a21o_1 _06530_ (.A1(net79),
    .A2(_02608_),
    .B1(_02609_),
    .X(_02625_));
 sky130_fd_sc_hd__a22o_1 _06531_ (.A1(net39),
    .A2(_02611_),
    .B1(_02612_),
    .B2(net7),
    .X(_02626_));
 sky130_fd_sc_hd__a22o_1 _06532_ (.A1(\u_reg.cfg_glb_ctrl[15] ),
    .A2(_02567_),
    .B1(_02599_),
    .B2(\u_async_wb.m_cmd_wr_data[68] ),
    .X(_02627_));
 sky130_fd_sc_hd__o32a_1 _06533_ (.A1(_02625_),
    .A2(_02626_),
    .A3(_02627_),
    .B1(_02615_),
    .B2(\u_reg.reg_rdata[15] ),
    .X(_00266_));
 sky130_fd_sc_hd__clkbuf_1 _06534_ (.A(_02549_),
    .X(_02628_));
 sky130_fd_sc_hd__a22o_1 _06535_ (.A1(\u_reg.cfg_clk_ctrl[0] ),
    .A2(_02557_),
    .B1(_02586_),
    .B2(net8),
    .X(_02629_));
 sky130_fd_sc_hd__a221o_1 _06536_ (.A1(net80),
    .A2(_02553_),
    .B1(_02628_),
    .B2(net40),
    .C1(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _06537_ (.A0(\u_reg.reg_rdata[16] ),
    .A1(_02630_),
    .S(_02565_),
    .X(_02631_));
 sky130_fd_sc_hd__clkbuf_1 _06538_ (.A(_02631_),
    .X(_00267_));
 sky130_fd_sc_hd__clkbuf_1 _06539_ (.A(_02169_),
    .X(_02632_));
 sky130_fd_sc_hd__a22o_1 _06540_ (.A1(\u_reg.cfg_clk_ctrl[1] ),
    .A2(_02632_),
    .B1(_02586_),
    .B2(net9),
    .X(_02633_));
 sky130_fd_sc_hd__a221o_1 _06541_ (.A1(net81),
    .A2(_02553_),
    .B1(_02628_),
    .B2(net41),
    .C1(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__mux2_1 _06542_ (.A0(\u_reg.reg_rdata[17] ),
    .A1(_02634_),
    .S(_02565_),
    .X(_02635_));
 sky130_fd_sc_hd__clkbuf_1 _06543_ (.A(_02635_),
    .X(_00268_));
 sky130_fd_sc_hd__clkbuf_1 _06544_ (.A(_02288_),
    .X(_02636_));
 sky130_fd_sc_hd__clkbuf_1 _06545_ (.A(_02545_),
    .X(_02637_));
 sky130_fd_sc_hd__a22o_1 _06546_ (.A1(\u_reg.cfg_clk_ctrl[2] ),
    .A2(_02632_),
    .B1(_02637_),
    .B2(net10),
    .X(_02638_));
 sky130_fd_sc_hd__a221o_1 _06547_ (.A1(net82),
    .A2(_02636_),
    .B1(_02628_),
    .B2(net42),
    .C1(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06548_ (.A(_02533_),
    .X(_02640_));
 sky130_fd_sc_hd__mux2_1 _06549_ (.A0(\u_reg.reg_rdata[18] ),
    .A1(_02639_),
    .S(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__clkbuf_1 _06550_ (.A(_02641_),
    .X(_00269_));
 sky130_fd_sc_hd__clkbuf_1 _06551_ (.A(_02549_),
    .X(_02642_));
 sky130_fd_sc_hd__a22o_1 _06552_ (.A1(\u_reg.cfg_clk_ctrl[3] ),
    .A2(_02632_),
    .B1(_02637_),
    .B2(net11),
    .X(_02643_));
 sky130_fd_sc_hd__a221o_1 _06553_ (.A1(net83),
    .A2(_02636_),
    .B1(_02642_),
    .B2(net43),
    .C1(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__mux2_1 _06554_ (.A0(\u_reg.reg_rdata[19] ),
    .A1(_02644_),
    .S(_02640_),
    .X(_02645_));
 sky130_fd_sc_hd__clkbuf_1 _06555_ (.A(_02645_),
    .X(_00270_));
 sky130_fd_sc_hd__a22o_1 _06556_ (.A1(\u_reg.cfg_clk_ctrl[4] ),
    .A2(_02632_),
    .B1(_02637_),
    .B2(net13),
    .X(_02646_));
 sky130_fd_sc_hd__a221o_1 _06557_ (.A1(net85),
    .A2(_02636_),
    .B1(_02642_),
    .B2(net45),
    .C1(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__mux2_1 _06558_ (.A0(\u_reg.reg_rdata[20] ),
    .A1(_02647_),
    .S(_02640_),
    .X(_02648_));
 sky130_fd_sc_hd__clkbuf_1 _06559_ (.A(_02648_),
    .X(_00271_));
 sky130_fd_sc_hd__a22o_1 _06560_ (.A1(\u_reg.cfg_clk_ctrl[5] ),
    .A2(_02543_),
    .B1(_02637_),
    .B2(net14),
    .X(_02649_));
 sky130_fd_sc_hd__a221o_1 _06561_ (.A1(net86),
    .A2(_02636_),
    .B1(_02642_),
    .B2(net46),
    .C1(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__mux2_1 _06562_ (.A0(\u_reg.reg_rdata[21] ),
    .A1(_02650_),
    .S(_02640_),
    .X(_02651_));
 sky130_fd_sc_hd__clkbuf_1 _06563_ (.A(_02651_),
    .X(_00272_));
 sky130_fd_sc_hd__a22o_1 _06564_ (.A1(\u_reg.cfg_clk_ctrl[6] ),
    .A2(_02543_),
    .B1(_02546_),
    .B2(net15),
    .X(_02652_));
 sky130_fd_sc_hd__a221o_1 _06565_ (.A1(net87),
    .A2(_02537_),
    .B1(_02642_),
    .B2(net47),
    .C1(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _06566_ (.A0(\u_reg.reg_rdata[22] ),
    .A1(_02653_),
    .S(_02534_),
    .X(_02654_));
 sky130_fd_sc_hd__clkbuf_1 _06567_ (.A(_02654_),
    .X(_00273_));
 sky130_fd_sc_hd__a22o_1 _06568_ (.A1(\u_reg.cfg_clk_ctrl[7] ),
    .A2(_02543_),
    .B1(_02546_),
    .B2(net16),
    .X(_02655_));
 sky130_fd_sc_hd__a221o_1 _06569_ (.A1(net88),
    .A2(_02537_),
    .B1(_02569_),
    .B2(net48),
    .C1(_02655_),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _06570_ (.A0(\u_reg.reg_rdata[23] ),
    .A1(_02656_),
    .S(_02534_),
    .X(_02657_));
 sky130_fd_sc_hd__clkbuf_1 _06571_ (.A(_02657_),
    .X(_00274_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06572_ (.A(_02535_),
    .X(_02658_));
 sky130_fd_sc_hd__clkbuf_1 _06573_ (.A(_02538_),
    .X(_02659_));
 sky130_fd_sc_hd__clkbuf_1 _06574_ (.A(_02612_),
    .X(_02660_));
 sky130_fd_sc_hd__a22o_1 _06575_ (.A1(net89),
    .A2(_02659_),
    .B1(_02660_),
    .B2(net17),
    .X(_02661_));
 sky130_fd_sc_hd__clkbuf_1 _06576_ (.A(_02611_),
    .X(_02662_));
 sky130_fd_sc_hd__a21o_1 _06577_ (.A1(net49),
    .A2(_02662_),
    .B1(_02603_),
    .X(_02663_));
 sky130_fd_sc_hd__o22a_1 _06578_ (.A1(\u_reg.reg_rdata[24] ),
    .A2(_02658_),
    .B1(_02661_),
    .B2(_02663_),
    .X(_00275_));
 sky130_fd_sc_hd__a21o_1 _06579_ (.A1(net90),
    .A2(_02659_),
    .B1(_02542_),
    .X(_02664_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06580_ (.A(_02628_),
    .X(_02665_));
 sky130_fd_sc_hd__a22o_1 _06581_ (.A1(net50),
    .A2(_02665_),
    .B1(_02660_),
    .B2(net18),
    .X(_02666_));
 sky130_fd_sc_hd__o22a_1 _06582_ (.A1(\u_reg.reg_rdata[25] ),
    .A2(_02658_),
    .B1(_02664_),
    .B2(_02666_),
    .X(_00276_));
 sky130_fd_sc_hd__a22o_1 _06583_ (.A1(net91),
    .A2(_02659_),
    .B1(_02660_),
    .B2(net19),
    .X(_02667_));
 sky130_fd_sc_hd__clkbuf_1 _06584_ (.A(_02541_),
    .X(_02668_));
 sky130_fd_sc_hd__a21o_1 _06585_ (.A1(net51),
    .A2(_02662_),
    .B1(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__o22a_1 _06586_ (.A1(\u_reg.reg_rdata[26] ),
    .A2(_02658_),
    .B1(_02667_),
    .B2(_02669_),
    .X(_00277_));
 sky130_fd_sc_hd__clkbuf_1 _06587_ (.A(_02538_),
    .X(_02670_));
 sky130_fd_sc_hd__clkbuf_1 _06588_ (.A(_02547_),
    .X(_02671_));
 sky130_fd_sc_hd__a22o_1 _06589_ (.A1(net92),
    .A2(_02670_),
    .B1(_02671_),
    .B2(net20),
    .X(_02672_));
 sky130_fd_sc_hd__a21o_1 _06590_ (.A1(net52),
    .A2(_02662_),
    .B1(_02668_),
    .X(_02673_));
 sky130_fd_sc_hd__o22a_1 _06591_ (.A1(\u_reg.reg_rdata[27] ),
    .A2(_02658_),
    .B1(_02672_),
    .B2(_02673_),
    .X(_00278_));
 sky130_fd_sc_hd__clkbuf_1 _06592_ (.A(_02535_),
    .X(_02674_));
 sky130_fd_sc_hd__a21o_1 _06593_ (.A1(net21),
    .A2(_02660_),
    .B1(_02542_),
    .X(_02675_));
 sky130_fd_sc_hd__a22o_1 _06594_ (.A1(net93),
    .A2(_02659_),
    .B1(_02665_),
    .B2(net53),
    .X(_02676_));
 sky130_fd_sc_hd__o22a_1 _06595_ (.A1(\u_reg.reg_rdata[28] ),
    .A2(_02674_),
    .B1(_02675_),
    .B2(_02676_),
    .X(_00279_));
 sky130_fd_sc_hd__a22o_1 _06596_ (.A1(net94),
    .A2(_02670_),
    .B1(_02671_),
    .B2(net22),
    .X(_02677_));
 sky130_fd_sc_hd__a21o_1 _06597_ (.A1(net54),
    .A2(_02662_),
    .B1(_02668_),
    .X(_02678_));
 sky130_fd_sc_hd__o22a_1 _06598_ (.A1(\u_reg.reg_rdata[29] ),
    .A2(_02674_),
    .B1(_02677_),
    .B2(_02678_),
    .X(_00280_));
 sky130_fd_sc_hd__a22o_1 _06599_ (.A1(net96),
    .A2(_02670_),
    .B1(_02671_),
    .B2(net24),
    .X(_02679_));
 sky130_fd_sc_hd__a21o_1 _06600_ (.A1(net56),
    .A2(_02665_),
    .B1(_02668_),
    .X(_02680_));
 sky130_fd_sc_hd__o22a_1 _06601_ (.A1(\u_reg.reg_rdata[30] ),
    .A2(_02674_),
    .B1(_02679_),
    .B2(_02680_),
    .X(_00281_));
 sky130_fd_sc_hd__a22o_1 _06602_ (.A1(net97),
    .A2(_02670_),
    .B1(_02671_),
    .B2(net25),
    .X(_02681_));
 sky130_fd_sc_hd__a21o_1 _06603_ (.A1(net57),
    .A2(_02665_),
    .B1(_02542_),
    .X(_02682_));
 sky130_fd_sc_hd__o22a_1 _06604_ (.A1(\u_reg.reg_rdata[31] ),
    .A2(_02674_),
    .B1(_02681_),
    .B2(_02682_),
    .X(_00282_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06605_ (.A(_01507_),
    .X(_02683_));
 sky130_fd_sc_hd__and2b_1 _06606_ (.A_N(_02683_),
    .B(_01790_),
    .X(_02684_));
 sky130_fd_sc_hd__and2b_1 _06607_ (.A_N(_01790_),
    .B(_02683_),
    .X(_02685_));
 sky130_fd_sc_hd__nor2_1 _06608_ (.A(_02684_),
    .B(_02685_),
    .Y(_00283_));
 sky130_fd_sc_hd__inv_2 _06609_ (.A(\u_async_wb.u_resp_if.rd_ptr[1] ),
    .Y(_02686_));
 sky130_fd_sc_hd__xnor2_1 _06610_ (.A(_02686_),
    .B(_02684_),
    .Y(_00284_));
 sky130_fd_sc_hd__clkbuf_1 _06611_ (.A(_01796_),
    .X(_02687_));
 sky130_fd_sc_hd__nor2_1 _06612_ (.A(_01797_),
    .B(strap_sticky[17]),
    .Y(_02688_));
 sky130_fd_sc_hd__a22o_1 _06613_ (.A1(_02687_),
    .A2(net226),
    .B1(_02688_),
    .B2(strap_sticky[16]),
    .X(_02689_));
 sky130_fd_sc_hd__or3b_2 _06614_ (.A(_01478_),
    .B(_02159_),
    .C_N(_02545_),
    .X(_02690_));
 sky130_fd_sc_hd__nand2_1 _06615_ (.A(_02414_),
    .B(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06616_ (.A(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__mux2_1 _06617_ (.A0(net12),
    .A1(_02689_),
    .S(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__clkbuf_1 _06618_ (.A(_02693_),
    .X(_00285_));
 sky130_fd_sc_hd__and2_1 _06619_ (.A(_01796_),
    .B(_02690_),
    .X(_02694_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06620_ (.A(_02694_),
    .X(_02695_));
 sky130_fd_sc_hd__nor2_1 _06621_ (.A(_02420_),
    .B(_02690_),
    .Y(_02696_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06622_ (.A(_02696_),
    .X(_02697_));
 sky130_fd_sc_hd__a221o_1 _06623_ (.A1(net23),
    .A2(_02695_),
    .B1(_02697_),
    .B2(_02259_),
    .C1(_02688_),
    .X(_00286_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06624_ (.A(_02692_),
    .X(_02698_));
 sky130_fd_sc_hd__or2_1 _06625_ (.A(_01106_),
    .B(_02690_),
    .X(_02699_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06626_ (.A(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__or3b_1 _06627_ (.A(_02519_),
    .B(strap_sticky[16]),
    .C_N(strap_sticky[17]),
    .X(_02701_));
 sky130_fd_sc_hd__o221a_1 _06628_ (.A1(net26),
    .A2(_02698_),
    .B1(_02700_),
    .B2(_02254_),
    .C1(_02701_),
    .X(_00287_));
 sky130_fd_sc_hd__nor2_1 _06629_ (.A(_01797_),
    .B(strap_sticky[19]),
    .Y(_02702_));
 sky130_fd_sc_hd__a22o_1 _06630_ (.A1(_02687_),
    .A2(net228),
    .B1(_02702_),
    .B2(strap_sticky[18]),
    .X(_02703_));
 sky130_fd_sc_hd__mux2_1 _06631_ (.A0(net28),
    .A1(_02703_),
    .S(_02692_),
    .X(_02704_));
 sky130_fd_sc_hd__clkbuf_1 _06632_ (.A(_02704_),
    .X(_00288_));
 sky130_fd_sc_hd__a221o_1 _06633_ (.A1(net29),
    .A2(_02695_),
    .B1(_02697_),
    .B2(_02473_),
    .C1(_02702_),
    .X(_00289_));
 sky130_fd_sc_hd__or3b_1 _06634_ (.A(_02519_),
    .B(strap_sticky[18]),
    .C_N(strap_sticky[19]),
    .X(_02705_));
 sky130_fd_sc_hd__o221a_1 _06635_ (.A1(net30),
    .A2(_02698_),
    .B1(_02700_),
    .B2(_02228_),
    .C1(_02705_),
    .X(_00290_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06636_ (.A(_02694_),
    .X(_02706_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06637_ (.A(_02706_),
    .X(_02707_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06638_ (.A(_02696_),
    .X(_02708_));
 sky130_fd_sc_hd__inv_2 _06639_ (.A(strap_sticky[20]),
    .Y(_02709_));
 sky130_fd_sc_hd__or2_1 _06640_ (.A(_02687_),
    .B(strap_sticky[21]),
    .X(_02710_));
 sky130_fd_sc_hd__nor2_1 _06641_ (.A(_02709_),
    .B(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__a221o_1 _06642_ (.A1(net32),
    .A2(_02707_),
    .B1(_02708_),
    .B2(_02181_),
    .C1(_02711_),
    .X(_00291_));
 sky130_fd_sc_hd__o221a_1 _06643_ (.A1(net2),
    .A2(_02698_),
    .B1(_02700_),
    .B2(_02187_),
    .C1(_02710_),
    .X(_00292_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06644_ (.A(_02691_),
    .X(_02712_));
 sky130_fd_sc_hd__clkbuf_1 _06645_ (.A(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__clkbuf_1 _06646_ (.A(_02699_),
    .X(_02714_));
 sky130_fd_sc_hd__clkbuf_1 _06647_ (.A(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__or3b_1 _06648_ (.A(_02519_),
    .B(_02709_),
    .C_N(strap_sticky[21]),
    .X(_02716_));
 sky130_fd_sc_hd__o221a_1 _06649_ (.A1(net3),
    .A2(_02713_),
    .B1(_02715_),
    .B2(_02485_),
    .C1(_02716_),
    .X(_00293_));
 sky130_fd_sc_hd__nor2_1 _06650_ (.A(_01797_),
    .B(strap_sticky[23]),
    .Y(_02717_));
 sky130_fd_sc_hd__a22o_1 _06651_ (.A1(_02414_),
    .A2(net229),
    .B1(_02717_),
    .B2(strap_sticky[22]),
    .X(_02718_));
 sky130_fd_sc_hd__mux2_1 _06652_ (.A0(net5),
    .A1(_02718_),
    .S(_02692_),
    .X(_02719_));
 sky130_fd_sc_hd__clkbuf_1 _06653_ (.A(_02719_),
    .X(_00294_));
 sky130_fd_sc_hd__a221o_1 _06654_ (.A1(net6),
    .A2(_02707_),
    .B1(_02708_),
    .B2(_02211_),
    .C1(_02717_),
    .X(_00295_));
 sky130_fd_sc_hd__clkinv_2 _06655_ (.A(strap_sticky[22]),
    .Y(_02720_));
 sky130_fd_sc_hd__and3_1 _06656_ (.A(_02466_),
    .B(_02720_),
    .C(strap_sticky[23]),
    .X(_02721_));
 sky130_fd_sc_hd__a221o_1 _06657_ (.A1(net7),
    .A2(_02707_),
    .B1(_02708_),
    .B2(_02493_),
    .C1(_02721_),
    .X(_00296_));
 sky130_fd_sc_hd__inv_2 _06658_ (.A(strap_sticky[25]),
    .Y(_02722_));
 sky130_fd_sc_hd__a21oi_1 _06659_ (.A1(_02722_),
    .A2(strap_sticky[24]),
    .B1(_01799_),
    .Y(_02723_));
 sky130_fd_sc_hd__a221o_1 _06660_ (.A1(net9),
    .A2(_02707_),
    .B1(_02708_),
    .B2(_02424_),
    .C1(_02723_),
    .X(_00297_));
 sky130_fd_sc_hd__o21ai_1 _06661_ (.A1(strap_sticky[25]),
    .A2(strap_sticky[24]),
    .B1(_02466_),
    .Y(_02724_));
 sky130_fd_sc_hd__o221a_1 _06662_ (.A1(net10),
    .A2(_02713_),
    .B1(_02715_),
    .B2(_02427_),
    .C1(_02724_),
    .X(_00298_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06663_ (.A(_02696_),
    .X(_02725_));
 sky130_fd_sc_hd__a21oi_1 _06664_ (.A1(strap_sticky[25]),
    .A2(strap_sticky[24]),
    .B1(_02724_),
    .Y(_02726_));
 sky130_fd_sc_hd__a221o_1 _06665_ (.A1(net11),
    .A2(_02706_),
    .B1(_02725_),
    .B2(_02430_),
    .C1(_02726_),
    .X(_00299_));
 sky130_fd_sc_hd__or3b_1 _06666_ (.A(_01798_),
    .B(strap_sticky[27]),
    .C_N(strap_sticky[26]),
    .X(_02727_));
 sky130_fd_sc_hd__o221a_1 _06667_ (.A1(net14),
    .A2(_02713_),
    .B1(_02715_),
    .B2(_02439_),
    .C1(_02727_),
    .X(_00300_));
 sky130_fd_sc_hd__or3_1 _06668_ (.A(_01798_),
    .B(strap_sticky[27]),
    .C(strap_sticky[26]),
    .X(_02728_));
 sky130_fd_sc_hd__o221a_1 _06669_ (.A1(net15),
    .A2(_02713_),
    .B1(_02715_),
    .B2(_02442_),
    .C1(_02728_),
    .X(_00301_));
 sky130_fd_sc_hd__a21o_1 _06670_ (.A1(strap_sticky[27]),
    .A2(strap_sticky[26]),
    .B1(_02460_),
    .X(_02729_));
 sky130_fd_sc_hd__o221a_1 _06671_ (.A1(net16),
    .A2(_02712_),
    .B1(_02714_),
    .B2(_02445_),
    .C1(_02729_),
    .X(_00302_));
 sky130_fd_sc_hd__inv_2 _06672_ (.A(strap_sticky[28]),
    .Y(_02730_));
 sky130_fd_sc_hd__or2_1 _06673_ (.A(_02687_),
    .B(strap_sticky[29]),
    .X(_02731_));
 sky130_fd_sc_hd__nor2_1 _06674_ (.A(_02730_),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__a221o_1 _06675_ (.A1(net18),
    .A2(_02706_),
    .B1(_02725_),
    .B2(_02515_),
    .C1(_02732_),
    .X(_00303_));
 sky130_fd_sc_hd__o221a_1 _06676_ (.A1(net19),
    .A2(_02712_),
    .B1(_02714_),
    .B2(_02521_),
    .C1(_02731_),
    .X(_00304_));
 sky130_fd_sc_hd__clkbuf_2 _06677_ (.A(_02390_),
    .X(_02733_));
 sky130_fd_sc_hd__and3_1 _06678_ (.A(_02466_),
    .B(strap_sticky[28]),
    .C(strap_sticky[29]),
    .X(_02734_));
 sky130_fd_sc_hd__a221o_1 _06679_ (.A1(net20),
    .A2(_02706_),
    .B1(_02725_),
    .B2(_02733_),
    .C1(_02734_),
    .X(_00305_));
 sky130_fd_sc_hd__inv_2 _06680_ (.A(\u_async_wb.u_resp_if.wr_ptr[0] ),
    .Y(_02735_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06681_ (.A(\u_async_wb.u_resp_if.wr_ptr[1] ),
    .X(_02736_));
 sky130_fd_sc_hd__inv_2 _06682_ (.A(\u_async_wb.u_resp_if.sync_rd_ptr_1[1] ),
    .Y(_02737_));
 sky130_fd_sc_hd__xnor2_1 _06683_ (.A(\u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(\u_async_wb.u_resp_if.sync_rd_ptr_1[0] ),
    .Y(_02738_));
 sky130_fd_sc_hd__o31ai_1 _06684_ (.A1(\u_async_wb.u_resp_if.wr_ptr[1] ),
    .A2(_02737_),
    .A3(_02738_),
    .B1(wbs_ack_i),
    .Y(_02739_));
 sky130_fd_sc_hd__a31o_1 _06685_ (.A1(_02736_),
    .A2(_02737_),
    .A3(_02738_),
    .B1(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__or3b_1 _06686_ (.A(_02740_),
    .B(net214),
    .C_N(net176),
    .X(_02741_));
 sky130_fd_sc_hd__nor2_1 _06687_ (.A(_02735_),
    .B(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__clkbuf_2 _06688_ (.A(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__mux2_1 _06689_ (.A0(\u_async_wb.u_resp_if.mem[1][0] ),
    .A1(wbs_dat_i[0]),
    .S(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__clkbuf_1 _06690_ (.A(_02744_),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _06691_ (.A0(\u_async_wb.u_resp_if.mem[1][1] ),
    .A1(wbs_dat_i[1]),
    .S(_02743_),
    .X(_02745_));
 sky130_fd_sc_hd__clkbuf_1 _06692_ (.A(_02745_),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _06693_ (.A0(\u_async_wb.u_resp_if.mem[1][2] ),
    .A1(wbs_dat_i[2]),
    .S(_02743_),
    .X(_02746_));
 sky130_fd_sc_hd__clkbuf_1 _06694_ (.A(_02746_),
    .X(_00308_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06695_ (.A(_02742_),
    .X(_02747_));
 sky130_fd_sc_hd__clkbuf_2 _06696_ (.A(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__mux2_1 _06697_ (.A0(\u_async_wb.u_resp_if.mem[1][3] ),
    .A1(wbs_dat_i[3]),
    .S(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__clkbuf_1 _06698_ (.A(_02749_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _06699_ (.A0(\u_async_wb.u_resp_if.mem[1][4] ),
    .A1(wbs_dat_i[4]),
    .S(_02748_),
    .X(_02750_));
 sky130_fd_sc_hd__clkbuf_1 _06700_ (.A(_02750_),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _06701_ (.A0(\u_async_wb.u_resp_if.mem[1][5] ),
    .A1(wbs_dat_i[5]),
    .S(_02748_),
    .X(_02751_));
 sky130_fd_sc_hd__clkbuf_1 _06702_ (.A(_02751_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _06703_ (.A0(\u_async_wb.u_resp_if.mem[1][6] ),
    .A1(wbs_dat_i[6]),
    .S(_02748_),
    .X(_02752_));
 sky130_fd_sc_hd__clkbuf_1 _06704_ (.A(_02752_),
    .X(_00312_));
 sky130_fd_sc_hd__clkbuf_2 _06705_ (.A(_02747_),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_1 _06706_ (.A0(\u_async_wb.u_resp_if.mem[1][7] ),
    .A1(wbs_dat_i[7]),
    .S(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__clkbuf_1 _06707_ (.A(_02754_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _06708_ (.A0(\u_async_wb.u_resp_if.mem[1][8] ),
    .A1(wbs_dat_i[8]),
    .S(_02753_),
    .X(_02755_));
 sky130_fd_sc_hd__clkbuf_1 _06709_ (.A(_02755_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _06710_ (.A0(\u_async_wb.u_resp_if.mem[1][9] ),
    .A1(wbs_dat_i[9]),
    .S(_02753_),
    .X(_02756_));
 sky130_fd_sc_hd__clkbuf_1 _06711_ (.A(_02756_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _06712_ (.A0(\u_async_wb.u_resp_if.mem[1][10] ),
    .A1(wbs_dat_i[10]),
    .S(_02753_),
    .X(_02757_));
 sky130_fd_sc_hd__clkbuf_1 _06713_ (.A(_02757_),
    .X(_00316_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06714_ (.A(_02742_),
    .X(_02758_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06715_ (.A(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__mux2_1 _06716_ (.A0(\u_async_wb.u_resp_if.mem[1][11] ),
    .A1(wbs_dat_i[11]),
    .S(_02759_),
    .X(_02760_));
 sky130_fd_sc_hd__clkbuf_1 _06717_ (.A(_02760_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _06718_ (.A0(\u_async_wb.u_resp_if.mem[1][12] ),
    .A1(wbs_dat_i[12]),
    .S(_02759_),
    .X(_02761_));
 sky130_fd_sc_hd__clkbuf_1 _06719_ (.A(_02761_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _06720_ (.A0(\u_async_wb.u_resp_if.mem[1][13] ),
    .A1(wbs_dat_i[13]),
    .S(_02759_),
    .X(_02762_));
 sky130_fd_sc_hd__clkbuf_1 _06721_ (.A(_02762_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _06722_ (.A0(\u_async_wb.u_resp_if.mem[1][14] ),
    .A1(wbs_dat_i[14]),
    .S(_02759_),
    .X(_02763_));
 sky130_fd_sc_hd__clkbuf_1 _06723_ (.A(_02763_),
    .X(_00320_));
 sky130_fd_sc_hd__clkbuf_2 _06724_ (.A(_02758_),
    .X(_02764_));
 sky130_fd_sc_hd__mux2_1 _06725_ (.A0(\u_async_wb.u_resp_if.mem[1][15] ),
    .A1(wbs_dat_i[15]),
    .S(_02764_),
    .X(_02765_));
 sky130_fd_sc_hd__clkbuf_1 _06726_ (.A(_02765_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _06727_ (.A0(\u_async_wb.u_resp_if.mem[1][16] ),
    .A1(wbs_dat_i[16]),
    .S(_02764_),
    .X(_02766_));
 sky130_fd_sc_hd__clkbuf_1 _06728_ (.A(_02766_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _06729_ (.A0(\u_async_wb.u_resp_if.mem[1][17] ),
    .A1(wbs_dat_i[17]),
    .S(_02764_),
    .X(_02767_));
 sky130_fd_sc_hd__clkbuf_1 _06730_ (.A(_02767_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _06731_ (.A0(\u_async_wb.u_resp_if.mem[1][18] ),
    .A1(wbs_dat_i[18]),
    .S(_02764_),
    .X(_02768_));
 sky130_fd_sc_hd__clkbuf_1 _06732_ (.A(_02768_),
    .X(_00324_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06733_ (.A(_02758_),
    .X(_02769_));
 sky130_fd_sc_hd__mux2_1 _06734_ (.A0(\u_async_wb.u_resp_if.mem[1][19] ),
    .A1(wbs_dat_i[19]),
    .S(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__clkbuf_1 _06735_ (.A(_02770_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _06736_ (.A0(\u_async_wb.u_resp_if.mem[1][20] ),
    .A1(wbs_dat_i[20]),
    .S(_02769_),
    .X(_02771_));
 sky130_fd_sc_hd__clkbuf_1 _06737_ (.A(_02771_),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _06738_ (.A0(\u_async_wb.u_resp_if.mem[1][21] ),
    .A1(wbs_dat_i[21]),
    .S(_02769_),
    .X(_02772_));
 sky130_fd_sc_hd__clkbuf_1 _06739_ (.A(_02772_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _06740_ (.A0(\u_async_wb.u_resp_if.mem[1][22] ),
    .A1(wbs_dat_i[22]),
    .S(_02769_),
    .X(_02773_));
 sky130_fd_sc_hd__clkbuf_1 _06741_ (.A(_02773_),
    .X(_00328_));
 sky130_fd_sc_hd__clkbuf_2 _06742_ (.A(_02758_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _06743_ (.A0(\u_async_wb.u_resp_if.mem[1][23] ),
    .A1(wbs_dat_i[23]),
    .S(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__clkbuf_1 _06744_ (.A(_02775_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _06745_ (.A0(\u_async_wb.u_resp_if.mem[1][24] ),
    .A1(wbs_dat_i[24]),
    .S(_02774_),
    .X(_02776_));
 sky130_fd_sc_hd__clkbuf_1 _06746_ (.A(_02776_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _06747_ (.A0(\u_async_wb.u_resp_if.mem[1][25] ),
    .A1(wbs_dat_i[25]),
    .S(_02774_),
    .X(_02777_));
 sky130_fd_sc_hd__clkbuf_1 _06748_ (.A(_02777_),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _06749_ (.A0(\u_async_wb.u_resp_if.mem[1][26] ),
    .A1(wbs_dat_i[26]),
    .S(_02774_),
    .X(_02778_));
 sky130_fd_sc_hd__clkbuf_1 _06750_ (.A(_02778_),
    .X(_00332_));
 sky130_fd_sc_hd__clkbuf_2 _06751_ (.A(_02742_),
    .X(_02779_));
 sky130_fd_sc_hd__mux2_1 _06752_ (.A0(\u_async_wb.u_resp_if.mem[1][27] ),
    .A1(wbs_dat_i[27]),
    .S(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__clkbuf_1 _06753_ (.A(_02780_),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _06754_ (.A0(\u_async_wb.u_resp_if.mem[1][28] ),
    .A1(wbs_dat_i[28]),
    .S(_02779_),
    .X(_02781_));
 sky130_fd_sc_hd__clkbuf_1 _06755_ (.A(_02781_),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _06756_ (.A0(\u_async_wb.u_resp_if.mem[1][29] ),
    .A1(wbs_dat_i[29]),
    .S(_02779_),
    .X(_02782_));
 sky130_fd_sc_hd__clkbuf_1 _06757_ (.A(_02782_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _06758_ (.A0(\u_async_wb.u_resp_if.mem[1][30] ),
    .A1(wbs_dat_i[30]),
    .S(_02779_),
    .X(_02783_));
 sky130_fd_sc_hd__clkbuf_1 _06759_ (.A(_02783_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _06760_ (.A0(\u_async_wb.u_resp_if.mem[1][31] ),
    .A1(wbs_dat_i[31]),
    .S(_02747_),
    .X(_02784_));
 sky130_fd_sc_hd__clkbuf_1 _06761_ (.A(_02784_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _06762_ (.A0(\u_async_wb.u_resp_if.mem[1][32] ),
    .A1(wbs_err_i),
    .S(_02747_),
    .X(_02785_));
 sky130_fd_sc_hd__clkbuf_1 _06763_ (.A(_02785_),
    .X(_00338_));
 sky130_fd_sc_hd__clkinv_2 _06764_ (.A(_01531_),
    .Y(_02786_));
 sky130_fd_sc_hd__inv_2 _06765_ (.A(wbs_ack_i),
    .Y(_02787_));
 sky130_fd_sc_hd__mux2_1 _06766_ (.A0(_02786_),
    .A1(\u_async_wb.u_cmd_if.grey_rd_ptr[0] ),
    .S(_02787_),
    .X(_02788_));
 sky130_fd_sc_hd__clkbuf_1 _06767_ (.A(_02788_),
    .X(_00339_));
 sky130_fd_sc_hd__clkbuf_1 _06768_ (.A(_01530_),
    .X(_02789_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06769_ (.A(_01528_),
    .X(_02790_));
 sky130_fd_sc_hd__o21ai_1 _06770_ (.A1(_02789_),
    .A2(_02790_),
    .B1(\u_async_wb.u_cmd_if.grey_rd_ptr[2] ),
    .Y(_02791_));
 sky130_fd_sc_hd__clkbuf_1 _06771_ (.A(wbs_ack_i),
    .X(_02792_));
 sky130_fd_sc_hd__o31a_1 _06772_ (.A1(_02789_),
    .A2(_02790_),
    .A3(\u_async_wb.u_cmd_if.grey_rd_ptr[2] ),
    .B1(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__a22o_1 _06773_ (.A1(_02787_),
    .A2(\u_async_wb.u_cmd_if.grey_rd_ptr[1] ),
    .B1(_02791_),
    .B2(_02793_),
    .X(_00340_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06774_ (.A(_01501_),
    .X(_02794_));
 sky130_fd_sc_hd__a22o_1 _06775_ (.A1(_02453_),
    .A2(_02794_),
    .B1(_01508_),
    .B2(\u_async_wb.PendingRd ),
    .X(_00341_));
 sky130_fd_sc_hd__nand2_1 _06776_ (.A(_01489_),
    .B(_01500_),
    .Y(_02795_));
 sky130_fd_sc_hd__or2_1 _06777_ (.A(_01489_),
    .B(_02794_),
    .X(_02796_));
 sky130_fd_sc_hd__and2_1 _06778_ (.A(_02795_),
    .B(_02796_),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_1 _06779_ (.A(_02797_),
    .X(_00342_));
 sky130_fd_sc_hd__clkbuf_1 _06780_ (.A(_01490_),
    .X(_02798_));
 sky130_fd_sc_hd__or2_2 _06781_ (.A(_02798_),
    .B(_02795_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_2 _06782_ (.A(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__clkbuf_2 _06783_ (.A(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__nand2_1 _06784_ (.A(_02798_),
    .B(_02795_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _06785_ (.A(_02801_),
    .B(_02802_),
    .Y(_00343_));
 sky130_fd_sc_hd__inv_2 _06786_ (.A(_02798_),
    .Y(_02803_));
 sky130_fd_sc_hd__mux2_1 _06787_ (.A0(\u_async_wb.u_cmd_if.grey_wr_ptr[0] ),
    .A1(_02803_),
    .S(_02794_),
    .X(_02804_));
 sky130_fd_sc_hd__clkbuf_1 _06788_ (.A(_02804_),
    .X(_00344_));
 sky130_fd_sc_hd__xnor2_1 _06789_ (.A(\u_async_wb.u_cmd_if.grey_wr_ptr[2] ),
    .B(_01491_),
    .Y(_02805_));
 sky130_fd_sc_hd__mux2_1 _06790_ (.A0(\u_async_wb.u_cmd_if.grey_wr_ptr[1] ),
    .A1(_02805_),
    .S(_02794_),
    .X(_02806_));
 sky130_fd_sc_hd__clkbuf_1 _06791_ (.A(_02806_),
    .X(_00345_));
 sky130_fd_sc_hd__or2_2 _06792_ (.A(_02803_),
    .B(_02795_),
    .X(_02807_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06793_ (.A(_02807_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_2 _06794_ (.A(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__xnor2_1 _06795_ (.A(\u_async_wb.u_cmd_if.grey_wr_ptr[2] ),
    .B(_02809_),
    .Y(_00346_));
 sky130_fd_sc_hd__or2_1 _06796_ (.A(\u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(_02741_),
    .X(_02810_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06797_ (.A(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_2 _06798_ (.A(_02811_),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_1 _06799_ (.A0(wbs_dat_i[0]),
    .A1(\u_async_wb.u_resp_if.mem[0][0] ),
    .S(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__clkbuf_1 _06800_ (.A(_02813_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _06801_ (.A0(wbs_dat_i[1]),
    .A1(\u_async_wb.u_resp_if.mem[0][1] ),
    .S(_02812_),
    .X(_02814_));
 sky130_fd_sc_hd__clkbuf_1 _06802_ (.A(_02814_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _06803_ (.A0(wbs_dat_i[2]),
    .A1(\u_async_wb.u_resp_if.mem[0][2] ),
    .S(_02812_),
    .X(_02815_));
 sky130_fd_sc_hd__clkbuf_1 _06804_ (.A(_02815_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _06805_ (.A0(wbs_dat_i[3]),
    .A1(\u_async_wb.u_resp_if.mem[0][3] ),
    .S(_02812_),
    .X(_02816_));
 sky130_fd_sc_hd__clkbuf_1 _06806_ (.A(_02816_),
    .X(_00350_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06807_ (.A(_02811_),
    .X(_02817_));
 sky130_fd_sc_hd__mux2_1 _06808_ (.A0(wbs_dat_i[4]),
    .A1(\u_async_wb.u_resp_if.mem[0][4] ),
    .S(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__clkbuf_1 _06809_ (.A(_02818_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _06810_ (.A0(wbs_dat_i[5]),
    .A1(\u_async_wb.u_resp_if.mem[0][5] ),
    .S(_02817_),
    .X(_02819_));
 sky130_fd_sc_hd__clkbuf_1 _06811_ (.A(_02819_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _06812_ (.A0(wbs_dat_i[6]),
    .A1(\u_async_wb.u_resp_if.mem[0][6] ),
    .S(_02817_),
    .X(_02820_));
 sky130_fd_sc_hd__clkbuf_1 _06813_ (.A(_02820_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _06814_ (.A0(wbs_dat_i[7]),
    .A1(\u_async_wb.u_resp_if.mem[0][7] ),
    .S(_02817_),
    .X(_02821_));
 sky130_fd_sc_hd__clkbuf_1 _06815_ (.A(_02821_),
    .X(_00354_));
 sky130_fd_sc_hd__clkbuf_2 _06816_ (.A(_02811_),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_1 _06817_ (.A0(wbs_dat_i[8]),
    .A1(\u_async_wb.u_resp_if.mem[0][8] ),
    .S(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_1 _06818_ (.A(_02823_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _06819_ (.A0(wbs_dat_i[9]),
    .A1(\u_async_wb.u_resp_if.mem[0][9] ),
    .S(_02822_),
    .X(_02824_));
 sky130_fd_sc_hd__clkbuf_1 _06820_ (.A(_02824_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _06821_ (.A0(wbs_dat_i[10]),
    .A1(\u_async_wb.u_resp_if.mem[0][10] ),
    .S(_02822_),
    .X(_02825_));
 sky130_fd_sc_hd__clkbuf_1 _06822_ (.A(_02825_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _06823_ (.A0(wbs_dat_i[11]),
    .A1(\u_async_wb.u_resp_if.mem[0][11] ),
    .S(_02822_),
    .X(_02826_));
 sky130_fd_sc_hd__clkbuf_1 _06824_ (.A(_02826_),
    .X(_00358_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06825_ (.A(_02810_),
    .X(_02827_));
 sky130_fd_sc_hd__clkbuf_2 _06826_ (.A(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _06827_ (.A0(wbs_dat_i[12]),
    .A1(\u_async_wb.u_resp_if.mem[0][12] ),
    .S(_02828_),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_1 _06828_ (.A(_02829_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _06829_ (.A0(wbs_dat_i[13]),
    .A1(\u_async_wb.u_resp_if.mem[0][13] ),
    .S(_02828_),
    .X(_02830_));
 sky130_fd_sc_hd__clkbuf_1 _06830_ (.A(_02830_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _06831_ (.A0(wbs_dat_i[14]),
    .A1(\u_async_wb.u_resp_if.mem[0][14] ),
    .S(_02828_),
    .X(_02831_));
 sky130_fd_sc_hd__clkbuf_1 _06832_ (.A(_02831_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _06833_ (.A0(wbs_dat_i[15]),
    .A1(\u_async_wb.u_resp_if.mem[0][15] ),
    .S(_02828_),
    .X(_02832_));
 sky130_fd_sc_hd__clkbuf_1 _06834_ (.A(_02832_),
    .X(_00362_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06835_ (.A(_02827_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _06836_ (.A0(wbs_dat_i[16]),
    .A1(\u_async_wb.u_resp_if.mem[0][16] ),
    .S(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__clkbuf_1 _06837_ (.A(_02834_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _06838_ (.A0(wbs_dat_i[17]),
    .A1(\u_async_wb.u_resp_if.mem[0][17] ),
    .S(_02833_),
    .X(_02835_));
 sky130_fd_sc_hd__clkbuf_1 _06839_ (.A(_02835_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _06840_ (.A0(wbs_dat_i[18]),
    .A1(\u_async_wb.u_resp_if.mem[0][18] ),
    .S(_02833_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _06841_ (.A(_02836_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _06842_ (.A0(wbs_dat_i[19]),
    .A1(\u_async_wb.u_resp_if.mem[0][19] ),
    .S(_02833_),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_1 _06843_ (.A(_02837_),
    .X(_00366_));
 sky130_fd_sc_hd__clkbuf_2 _06844_ (.A(_02827_),
    .X(_02838_));
 sky130_fd_sc_hd__mux2_1 _06845_ (.A0(wbs_dat_i[20]),
    .A1(\u_async_wb.u_resp_if.mem[0][20] ),
    .S(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__clkbuf_1 _06846_ (.A(_02839_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _06847_ (.A0(wbs_dat_i[21]),
    .A1(\u_async_wb.u_resp_if.mem[0][21] ),
    .S(_02838_),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_1 _06848_ (.A(_02840_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _06849_ (.A0(wbs_dat_i[22]),
    .A1(\u_async_wb.u_resp_if.mem[0][22] ),
    .S(_02838_),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_1 _06850_ (.A(_02841_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _06851_ (.A0(wbs_dat_i[23]),
    .A1(\u_async_wb.u_resp_if.mem[0][23] ),
    .S(_02838_),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _06852_ (.A(_02842_),
    .X(_00370_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06853_ (.A(_02827_),
    .X(_02843_));
 sky130_fd_sc_hd__mux2_1 _06854_ (.A0(wbs_dat_i[24]),
    .A1(\u_async_wb.u_resp_if.mem[0][24] ),
    .S(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _06855_ (.A(_02844_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _06856_ (.A0(wbs_dat_i[25]),
    .A1(\u_async_wb.u_resp_if.mem[0][25] ),
    .S(_02843_),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _06857_ (.A(_02845_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _06858_ (.A0(wbs_dat_i[26]),
    .A1(\u_async_wb.u_resp_if.mem[0][26] ),
    .S(_02843_),
    .X(_02846_));
 sky130_fd_sc_hd__clkbuf_1 _06859_ (.A(_02846_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _06860_ (.A0(wbs_dat_i[27]),
    .A1(\u_async_wb.u_resp_if.mem[0][27] ),
    .S(_02843_),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _06861_ (.A(_02847_),
    .X(_00374_));
 sky130_fd_sc_hd__clkbuf_2 _06862_ (.A(_02810_),
    .X(_02848_));
 sky130_fd_sc_hd__mux2_1 _06863_ (.A0(wbs_dat_i[28]),
    .A1(\u_async_wb.u_resp_if.mem[0][28] ),
    .S(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _06864_ (.A(_02849_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _06865_ (.A0(wbs_dat_i[29]),
    .A1(\u_async_wb.u_resp_if.mem[0][29] ),
    .S(_02848_),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _06866_ (.A(_02850_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _06867_ (.A0(wbs_dat_i[30]),
    .A1(\u_async_wb.u_resp_if.mem[0][30] ),
    .S(_02848_),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _06868_ (.A(_02851_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _06869_ (.A0(wbs_dat_i[31]),
    .A1(\u_async_wb.u_resp_if.mem[0][31] ),
    .S(_02848_),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _06870_ (.A(_02852_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _06871_ (.A0(wbs_err_i),
    .A1(\u_async_wb.u_resp_if.mem[0][32] ),
    .S(_02811_),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _06872_ (.A(_02853_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _06873_ (.A0(_02686_),
    .A1(\u_async_wb.u_resp_if.grey_rd_ptr[0] ),
    .S(_02683_),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _06874_ (.A(_02854_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _06875_ (.A0(_01505_),
    .A1(\u_async_wb.u_resp_if.grey_rd_ptr[1] ),
    .S(_02683_),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _06876_ (.A(_02855_),
    .X(_00381_));
 sky130_fd_sc_hd__xor2_1 _06877_ (.A(_02790_),
    .B(_02792_),
    .X(_00382_));
 sky130_fd_sc_hd__a21oi_1 _06878_ (.A1(_02790_),
    .A2(_02792_),
    .B1(_02789_),
    .Y(_02856_));
 sky130_fd_sc_hd__and3_1 _06879_ (.A(_02789_),
    .B(_01528_),
    .C(_02792_),
    .X(_02857_));
 sky130_fd_sc_hd__nor2_1 _06880_ (.A(_02856_),
    .B(_02857_),
    .Y(_00383_));
 sky130_fd_sc_hd__xor2_1 _06881_ (.A(\u_async_wb.u_cmd_if.grey_rd_ptr[2] ),
    .B(_02857_),
    .X(_00384_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06882_ (.A(_02741_),
    .X(_02858_));
 sky130_fd_sc_hd__and2_1 _06883_ (.A(_02735_),
    .B(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__nor2_1 _06884_ (.A(_02743_),
    .B(_02859_),
    .Y(_00385_));
 sky130_fd_sc_hd__xor2_1 _06885_ (.A(\u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(_02736_),
    .X(_02860_));
 sky130_fd_sc_hd__mux2_1 _06886_ (.A0(_02860_),
    .A1(_02736_),
    .S(_02858_),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_1 _06887_ (.A(_02861_),
    .X(_00386_));
 sky130_fd_sc_hd__clkinv_2 _06888_ (.A(_02736_),
    .Y(_02862_));
 sky130_fd_sc_hd__mux2_1 _06889_ (.A0(_02862_),
    .A1(\u_async_wb.u_resp_if.grey_wr_ptr[0] ),
    .S(_02858_),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _06890_ (.A(_02863_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _06891_ (.A0(_02860_),
    .A1(\u_async_wb.u_resp_if.grey_wr_ptr[1] ),
    .S(_02858_),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_1 _06892_ (.A(_02864_),
    .X(_00388_));
 sky130_fd_sc_hd__nand2_1 _06893_ (.A(wbm_cyc_i),
    .B(net367),
    .Y(_02865_));
 sky130_fd_sc_hd__a21oi_1 _06894_ (.A1(wbm_cyc_i),
    .A2(wbm_stb_i),
    .B1(\u_uart2wb.u_async_reg_bus.out_reg_cs ),
    .Y(_02866_));
 sky130_fd_sc_hd__or2_1 _06895_ (.A(_01733_),
    .B(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__a31o_1 _06896_ (.A1(_01472_),
    .A2(_01731_),
    .A3(_02867_),
    .B1(_01740_),
    .X(_02868_));
 sky130_fd_sc_hd__inv_2 _06897_ (.A(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__a21o_1 _06898_ (.A1(_02865_),
    .A2(_01732_),
    .B1(_02868_),
    .X(_02870_));
 sky130_fd_sc_hd__a32o_1 _06899_ (.A1(\u_uart2wb.u_async_reg_bus.out_reg_cs ),
    .A2(_02865_),
    .A3(_02869_),
    .B1(_02870_),
    .B2(\u_arb.gnt[0] ),
    .X(_00389_));
 sky130_fd_sc_hd__nor2_1 _06900_ (.A(_01732_),
    .B(_02868_),
    .Y(_02871_));
 sky130_fd_sc_hd__o22a_1 _06901_ (.A1(_02866_),
    .A2(_02868_),
    .B1(_02871_),
    .B2(_01731_),
    .X(_00390_));
 sky130_fd_sc_hd__and4_1 _06902_ (.A(\u_uart2wb.u_msg.wait_cnt[0] ),
    .B(\u_uart2wb.u_msg.wait_cnt[1] ),
    .C(\u_uart2wb.u_msg.wait_cnt[3] ),
    .D(\u_uart2wb.u_msg.wait_cnt[2] ),
    .X(_02872_));
 sky130_fd_sc_hd__and4_1 _06903_ (.A(\u_uart2wb.u_msg.wait_cnt[5] ),
    .B(\u_uart2wb.u_msg.wait_cnt[4] ),
    .C(\u_uart2wb.u_msg.wait_cnt[6] ),
    .D(_02872_),
    .X(_02873_));
 sky130_fd_sc_hd__and2_1 _06904_ (.A(\u_uart2wb.u_msg.wait_cnt[7] ),
    .B(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__or2_1 _06905_ (.A(\u_uart2wb.u_msg.State[1] ),
    .B(\u_uart2wb.u_msg.State[0] ),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_1 _06906_ (.A(\u_uart2wb.u_msg.State[2] ),
    .X(_02876_));
 sky130_fd_sc_hd__clkbuf_1 _06907_ (.A(\u_uart2wb.u_msg.State[3] ),
    .X(_02877_));
 sky130_fd_sc_hd__or2_1 _06908_ (.A(_02876_),
    .B(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__clkbuf_2 _06909_ (.A(_02878_),
    .X(_02879_));
 sky130_fd_sc_hd__nor2_2 _06910_ (.A(_02875_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__and3b_1 _06911_ (.A_N(_02874_),
    .B(_02880_),
    .C(_01158_),
    .X(_02881_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06912_ (.A(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__xor2_1 _06913_ (.A(\u_uart2wb.u_msg.wait_cnt[0] ),
    .B(_02882_),
    .X(_00391_));
 sky130_fd_sc_hd__and3_1 _06914_ (.A(\u_uart2wb.u_msg.wait_cnt[0] ),
    .B(\u_uart2wb.u_msg.wait_cnt[1] ),
    .C(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__a21oi_1 _06915_ (.A1(\u_uart2wb.u_msg.wait_cnt[0] ),
    .A2(_02882_),
    .B1(\u_uart2wb.u_msg.wait_cnt[1] ),
    .Y(_02884_));
 sky130_fd_sc_hd__nor2_1 _06916_ (.A(_02883_),
    .B(_02884_),
    .Y(_00392_));
 sky130_fd_sc_hd__xor2_1 _06917_ (.A(\u_uart2wb.u_msg.wait_cnt[2] ),
    .B(_02883_),
    .X(_00393_));
 sky130_fd_sc_hd__and3_1 _06918_ (.A(\u_uart2wb.u_msg.wait_cnt[3] ),
    .B(\u_uart2wb.u_msg.wait_cnt[2] ),
    .C(_02883_),
    .X(_02885_));
 sky130_fd_sc_hd__a21oi_1 _06919_ (.A1(\u_uart2wb.u_msg.wait_cnt[2] ),
    .A2(_02883_),
    .B1(\u_uart2wb.u_msg.wait_cnt[3] ),
    .Y(_02886_));
 sky130_fd_sc_hd__nor2_1 _06920_ (.A(_02885_),
    .B(_02886_),
    .Y(_00394_));
 sky130_fd_sc_hd__xor2_1 _06921_ (.A(\u_uart2wb.u_msg.wait_cnt[4] ),
    .B(_02885_),
    .X(_00395_));
 sky130_fd_sc_hd__and3_1 _06922_ (.A(\u_uart2wb.u_msg.wait_cnt[5] ),
    .B(\u_uart2wb.u_msg.wait_cnt[4] ),
    .C(_02885_),
    .X(_02887_));
 sky130_fd_sc_hd__a21oi_1 _06923_ (.A1(\u_uart2wb.u_msg.wait_cnt[4] ),
    .A2(_02885_),
    .B1(\u_uart2wb.u_msg.wait_cnt[5] ),
    .Y(_02888_));
 sky130_fd_sc_hd__nor2_1 _06924_ (.A(_02887_),
    .B(_02888_),
    .Y(_00396_));
 sky130_fd_sc_hd__o2bb2a_1 _06925_ (.A1_N(_02873_),
    .A2_N(_02882_),
    .B1(_02887_),
    .B2(\u_uart2wb.u_msg.wait_cnt[6] ),
    .X(_00397_));
 sky130_fd_sc_hd__a31o_1 _06926_ (.A1(_01159_),
    .A2(_02873_),
    .A3(_02880_),
    .B1(\u_uart2wb.u_msg.wait_cnt[7] ),
    .X(_00398_));
 sky130_fd_sc_hd__inv_2 _06927_ (.A(net335),
    .Y(_00036_));
 sky130_fd_sc_hd__inv_2 _06928_ (.A(net335),
    .Y(_00037_));
 sky130_fd_sc_hd__inv_2 _06929_ (.A(\u_uart2wb.u_msg.State[1] ),
    .Y(_02889_));
 sky130_fd_sc_hd__or2_1 _06930_ (.A(_02889_),
    .B(\u_uart2wb.u_msg.State[0] ),
    .X(_02890_));
 sky130_fd_sc_hd__inv_2 _06931_ (.A(\u_uart2wb.u_msg.State[3] ),
    .Y(_02891_));
 sky130_fd_sc_hd__or2_1 _06932_ (.A(\u_uart2wb.u_msg.State[2] ),
    .B(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__clkbuf_1 _06933_ (.A(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__nor2_1 _06934_ (.A(_02890_),
    .B(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__clkbuf_1 _06935_ (.A(_02894_),
    .X(_02895_));
 sky130_fd_sc_hd__nor2_1 _06936_ (.A(_02875_),
    .B(_02892_),
    .Y(_02896_));
 sky130_fd_sc_hd__nand2_1 _06937_ (.A(_02889_),
    .B(\u_uart2wb.u_msg.State[0] ),
    .Y(_02897_));
 sky130_fd_sc_hd__clkbuf_1 _06938_ (.A(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__and2_1 _06939_ (.A(_02890_),
    .B(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__nor2_1 _06940_ (.A(_02878_),
    .B(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__clkbuf_1 _06941_ (.A(\u_uart2wb.u_msg.State[1] ),
    .X(_02901_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06942_ (.A(\u_uart2wb.u_msg.State[0] ),
    .X(_02902_));
 sky130_fd_sc_hd__nand2_1 _06943_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__clkbuf_1 _06944_ (.A(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__nor2_1 _06945_ (.A(_02877_),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__nor2_1 _06946_ (.A(_02893_),
    .B(_02898_),
    .Y(_02906_));
 sky130_fd_sc_hd__or2_1 _06947_ (.A(_02905_),
    .B(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__or3_2 _06948_ (.A(_02896_),
    .B(_02900_),
    .C(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__nor2_1 _06949_ (.A(_02895_),
    .B(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__or3_1 _06950_ (.A(\u_uart2wb.u_msg.TxMsgSize[1] ),
    .B(\u_uart2wb.u_msg.TxMsgSize[0] ),
    .C(\u_uart2wb.u_msg.TxMsgSize[2] ),
    .X(_02910_));
 sky130_fd_sc_hd__or2_1 _06951_ (.A(\u_uart2wb.u_msg.TxMsgSize[3] ),
    .B(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__o21ai_1 _06952_ (.A1(\u_uart2wb.u_msg.TxMsgSize[4] ),
    .A2(_02911_),
    .B1(\u_uart2wb.tx_rd ),
    .Y(_02912_));
 sky130_fd_sc_hd__nand2_1 _06953_ (.A(_02876_),
    .B(_02891_),
    .Y(_02913_));
 sky130_fd_sc_hd__clkbuf_1 _06954_ (.A(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__nor2_1 _06955_ (.A(_02903_),
    .B(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__nor2_1 _06956_ (.A(_02896_),
    .B(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__nor2_2 _06957_ (.A(\u_uart2wb.reg_ack ),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__inv_2 _06958_ (.A(net243),
    .Y(_02918_));
 sky130_fd_sc_hd__a211o_1 _06959_ (.A1(_02894_),
    .A2(_02912_),
    .B1(_02917_),
    .C1(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_1 _06960_ (.A(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__or2_1 _06961_ (.A(_02909_),
    .B(_02920_),
    .X(_02921_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06962_ (.A(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__inv_2 _06963_ (.A(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06964_ (.A(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06965_ (.A(_02924_),
    .X(_02925_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06966_ (.A(_02895_),
    .X(_02926_));
 sky130_fd_sc_hd__clkbuf_2 _06967_ (.A(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_1 _06968_ (.A(_02927_),
    .X(_02928_));
 sky130_fd_sc_hd__clkbuf_1 _06969_ (.A(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__clkbuf_2 _06970_ (.A(_02915_),
    .X(_02930_));
 sky130_fd_sc_hd__clkbuf_2 _06971_ (.A(_02930_),
    .X(_02931_));
 sky130_fd_sc_hd__clkbuf_1 _06972_ (.A(_02922_),
    .X(_02932_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06973_ (.A(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__a211o_1 _06974_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[48] ),
    .A2(_02929_),
    .B1(_02931_),
    .C1(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__o21a_1 _06975_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[56] ),
    .A2(_02925_),
    .B1(_02934_),
    .X(_00399_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06976_ (.A(_02890_),
    .X(_02935_));
 sky130_fd_sc_hd__or2_1 _06977_ (.A(_02935_),
    .B(_02893_),
    .X(_02936_));
 sky130_fd_sc_hd__or2_1 _06978_ (.A(_02893_),
    .B(_02898_),
    .X(_02937_));
 sky130_fd_sc_hd__nand2_1 _06979_ (.A(_02936_),
    .B(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__clkbuf_1 _06980_ (.A(_02905_),
    .X(_02939_));
 sky130_fd_sc_hd__nor2_2 _06981_ (.A(_02879_),
    .B(_02935_),
    .Y(_02940_));
 sky130_fd_sc_hd__or2_1 _06982_ (.A(_02939_),
    .B(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__nor2_1 _06983_ (.A(_02938_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__clkbuf_2 _06984_ (.A(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06985_ (.A(_02906_),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_1 _06986_ (.A(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__clkbuf_2 _06987_ (.A(_02945_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_2 _06988_ (.A(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06989_ (.A(_02921_),
    .X(_02948_));
 sky130_fd_sc_hd__clkbuf_2 _06990_ (.A(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__nor2_2 _06991_ (.A(_02879_),
    .B(_02904_),
    .Y(_02950_));
 sky130_fd_sc_hd__a2111o_1 _06992_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[49] ),
    .A2(_02928_),
    .B1(_02947_),
    .C1(_02949_),
    .D1(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__o22a_1 _06993_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[57] ),
    .A2(_02924_),
    .B1(_02943_),
    .B2(_02951_),
    .X(_00400_));
 sky130_fd_sc_hd__nor2_2 _06994_ (.A(_02889_),
    .B(_02902_),
    .Y(_02952_));
 sky130_fd_sc_hd__clkbuf_2 _06995_ (.A(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__clkbuf_1 _06996_ (.A(_02876_),
    .X(_02954_));
 sky130_fd_sc_hd__or3b_2 _06997_ (.A(_02954_),
    .B(_02891_),
    .C_N(_02904_),
    .X(_02955_));
 sky130_fd_sc_hd__a211o_1 _06998_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[50] ),
    .A2(_02953_),
    .B1(_02933_),
    .C1(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__o21a_1 _06999_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[58] ),
    .A2(_02925_),
    .B1(_02956_),
    .X(_00401_));
 sky130_fd_sc_hd__clkbuf_1 _07000_ (.A(_02926_),
    .X(_02957_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07001_ (.A(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07002_ (.A(_02945_),
    .X(_02959_));
 sky130_fd_sc_hd__clkbuf_2 _07003_ (.A(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07004_ (.A(_02896_),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_2 _07005_ (.A(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__nor2_1 _07006_ (.A(_02889_),
    .B(_02879_),
    .Y(_02963_));
 sky130_fd_sc_hd__or2_1 _07007_ (.A(_02962_),
    .B(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__clkbuf_2 _07008_ (.A(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__a211o_1 _07009_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[51] ),
    .A2(_02958_),
    .B1(_02960_),
    .C1(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07010_ (.A(_02932_),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_1 _07011_ (.A0(_02966_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[59] ),
    .S(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__clkbuf_1 _07012_ (.A(_02968_),
    .X(_00402_));
 sky130_fd_sc_hd__clkbuf_1 _07013_ (.A(_02932_),
    .X(_02969_));
 sky130_fd_sc_hd__a211o_1 _07014_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[52] ),
    .A2(_02929_),
    .B1(_02969_),
    .C1(_02965_),
    .X(_02970_));
 sky130_fd_sc_hd__o21a_1 _07015_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[60] ),
    .A2(_02925_),
    .B1(_02970_),
    .X(_00403_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07016_ (.A(_02928_),
    .X(_02971_));
 sky130_fd_sc_hd__or2_1 _07017_ (.A(_02961_),
    .B(_02941_),
    .X(_02972_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07018_ (.A(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__a211o_1 _07019_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[53] ),
    .A2(_02971_),
    .B1(_02969_),
    .C1(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__o21a_1 _07020_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[61] ),
    .A2(_02925_),
    .B1(_02974_),
    .X(_00404_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07021_ (.A(_02923_),
    .X(_02975_));
 sky130_fd_sc_hd__nor2_2 _07022_ (.A(_02938_),
    .B(_02972_),
    .Y(_02976_));
 sky130_fd_sc_hd__or2_1 _07023_ (.A(_02930_),
    .B(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__a211o_1 _07024_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[54] ),
    .A2(_02971_),
    .B1(_02969_),
    .C1(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__o21a_1 _07025_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[62] ),
    .A2(_02975_),
    .B1(_02978_),
    .X(_00405_));
 sky130_fd_sc_hd__clkbuf_1 _07026_ (.A(_02922_),
    .X(_02979_));
 sky130_fd_sc_hd__clkbuf_1 _07027_ (.A(_02940_),
    .X(_02980_));
 sky130_fd_sc_hd__clkbuf_1 _07028_ (.A(_02894_),
    .X(_02981_));
 sky130_fd_sc_hd__clkbuf_2 _07029_ (.A(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__clkbuf_2 _07030_ (.A(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__nor2_1 _07031_ (.A(\u_uart2wb.reg_rdata[29] ),
    .B(\u_uart2wb.reg_rdata[30] ),
    .Y(_02984_));
 sky130_fd_sc_hd__clkbuf_1 _07032_ (.A(\u_uart2wb.reg_rdata[31] ),
    .X(_02985_));
 sky130_fd_sc_hd__and3b_1 _07033_ (.A_N(_02984_),
    .B(_02944_),
    .C(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__inv_2 _07034_ (.A(\u_uart2wb.reg_rdata[31] ),
    .Y(_02987_));
 sky130_fd_sc_hd__o21a_1 _07035_ (.A1(_02987_),
    .A2(_02984_),
    .B1(_02944_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _07036_ (.A0(_02986_),
    .A1(_02988_),
    .S(\u_uart2wb.reg_rdata[28] ),
    .X(_02989_));
 sky130_fd_sc_hd__a21o_1 _07037_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[112] ),
    .A2(_02983_),
    .B1(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__or4_1 _07038_ (.A(_02979_),
    .B(_02980_),
    .C(_02977_),
    .D(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__o21a_1 _07039_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[120] ),
    .A2(_02975_),
    .B1(_02991_),
    .X(_00406_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07040_ (.A(_02948_),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _07041_ (.A(_02906_),
    .X(_02993_));
 sky130_fd_sc_hd__nor2_1 _07042_ (.A(_02981_),
    .B(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07043_ (.A(_02994_),
    .X(_02995_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07044_ (.A(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_1 _07045_ (.A(_02952_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_1 _07046_ (.A(_02945_),
    .X(_02998_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07047_ (.A(_02998_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_1 _07048_ (.A(\u_uart2wb.reg_rdata[29] ),
    .X(_03000_));
 sky130_fd_sc_hd__or2_1 _07049_ (.A(\u_uart2wb.reg_rdata[28] ),
    .B(_02987_),
    .X(_03001_));
 sky130_fd_sc_hd__and4bb_1 _07050_ (.A_N(\u_uart2wb.reg_rdata[28] ),
    .B_N(_03000_),
    .C(\u_uart2wb.reg_rdata[30] ),
    .D(_02985_),
    .X(_03002_));
 sky130_fd_sc_hd__a21o_1 _07051_ (.A1(_03000_),
    .A2(_03001_),
    .B1(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__a22o_1 _07052_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[113] ),
    .A2(_02997_),
    .B1(_02999_),
    .B2(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__or3_1 _07053_ (.A(_02992_),
    .B(_02996_),
    .C(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__o21a_1 _07054_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[121] ),
    .A2(_02975_),
    .B1(_03005_),
    .X(_00407_));
 sky130_fd_sc_hd__o211a_1 _07055_ (.A1(_03000_),
    .A2(_03001_),
    .B1(_02946_),
    .C1(\u_uart2wb.reg_rdata[30] ),
    .X(_03006_));
 sky130_fd_sc_hd__a211o_1 _07056_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[114] ),
    .A2(_02958_),
    .B1(_02940_),
    .C1(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__mux2_1 _07057_ (.A0(_03007_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[122] ),
    .S(_02967_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_1 _07058_ (.A(_03008_),
    .X(_00408_));
 sky130_fd_sc_hd__a32o_1 _07059_ (.A1(_02985_),
    .A2(_02960_),
    .A3(_02984_),
    .B1(\u_uart2wb.u_msg.TxMsgBuf[115] ),
    .B2(_02958_),
    .X(_03009_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07060_ (.A(_02932_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_1 _07061_ (.A0(_03009_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[123] ),
    .S(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__clkbuf_1 _07062_ (.A(_03011_),
    .X(_00409_));
 sky130_fd_sc_hd__a211o_1 _07063_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[116] ),
    .A2(_02958_),
    .B1(_02965_),
    .C1(_02988_),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_1 _07064_ (.A0(_03012_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[124] ),
    .S(_03010_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_1 _07065_ (.A(_03013_),
    .X(_00410_));
 sky130_fd_sc_hd__clkbuf_1 _07066_ (.A(_02926_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_2 _07067_ (.A(_03014_),
    .X(_03015_));
 sky130_fd_sc_hd__a211o_1 _07068_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[117] ),
    .A2(_03015_),
    .B1(_02941_),
    .C1(_02988_),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_1 _07069_ (.A0(_03016_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[125] ),
    .S(_03010_),
    .X(_03017_));
 sky130_fd_sc_hd__clkbuf_1 _07070_ (.A(_03017_),
    .X(_00411_));
 sky130_fd_sc_hd__a211o_1 _07071_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[118] ),
    .A2(_03015_),
    .B1(_02996_),
    .C1(_02986_),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_1 _07072_ (.A0(_03018_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[126] ),
    .S(_03010_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_1 _07073_ (.A(_03019_),
    .X(_00412_));
 sky130_fd_sc_hd__or2_1 _07074_ (.A(_02961_),
    .B(_02915_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_1 _07075_ (.A(_03020_),
    .X(_03021_));
 sky130_fd_sc_hd__o21a_1 _07076_ (.A1(\u_uart2wb.reg_rdata[5] ),
    .A2(\u_uart2wb.reg_rdata[6] ),
    .B1(\u_uart2wb.reg_rdata[7] ),
    .X(_03022_));
 sky130_fd_sc_hd__and2_1 _07077_ (.A(_02993_),
    .B(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_2 _07078_ (.A(_02937_),
    .X(_03024_));
 sky130_fd_sc_hd__nor2_1 _07079_ (.A(_03024_),
    .B(_03022_),
    .Y(_03025_));
 sky130_fd_sc_hd__mux2_1 _07080_ (.A0(_03023_),
    .A1(_03025_),
    .S(\u_uart2wb.reg_rdata[4] ),
    .X(_03026_));
 sky130_fd_sc_hd__a211o_1 _07081_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[64] ),
    .A2(_03015_),
    .B1(_03021_),
    .C1(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07082_ (.A(_02922_),
    .X(_03028_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07083_ (.A(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__mux2_1 _07084_ (.A0(_03027_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[72] ),
    .S(_03029_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _07085_ (.A(_03030_),
    .X(_00413_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07086_ (.A(\u_uart2wb.reg_rdata[6] ),
    .X(_03031_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07087_ (.A(\u_uart2wb.reg_rdata[5] ),
    .X(_03032_));
 sky130_fd_sc_hd__or2b_1 _07088_ (.A(\u_uart2wb.reg_rdata[4] ),
    .B_N(\u_uart2wb.reg_rdata[7] ),
    .X(_03033_));
 sky130_fd_sc_hd__nor2_1 _07089_ (.A(_03032_),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__and3_1 _07090_ (.A(_03031_),
    .B(_02946_),
    .C(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__a32o_1 _07091_ (.A1(_03032_),
    .A2(_02946_),
    .A3(_03033_),
    .B1(\u_uart2wb.u_msg.TxMsgBuf[65] ),
    .B2(_02983_),
    .X(_03036_));
 sky130_fd_sc_hd__or4_1 _07092_ (.A(_02979_),
    .B(_02972_),
    .C(_03035_),
    .D(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__o21a_1 _07093_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[73] ),
    .A2(_02975_),
    .B1(_03037_),
    .X(_00414_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07094_ (.A(_02945_),
    .X(_03038_));
 sky130_fd_sc_hd__and3b_1 _07095_ (.A_N(_03034_),
    .B(_03038_),
    .C(_03031_),
    .X(_03039_));
 sky130_fd_sc_hd__nor2_1 _07096_ (.A(_03020_),
    .B(_02938_),
    .Y(_03040_));
 sky130_fd_sc_hd__a211o_1 _07097_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[66] ),
    .A2(_03015_),
    .B1(_03039_),
    .C1(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__mux2_1 _07098_ (.A0(_03041_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[74] ),
    .S(_03029_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _07099_ (.A(_03042_),
    .X(_00415_));
 sky130_fd_sc_hd__clkbuf_1 _07100_ (.A(_03014_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _07101_ (.A(_02944_),
    .X(_03044_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07102_ (.A(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__and4bb_1 _07103_ (.A_N(_03032_),
    .B_N(_03031_),
    .C(_03045_),
    .D(\u_uart2wb.reg_rdata[7] ),
    .X(_03046_));
 sky130_fd_sc_hd__a211o_1 _07104_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[67] ),
    .A2(_03043_),
    .B1(_02963_),
    .C1(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__mux2_1 _07105_ (.A0(_03047_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[75] ),
    .S(_03029_),
    .X(_03048_));
 sky130_fd_sc_hd__clkbuf_1 _07106_ (.A(_03048_),
    .X(_00416_));
 sky130_fd_sc_hd__a211o_1 _07107_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[68] ),
    .A2(_03043_),
    .B1(_02964_),
    .C1(_03025_),
    .X(_03049_));
 sky130_fd_sc_hd__mux2_1 _07108_ (.A0(_03049_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[76] ),
    .S(_03029_),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_1 _07109_ (.A(_03050_),
    .X(_00417_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07110_ (.A(_02994_),
    .X(_03051_));
 sky130_fd_sc_hd__a211o_1 _07111_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[69] ),
    .A2(_03043_),
    .B1(_03051_),
    .C1(_03025_),
    .X(_03052_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07112_ (.A(_03028_),
    .X(_03053_));
 sky130_fd_sc_hd__mux2_1 _07113_ (.A0(_03052_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[77] ),
    .S(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _07114_ (.A(_03054_),
    .X(_00418_));
 sky130_fd_sc_hd__or2_1 _07115_ (.A(_02915_),
    .B(_02942_),
    .X(_03055_));
 sky130_fd_sc_hd__a211o_1 _07116_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[70] ),
    .A2(_03043_),
    .B1(_03023_),
    .C1(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__mux2_1 _07117_ (.A0(_03056_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[78] ),
    .S(_03053_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_1 _07118_ (.A(_03057_),
    .X(_00419_));
 sky130_fd_sc_hd__clkbuf_1 _07119_ (.A(_03014_),
    .X(_03058_));
 sky130_fd_sc_hd__o21a_1 _07120_ (.A1(\u_uart2wb.reg_rdata[9] ),
    .A2(\u_uart2wb.reg_rdata[10] ),
    .B1(\u_uart2wb.reg_rdata[11] ),
    .X(_03059_));
 sky130_fd_sc_hd__and2_1 _07121_ (.A(_03044_),
    .B(_03059_),
    .X(_03060_));
 sky130_fd_sc_hd__nor2_1 _07122_ (.A(_03024_),
    .B(_03059_),
    .Y(_03061_));
 sky130_fd_sc_hd__mux2_1 _07123_ (.A0(_03060_),
    .A1(_03061_),
    .S(\u_uart2wb.reg_rdata[8] ),
    .X(_03062_));
 sky130_fd_sc_hd__a211o_1 _07124_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[72] ),
    .A2(_03058_),
    .B1(_02931_),
    .C1(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_1 _07125_ (.A0(_03063_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[80] ),
    .S(_03053_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _07126_ (.A(_03064_),
    .X(_00420_));
 sky130_fd_sc_hd__clkbuf_2 _07127_ (.A(_02923_),
    .X(_03065_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07128_ (.A(\u_uart2wb.reg_rdata[10] ),
    .X(_03066_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07129_ (.A(_03038_),
    .X(_03067_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07130_ (.A(\u_uart2wb.reg_rdata[9] ),
    .X(_03068_));
 sky130_fd_sc_hd__or2b_1 _07131_ (.A(\u_uart2wb.reg_rdata[8] ),
    .B_N(\u_uart2wb.reg_rdata[11] ),
    .X(_03069_));
 sky130_fd_sc_hd__nor2_1 _07132_ (.A(_03068_),
    .B(_03069_),
    .Y(_03070_));
 sky130_fd_sc_hd__clkbuf_2 _07133_ (.A(_02993_),
    .X(_03071_));
 sky130_fd_sc_hd__clkbuf_2 _07134_ (.A(_02981_),
    .X(_03072_));
 sky130_fd_sc_hd__a32o_1 _07135_ (.A1(_03068_),
    .A2(_03071_),
    .A3(_03069_),
    .B1(\u_uart2wb.u_msg.TxMsgBuf[73] ),
    .B2(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__a31o_1 _07136_ (.A1(_03066_),
    .A2(_03067_),
    .A3(_03070_),
    .B1(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__or3_1 _07137_ (.A(_02992_),
    .B(_02943_),
    .C(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__o21a_1 _07138_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[81] ),
    .A2(_03065_),
    .B1(_03075_),
    .X(_00421_));
 sky130_fd_sc_hd__and3b_1 _07139_ (.A_N(_03070_),
    .B(_02998_),
    .C(_03066_),
    .X(_03076_));
 sky130_fd_sc_hd__a211o_1 _07140_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[74] ),
    .A2(_02953_),
    .B1(_03051_),
    .C1(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_1 _07141_ (.A0(_03077_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[82] ),
    .S(_03053_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_1 _07142_ (.A(_03078_),
    .X(_00422_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07143_ (.A(_03044_),
    .X(_03079_));
 sky130_fd_sc_hd__and4bb_1 _07144_ (.A_N(_03068_),
    .B_N(_03066_),
    .C(_03079_),
    .D(\u_uart2wb.reg_rdata[11] ),
    .X(_03080_));
 sky130_fd_sc_hd__a211o_1 _07145_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[75] ),
    .A2(_03058_),
    .B1(_02943_),
    .C1(_03080_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_2 _07146_ (.A(_03028_),
    .X(_03082_));
 sky130_fd_sc_hd__mux2_1 _07147_ (.A0(_03081_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[83] ),
    .S(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_1 _07148_ (.A(_03083_),
    .X(_00423_));
 sky130_fd_sc_hd__a211o_1 _07149_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[76] ),
    .A2(_03058_),
    .B1(_02931_),
    .C1(_03061_),
    .X(_03084_));
 sky130_fd_sc_hd__mux2_1 _07150_ (.A0(_03084_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[84] ),
    .S(_03082_),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_1 _07151_ (.A(_03085_),
    .X(_00424_));
 sky130_fd_sc_hd__a211o_1 _07152_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[77] ),
    .A2(_03058_),
    .B1(_03051_),
    .C1(_03061_),
    .X(_03086_));
 sky130_fd_sc_hd__mux2_1 _07153_ (.A0(_03086_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[85] ),
    .S(_03082_),
    .X(_03087_));
 sky130_fd_sc_hd__clkbuf_1 _07154_ (.A(_03087_),
    .X(_00425_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07155_ (.A(_03014_),
    .X(_03088_));
 sky130_fd_sc_hd__a211o_1 _07156_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[78] ),
    .A2(_03088_),
    .B1(_03051_),
    .C1(_03060_),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_1 _07157_ (.A0(_03089_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[86] ),
    .S(_03082_),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _07158_ (.A(_03090_),
    .X(_00426_));
 sky130_fd_sc_hd__clkbuf_2 _07159_ (.A(_02937_),
    .X(_03091_));
 sky130_fd_sc_hd__o21a_1 _07160_ (.A1(\u_uart2wb.reg_rdata[17] ),
    .A2(\u_uart2wb.reg_rdata[18] ),
    .B1(\u_uart2wb.reg_rdata[19] ),
    .X(_03092_));
 sky130_fd_sc_hd__nor2_1 _07161_ (.A(_03091_),
    .B(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__inv_2 _07162_ (.A(\u_uart2wb.reg_rdata[16] ),
    .Y(_03094_));
 sky130_fd_sc_hd__a32o_1 _07163_ (.A1(_03094_),
    .A2(_03045_),
    .A3(_03092_),
    .B1(_03072_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[88] ),
    .X(_03095_));
 sky130_fd_sc_hd__a211o_1 _07164_ (.A1(\u_uart2wb.reg_rdata[16] ),
    .A2(_03093_),
    .B1(_03095_),
    .C1(_02976_),
    .X(_03096_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07165_ (.A(_03028_),
    .X(_03097_));
 sky130_fd_sc_hd__mux2_1 _07166_ (.A0(_03096_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[96] ),
    .S(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__clkbuf_1 _07167_ (.A(_03098_),
    .X(_00427_));
 sky130_fd_sc_hd__clkbuf_1 _07168_ (.A(\u_uart2wb.reg_rdata[18] ),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _07169_ (.A(\u_uart2wb.reg_rdata[17] ),
    .X(_03100_));
 sky130_fd_sc_hd__nand2_1 _07170_ (.A(_03094_),
    .B(\u_uart2wb.reg_rdata[19] ),
    .Y(_03101_));
 sky130_fd_sc_hd__nor2_1 _07171_ (.A(_03100_),
    .B(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__a32o_1 _07172_ (.A1(_03100_),
    .A2(_02998_),
    .A3(_03101_),
    .B1(\u_uart2wb.u_msg.TxMsgBuf[89] ),
    .B2(_02927_),
    .X(_03103_));
 sky130_fd_sc_hd__a31o_1 _07173_ (.A1(_03099_),
    .A2(_02947_),
    .A3(_03102_),
    .B1(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_1 _07174_ (.A0(_03104_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[97] ),
    .S(_03097_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _07175_ (.A(_03105_),
    .X(_00428_));
 sky130_fd_sc_hd__and3b_1 _07176_ (.A_N(_03102_),
    .B(_02998_),
    .C(_03099_),
    .X(_03106_));
 sky130_fd_sc_hd__a211o_1 _07177_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[90] ),
    .A2(_03088_),
    .B1(_03040_),
    .C1(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__mux2_1 _07178_ (.A0(_03107_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[98] ),
    .S(_03097_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _07179_ (.A(_03108_),
    .X(_00429_));
 sky130_fd_sc_hd__and4bb_1 _07180_ (.A_N(_03100_),
    .B_N(_03099_),
    .C(_03079_),
    .D(\u_uart2wb.reg_rdata[19] ),
    .X(_03109_));
 sky130_fd_sc_hd__a211o_1 _07181_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[91] ),
    .A2(_03088_),
    .B1(_03040_),
    .C1(_03109_),
    .X(_03110_));
 sky130_fd_sc_hd__mux2_1 _07182_ (.A0(_03110_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[99] ),
    .S(_03097_),
    .X(_03111_));
 sky130_fd_sc_hd__clkbuf_1 _07183_ (.A(_03111_),
    .X(_00430_));
 sky130_fd_sc_hd__a211o_1 _07184_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[92] ),
    .A2(_03088_),
    .B1(_02964_),
    .C1(_03093_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_1 _07185_ (.A(_02921_),
    .X(_03113_));
 sky130_fd_sc_hd__clkbuf_2 _07186_ (.A(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_1 _07187_ (.A0(_03112_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[100] ),
    .S(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__clkbuf_1 _07188_ (.A(_03115_),
    .X(_00431_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07189_ (.A(_02994_),
    .X(_03116_));
 sky130_fd_sc_hd__a211o_1 _07190_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[93] ),
    .A2(_02953_),
    .B1(_03116_),
    .C1(_03093_),
    .X(_03117_));
 sky130_fd_sc_hd__mux2_1 _07191_ (.A0(_03117_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[101] ),
    .S(_03114_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_1 _07192_ (.A(_03118_),
    .X(_00432_));
 sky130_fd_sc_hd__a221o_1 _07193_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[94] ),
    .A2(_02983_),
    .B1(_02999_),
    .B2(_03092_),
    .C1(_02942_),
    .X(_03119_));
 sky130_fd_sc_hd__mux2_1 _07194_ (.A0(_03119_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[102] ),
    .S(_03114_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_1 _07195_ (.A(_03120_),
    .X(_00433_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07196_ (.A(_02957_),
    .X(_03121_));
 sky130_fd_sc_hd__o21a_1 _07197_ (.A1(\u_uart2wb.reg_rdata[21] ),
    .A2(\u_uart2wb.reg_rdata[22] ),
    .B1(\u_uart2wb.reg_rdata[23] ),
    .X(_03122_));
 sky130_fd_sc_hd__and2_1 _07198_ (.A(_03044_),
    .B(_03122_),
    .X(_03123_));
 sky130_fd_sc_hd__nor2_1 _07199_ (.A(_03024_),
    .B(_03122_),
    .Y(_03124_));
 sky130_fd_sc_hd__mux2_1 _07200_ (.A0(_03123_),
    .A1(_03124_),
    .S(\u_uart2wb.reg_rdata[20] ),
    .X(_03125_));
 sky130_fd_sc_hd__a211o_1 _07201_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[96] ),
    .A2(_03121_),
    .B1(_02943_),
    .C1(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__mux2_1 _07202_ (.A0(_03126_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[104] ),
    .S(_03114_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_1 _07203_ (.A(_03127_),
    .X(_00434_));
 sky130_fd_sc_hd__clkbuf_1 _07204_ (.A(\u_uart2wb.reg_rdata[22] ),
    .X(_03128_));
 sky130_fd_sc_hd__clkbuf_1 _07205_ (.A(\u_uart2wb.reg_rdata[21] ),
    .X(_03129_));
 sky130_fd_sc_hd__or2b_1 _07206_ (.A(\u_uart2wb.reg_rdata[20] ),
    .B_N(\u_uart2wb.reg_rdata[23] ),
    .X(_03130_));
 sky130_fd_sc_hd__nor2_1 _07207_ (.A(_03129_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__clkbuf_2 _07208_ (.A(_02981_),
    .X(_03132_));
 sky130_fd_sc_hd__a21o_1 _07209_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[97] ),
    .A2(_03132_),
    .B1(_02962_),
    .X(_03133_));
 sky130_fd_sc_hd__a31o_1 _07210_ (.A1(_03129_),
    .A2(_02959_),
    .A3(_03130_),
    .B1(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__a31o_1 _07211_ (.A1(_03128_),
    .A2(_02960_),
    .A3(_03131_),
    .B1(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07212_ (.A(_03113_),
    .X(_03136_));
 sky130_fd_sc_hd__mux2_1 _07213_ (.A0(_03135_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[105] ),
    .S(_03136_),
    .X(_03137_));
 sky130_fd_sc_hd__clkbuf_1 _07214_ (.A(_03137_),
    .X(_00435_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07215_ (.A(_03072_),
    .X(_03138_));
 sky130_fd_sc_hd__clkbuf_2 _07216_ (.A(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__and3b_1 _07217_ (.A_N(_03131_),
    .B(_03067_),
    .C(_03128_),
    .X(_03140_));
 sky130_fd_sc_hd__a211o_1 _07218_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[98] ),
    .A2(_03139_),
    .B1(_02967_),
    .C1(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__o22a_1 _07219_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[106] ),
    .A2(_02924_),
    .B1(_02977_),
    .B2(_03141_),
    .X(_00436_));
 sky130_fd_sc_hd__and4bb_1 _07220_ (.A_N(_03129_),
    .B_N(_03128_),
    .C(_03079_),
    .D(\u_uart2wb.reg_rdata[23] ),
    .X(_03142_));
 sky130_fd_sc_hd__a211o_1 _07221_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[99] ),
    .A2(_03121_),
    .B1(_02976_),
    .C1(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__mux2_1 _07222_ (.A0(_03143_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[107] ),
    .S(_03136_),
    .X(_03144_));
 sky130_fd_sc_hd__clkbuf_1 _07223_ (.A(_03144_),
    .X(_00437_));
 sky130_fd_sc_hd__clkbuf_2 _07224_ (.A(_02962_),
    .X(_03145_));
 sky130_fd_sc_hd__a211o_1 _07225_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[100] ),
    .A2(_03121_),
    .B1(_03145_),
    .C1(_03124_),
    .X(_03146_));
 sky130_fd_sc_hd__mux2_1 _07226_ (.A0(_03146_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[108] ),
    .S(_03136_),
    .X(_03147_));
 sky130_fd_sc_hd__clkbuf_1 _07227_ (.A(_03147_),
    .X(_00438_));
 sky130_fd_sc_hd__a211o_1 _07228_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[101] ),
    .A2(_02953_),
    .B1(_03116_),
    .C1(_03124_),
    .X(_03148_));
 sky130_fd_sc_hd__mux2_1 _07229_ (.A0(_03148_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[109] ),
    .S(_03136_),
    .X(_03149_));
 sky130_fd_sc_hd__clkbuf_1 _07230_ (.A(_03149_),
    .X(_00439_));
 sky130_fd_sc_hd__a211o_1 _07231_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[102] ),
    .A2(_03121_),
    .B1(_03055_),
    .C1(_03123_),
    .X(_03150_));
 sky130_fd_sc_hd__clkbuf_2 _07232_ (.A(_03113_),
    .X(_03151_));
 sky130_fd_sc_hd__mux2_1 _07233_ (.A0(_03150_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[110] ),
    .S(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__clkbuf_1 _07234_ (.A(_03152_),
    .X(_00440_));
 sky130_fd_sc_hd__o21a_1 _07235_ (.A1(\u_uart2wb.reg_rdata[25] ),
    .A2(\u_uart2wb.reg_rdata[26] ),
    .B1(\u_uart2wb.reg_rdata[27] ),
    .X(_03153_));
 sky130_fd_sc_hd__xor2_1 _07236_ (.A(\u_uart2wb.reg_rdata[24] ),
    .B(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__a221o_1 _07237_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[104] ),
    .A2(_02997_),
    .B1(_02999_),
    .B2(_03154_),
    .C1(_02995_),
    .X(_03155_));
 sky130_fd_sc_hd__mux2_1 _07238_ (.A0(_03155_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[112] ),
    .S(_03151_),
    .X(_03156_));
 sky130_fd_sc_hd__clkbuf_1 _07239_ (.A(_03156_),
    .X(_00441_));
 sky130_fd_sc_hd__clkbuf_1 _07240_ (.A(\u_uart2wb.reg_rdata[26] ),
    .X(_03157_));
 sky130_fd_sc_hd__clkbuf_1 _07241_ (.A(\u_uart2wb.reg_rdata[25] ),
    .X(_03158_));
 sky130_fd_sc_hd__or2b_1 _07242_ (.A(\u_uart2wb.reg_rdata[24] ),
    .B_N(\u_uart2wb.reg_rdata[27] ),
    .X(_03159_));
 sky130_fd_sc_hd__nor2_1 _07243_ (.A(_03158_),
    .B(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__a32o_1 _07244_ (.A1(_03158_),
    .A2(_03071_),
    .A3(_03159_),
    .B1(\u_uart2wb.u_msg.TxMsgBuf[105] ),
    .B2(_02982_),
    .X(_03161_));
 sky130_fd_sc_hd__a31o_1 _07245_ (.A1(_03157_),
    .A2(_03067_),
    .A3(_03160_),
    .B1(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__or3_1 _07246_ (.A(_02949_),
    .B(_02976_),
    .C(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__o21a_1 _07247_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[113] ),
    .A2(_03065_),
    .B1(_03163_),
    .X(_00442_));
 sky130_fd_sc_hd__and3b_1 _07248_ (.A_N(_03160_),
    .B(_03038_),
    .C(_03157_),
    .X(_03164_));
 sky130_fd_sc_hd__a211o_1 _07249_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[106] ),
    .A2(_02997_),
    .B1(_03116_),
    .C1(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__mux2_1 _07250_ (.A0(_03165_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[114] ),
    .S(_03151_),
    .X(_03166_));
 sky130_fd_sc_hd__clkbuf_1 _07251_ (.A(_03166_),
    .X(_00443_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07252_ (.A(_02957_),
    .X(_03167_));
 sky130_fd_sc_hd__and4bb_1 _07253_ (.A_N(_03158_),
    .B_N(_03157_),
    .C(_03079_),
    .D(\u_uart2wb.reg_rdata[27] ),
    .X(_03168_));
 sky130_fd_sc_hd__a211o_1 _07254_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[107] ),
    .A2(_03167_),
    .B1(_02955_),
    .C1(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__mux2_1 _07255_ (.A0(_03169_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[115] ),
    .S(_03151_),
    .X(_03170_));
 sky130_fd_sc_hd__clkbuf_1 _07256_ (.A(_03170_),
    .X(_00444_));
 sky130_fd_sc_hd__nor2_1 _07257_ (.A(_03091_),
    .B(_03153_),
    .Y(_03171_));
 sky130_fd_sc_hd__a211o_1 _07258_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[108] ),
    .A2(_02971_),
    .B1(_02969_),
    .C1(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__o21a_1 _07259_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[116] ),
    .A2(_03065_),
    .B1(_03172_),
    .X(_00445_));
 sky130_fd_sc_hd__a211o_1 _07260_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[109] ),
    .A2(_03167_),
    .B1(_03116_),
    .C1(_03171_),
    .X(_03173_));
 sky130_fd_sc_hd__clkbuf_2 _07261_ (.A(_03113_),
    .X(_03174_));
 sky130_fd_sc_hd__mux2_1 _07262_ (.A0(_03173_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[117] ),
    .S(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__clkbuf_1 _07263_ (.A(_03175_),
    .X(_00446_));
 sky130_fd_sc_hd__a221o_1 _07264_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[110] ),
    .A2(_02997_),
    .B1(_02999_),
    .B2(_03153_),
    .C1(_02995_),
    .X(_03176_));
 sky130_fd_sc_hd__mux2_1 _07265_ (.A0(_03176_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[118] ),
    .S(_03174_),
    .X(_03177_));
 sky130_fd_sc_hd__clkbuf_1 _07266_ (.A(_03177_),
    .X(_00447_));
 sky130_fd_sc_hd__o22a_1 _07267_ (.A1(_02156_),
    .A2(\u_spi2wb.reg_be[0] ),
    .B1(_02157_),
    .B2(wbm_sel_i[0]),
    .X(_03178_));
 sky130_fd_sc_hd__clkbuf_1 _07268_ (.A(_03178_),
    .X(_03179_));
 sky130_fd_sc_hd__mux2_1 _07269_ (.A0(_03179_),
    .A1(\u_async_wb.u_cmd_if.mem[3][0] ),
    .S(_02809_),
    .X(_03180_));
 sky130_fd_sc_hd__clkbuf_1 _07270_ (.A(_03180_),
    .X(_00448_));
 sky130_fd_sc_hd__clkbuf_1 _07271_ (.A(_02158_),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_1 _07272_ (.A0(_03181_),
    .A1(\u_async_wb.u_cmd_if.mem[3][1] ),
    .S(_02809_),
    .X(_03182_));
 sky130_fd_sc_hd__clkbuf_1 _07273_ (.A(_03182_),
    .X(_00449_));
 sky130_fd_sc_hd__clkbuf_1 _07274_ (.A(_02415_),
    .X(_03183_));
 sky130_fd_sc_hd__mux2_1 _07275_ (.A0(_03183_),
    .A1(\u_async_wb.u_cmd_if.mem[3][2] ),
    .S(_02809_),
    .X(_03184_));
 sky130_fd_sc_hd__clkbuf_1 _07276_ (.A(_03184_),
    .X(_00450_));
 sky130_fd_sc_hd__o22a_2 _07277_ (.A1(_02156_),
    .A2(\u_spi2wb.reg_be[3] ),
    .B1(wbm_sel_i[3]),
    .B2(_02157_),
    .X(_03185_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07278_ (.A(_02808_),
    .X(_03186_));
 sky130_fd_sc_hd__mux2_1 _07279_ (.A0(_03185_),
    .A1(\u_async_wb.u_cmd_if.mem[3][3] ),
    .S(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__clkbuf_1 _07280_ (.A(_03187_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _07281_ (.A0(_02286_),
    .A1(\u_async_wb.u_cmd_if.mem[3][4] ),
    .S(_03186_),
    .X(_03188_));
 sky130_fd_sc_hd__clkbuf_1 _07282_ (.A(_03188_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _07283_ (.A0(_02266_),
    .A1(\u_async_wb.u_cmd_if.mem[3][5] ),
    .S(_03186_),
    .X(_03189_));
 sky130_fd_sc_hd__clkbuf_1 _07284_ (.A(_03189_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _07285_ (.A0(_02259_),
    .A1(\u_async_wb.u_cmd_if.mem[3][6] ),
    .S(_03186_),
    .X(_03190_));
 sky130_fd_sc_hd__clkbuf_1 _07286_ (.A(_03190_),
    .X(_00454_));
 sky130_fd_sc_hd__clkbuf_2 _07287_ (.A(_02807_),
    .X(_03191_));
 sky130_fd_sc_hd__clkbuf_2 _07288_ (.A(_03191_),
    .X(_03192_));
 sky130_fd_sc_hd__clkbuf_2 _07289_ (.A(_03192_),
    .X(_03193_));
 sky130_fd_sc_hd__mux2_1 _07290_ (.A0(_02254_),
    .A1(\u_async_wb.u_cmd_if.mem[3][7] ),
    .S(_03193_),
    .X(_03194_));
 sky130_fd_sc_hd__clkbuf_1 _07291_ (.A(_03194_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _07292_ (.A0(_02246_),
    .A1(\u_async_wb.u_cmd_if.mem[3][8] ),
    .S(_03193_),
    .X(_03195_));
 sky130_fd_sc_hd__clkbuf_1 _07293_ (.A(_03195_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _07294_ (.A0(_02239_),
    .A1(\u_async_wb.u_cmd_if.mem[3][9] ),
    .S(_03193_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_1 _07295_ (.A(_03196_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _07296_ (.A0(_02473_),
    .A1(\u_async_wb.u_cmd_if.mem[3][10] ),
    .S(_03193_),
    .X(_03197_));
 sky130_fd_sc_hd__clkbuf_1 _07297_ (.A(_03197_),
    .X(_00458_));
 sky130_fd_sc_hd__clkbuf_2 _07298_ (.A(_03192_),
    .X(_03198_));
 sky130_fd_sc_hd__mux2_1 _07299_ (.A0(_02228_),
    .A1(\u_async_wb.u_cmd_if.mem[3][11] ),
    .S(_03198_),
    .X(_03199_));
 sky130_fd_sc_hd__clkbuf_1 _07300_ (.A(_03199_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _07301_ (.A0(_02477_),
    .A1(\u_async_wb.u_cmd_if.mem[3][12] ),
    .S(_03198_),
    .X(_03200_));
 sky130_fd_sc_hd__clkbuf_1 _07302_ (.A(_03200_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _07303_ (.A0(_02181_),
    .A1(\u_async_wb.u_cmd_if.mem[3][13] ),
    .S(_03198_),
    .X(_03201_));
 sky130_fd_sc_hd__clkbuf_1 _07304_ (.A(_03201_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _07305_ (.A0(_02187_),
    .A1(\u_async_wb.u_cmd_if.mem[3][14] ),
    .S(_03198_),
    .X(_03202_));
 sky130_fd_sc_hd__clkbuf_1 _07306_ (.A(_03202_),
    .X(_00462_));
 sky130_fd_sc_hd__clkbuf_2 _07307_ (.A(_03192_),
    .X(_03203_));
 sky130_fd_sc_hd__mux2_1 _07308_ (.A0(_02485_),
    .A1(\u_async_wb.u_cmd_if.mem[3][15] ),
    .S(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__clkbuf_1 _07309_ (.A(_03204_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _07310_ (.A0(_02200_),
    .A1(\u_async_wb.u_cmd_if.mem[3][16] ),
    .S(_03203_),
    .X(_03205_));
 sky130_fd_sc_hd__clkbuf_1 _07311_ (.A(_03205_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _07312_ (.A0(_02206_),
    .A1(\u_async_wb.u_cmd_if.mem[3][17] ),
    .S(_03203_),
    .X(_03206_));
 sky130_fd_sc_hd__clkbuf_1 _07313_ (.A(_03206_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _07314_ (.A0(_02211_),
    .A1(\u_async_wb.u_cmd_if.mem[3][18] ),
    .S(_03203_),
    .X(_03207_));
 sky130_fd_sc_hd__clkbuf_1 _07315_ (.A(_03207_),
    .X(_00466_));
 sky130_fd_sc_hd__clkbuf_2 _07316_ (.A(_03192_),
    .X(_03208_));
 sky130_fd_sc_hd__mux2_1 _07317_ (.A0(_02493_),
    .A1(\u_async_wb.u_cmd_if.mem[3][19] ),
    .S(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__clkbuf_1 _07318_ (.A(_03209_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _07319_ (.A0(_02413_),
    .A1(\u_async_wb.u_cmd_if.mem[3][20] ),
    .S(_03208_),
    .X(_03210_));
 sky130_fd_sc_hd__clkbuf_1 _07320_ (.A(_03210_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _07321_ (.A0(_02424_),
    .A1(\u_async_wb.u_cmd_if.mem[3][21] ),
    .S(_03208_),
    .X(_03211_));
 sky130_fd_sc_hd__clkbuf_1 _07322_ (.A(_03211_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _07323_ (.A0(_02427_),
    .A1(\u_async_wb.u_cmd_if.mem[3][22] ),
    .S(_03208_),
    .X(_03212_));
 sky130_fd_sc_hd__clkbuf_1 _07324_ (.A(_03212_),
    .X(_00470_));
 sky130_fd_sc_hd__clkbuf_1 _07325_ (.A(_02807_),
    .X(_03213_));
 sky130_fd_sc_hd__clkbuf_2 _07326_ (.A(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__mux2_1 _07327_ (.A0(_02430_),
    .A1(\u_async_wb.u_cmd_if.mem[3][23] ),
    .S(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_1 _07328_ (.A(_03215_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _07329_ (.A0(_02433_),
    .A1(\u_async_wb.u_cmd_if.mem[3][24] ),
    .S(_03214_),
    .X(_03216_));
 sky130_fd_sc_hd__clkbuf_1 _07330_ (.A(_03216_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _07331_ (.A0(_02439_),
    .A1(\u_async_wb.u_cmd_if.mem[3][25] ),
    .S(_03214_),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_1 _07332_ (.A(_03217_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _07333_ (.A0(_02442_),
    .A1(\u_async_wb.u_cmd_if.mem[3][26] ),
    .S(_03214_),
    .X(_03218_));
 sky130_fd_sc_hd__clkbuf_1 _07334_ (.A(_03218_),
    .X(_00474_));
 sky130_fd_sc_hd__clkbuf_2 _07335_ (.A(_03213_),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_1 _07336_ (.A0(_02445_),
    .A1(\u_async_wb.u_cmd_if.mem[3][27] ),
    .S(_03219_),
    .X(_03220_));
 sky130_fd_sc_hd__clkbuf_1 _07337_ (.A(_03220_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _07338_ (.A0(_02513_),
    .A1(\u_async_wb.u_cmd_if.mem[3][28] ),
    .S(_03219_),
    .X(_03221_));
 sky130_fd_sc_hd__clkbuf_1 _07339_ (.A(_03221_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _07340_ (.A0(_02515_),
    .A1(\u_async_wb.u_cmd_if.mem[3][29] ),
    .S(_03219_),
    .X(_03222_));
 sky130_fd_sc_hd__clkbuf_1 _07341_ (.A(_03222_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _07342_ (.A0(_02521_),
    .A1(\u_async_wb.u_cmd_if.mem[3][30] ),
    .S(_03219_),
    .X(_03223_));
 sky130_fd_sc_hd__clkbuf_1 _07343_ (.A(_03223_),
    .X(_00478_));
 sky130_fd_sc_hd__clkbuf_2 _07344_ (.A(_03213_),
    .X(_03224_));
 sky130_fd_sc_hd__mux2_1 _07345_ (.A0(_02733_),
    .A1(\u_async_wb.u_cmd_if.mem[3][31] ),
    .S(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__clkbuf_1 _07346_ (.A(_03225_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _07347_ (.A0(_02525_),
    .A1(\u_async_wb.u_cmd_if.mem[3][32] ),
    .S(_03224_),
    .X(_03226_));
 sky130_fd_sc_hd__clkbuf_1 _07348_ (.A(_03226_),
    .X(_00480_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07349_ (.A(_02399_),
    .X(_03227_));
 sky130_fd_sc_hd__mux2_1 _07350_ (.A0(_03227_),
    .A1(\u_async_wb.u_cmd_if.mem[3][33] ),
    .S(_03224_),
    .X(_03228_));
 sky130_fd_sc_hd__clkbuf_1 _07351_ (.A(_03228_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _07352_ (.A0(_02529_),
    .A1(\u_async_wb.u_cmd_if.mem[3][34] ),
    .S(_03224_),
    .X(_03229_));
 sky130_fd_sc_hd__clkbuf_1 _07353_ (.A(_03229_),
    .X(_00482_));
 sky130_fd_sc_hd__clkbuf_2 _07354_ (.A(_03213_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _07355_ (.A0(_02531_),
    .A1(\u_async_wb.u_cmd_if.mem[3][35] ),
    .S(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__clkbuf_1 _07356_ (.A(_03231_),
    .X(_00483_));
 sky130_fd_sc_hd__clkbuf_1 _07357_ (.A(_01485_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_1 _07358_ (.A0(_03232_),
    .A1(\u_async_wb.u_cmd_if.mem[3][36] ),
    .S(_03230_),
    .X(_03233_));
 sky130_fd_sc_hd__clkbuf_1 _07359_ (.A(_03233_),
    .X(_00484_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07360_ (.A(_02372_),
    .X(_03234_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07361_ (.A(_01730_),
    .X(_03235_));
 sky130_fd_sc_hd__and2_1 _07362_ (.A(_03235_),
    .B(\u_spi2wb.reg_addr[0] ),
    .X(_03236_));
 sky130_fd_sc_hd__a221o_4 _07363_ (.A1(wbm_adr_i[0]),
    .A2(_01776_),
    .B1(_03234_),
    .B2(\u_uart2wb.reg_addr[0] ),
    .C1(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__mux2_1 _07364_ (.A0(_03237_),
    .A1(\u_async_wb.u_cmd_if.mem[3][37] ),
    .S(_03230_),
    .X(_03238_));
 sky130_fd_sc_hd__clkbuf_1 _07365_ (.A(_03238_),
    .X(_00485_));
 sky130_fd_sc_hd__clkbuf_1 _07366_ (.A(_01730_),
    .X(_03239_));
 sky130_fd_sc_hd__and2_1 _07367_ (.A(_03239_),
    .B(\u_spi2wb.reg_addr[1] ),
    .X(_03240_));
 sky130_fd_sc_hd__a221o_4 _07368_ (.A1(wbm_adr_i[1]),
    .A2(_01776_),
    .B1(_03234_),
    .B2(\u_uart2wb.reg_addr[1] ),
    .C1(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__mux2_1 _07369_ (.A0(_03241_),
    .A1(\u_async_wb.u_cmd_if.mem[3][38] ),
    .S(_03230_),
    .X(_03242_));
 sky130_fd_sc_hd__clkbuf_1 _07370_ (.A(_03242_),
    .X(_00486_));
 sky130_fd_sc_hd__clkbuf_1 _07371_ (.A(_02162_),
    .X(_03243_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07372_ (.A(_02807_),
    .X(_03244_));
 sky130_fd_sc_hd__clkbuf_2 _07373_ (.A(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_1 _07374_ (.A0(_03243_),
    .A1(\u_async_wb.u_cmd_if.mem[3][39] ),
    .S(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__clkbuf_1 _07375_ (.A(_03246_),
    .X(_00487_));
 sky130_fd_sc_hd__clkbuf_1 _07376_ (.A(_02165_),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_1 _07377_ (.A0(_03247_),
    .A1(\u_async_wb.u_cmd_if.mem[3][40] ),
    .S(_03245_),
    .X(_03248_));
 sky130_fd_sc_hd__clkbuf_1 _07378_ (.A(_03248_),
    .X(_00488_));
 sky130_fd_sc_hd__clkbuf_1 _07379_ (.A(_02168_),
    .X(_03249_));
 sky130_fd_sc_hd__mux2_1 _07380_ (.A0(_03249_),
    .A1(\u_async_wb.u_cmd_if.mem[3][41] ),
    .S(_03245_),
    .X(_03250_));
 sky130_fd_sc_hd__clkbuf_1 _07381_ (.A(_03250_),
    .X(_00489_));
 sky130_fd_sc_hd__clkbuf_1 _07382_ (.A(_01775_),
    .X(_03251_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07383_ (.A(_02372_),
    .X(_03252_));
 sky130_fd_sc_hd__and2_1 _07384_ (.A(_03239_),
    .B(\u_spi2wb.reg_addr[5] ),
    .X(_03253_));
 sky130_fd_sc_hd__a221o_2 _07385_ (.A1(wbm_adr_i[5]),
    .A2(_03251_),
    .B1(_03252_),
    .B2(\u_uart2wb.reg_addr[5] ),
    .C1(_03253_),
    .X(_03254_));
 sky130_fd_sc_hd__mux2_1 _07386_ (.A0(_03254_),
    .A1(\u_async_wb.u_cmd_if.mem[3][42] ),
    .S(_03245_),
    .X(_03255_));
 sky130_fd_sc_hd__clkbuf_1 _07387_ (.A(_03255_),
    .X(_00490_));
 sky130_fd_sc_hd__and2_1 _07388_ (.A(_03239_),
    .B(\u_spi2wb.reg_addr[6] ),
    .X(_03256_));
 sky130_fd_sc_hd__a221o_2 _07389_ (.A1(wbm_adr_i[6]),
    .A2(_03251_),
    .B1(_03252_),
    .B2(\u_uart2wb.reg_addr[6] ),
    .C1(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__clkbuf_2 _07390_ (.A(_03244_),
    .X(_03258_));
 sky130_fd_sc_hd__mux2_1 _07391_ (.A0(_03257_),
    .A1(\u_async_wb.u_cmd_if.mem[3][43] ),
    .S(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__clkbuf_1 _07392_ (.A(_03259_),
    .X(_00491_));
 sky130_fd_sc_hd__and2_1 _07393_ (.A(_03239_),
    .B(\u_spi2wb.reg_addr[7] ),
    .X(_03260_));
 sky130_fd_sc_hd__a221o_2 _07394_ (.A1(wbm_adr_i[7]),
    .A2(_03251_),
    .B1(_03252_),
    .B2(\u_uart2wb.reg_addr[7] ),
    .C1(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__mux2_1 _07395_ (.A0(_03261_),
    .A1(\u_async_wb.u_cmd_if.mem[3][44] ),
    .S(_03258_),
    .X(_03262_));
 sky130_fd_sc_hd__clkbuf_1 _07396_ (.A(_03262_),
    .X(_00492_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07397_ (.A(_02250_),
    .X(_03263_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07398_ (.A(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__clkbuf_1 _07399_ (.A(_01736_),
    .X(_03265_));
 sky130_fd_sc_hd__a22o_1 _07400_ (.A1(_01731_),
    .A2(\u_spi2wb.reg_addr[8] ),
    .B1(wbm_adr_i[8]),
    .B2(_03265_),
    .X(_03266_));
 sky130_fd_sc_hd__a21o_1 _07401_ (.A1(\u_uart2wb.reg_addr[8] ),
    .A2(_03264_),
    .B1(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__mux2_1 _07402_ (.A0(_03267_),
    .A1(\u_async_wb.u_cmd_if.mem[3][45] ),
    .S(_03258_),
    .X(_03268_));
 sky130_fd_sc_hd__clkbuf_1 _07403_ (.A(_03268_),
    .X(_00493_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07404_ (.A(_02349_),
    .X(_03269_));
 sky130_fd_sc_hd__and2_1 _07405_ (.A(_03269_),
    .B(\u_spi2wb.reg_addr[9] ),
    .X(_03270_));
 sky130_fd_sc_hd__a221o_2 _07406_ (.A1(wbm_adr_i[9]),
    .A2(_03251_),
    .B1(_03252_),
    .B2(\u_uart2wb.reg_addr[9] ),
    .C1(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__mux2_1 _07407_ (.A0(_03271_),
    .A1(\u_async_wb.u_cmd_if.mem[3][46] ),
    .S(_03258_),
    .X(_03272_));
 sky130_fd_sc_hd__clkbuf_1 _07408_ (.A(_03272_),
    .X(_00494_));
 sky130_fd_sc_hd__clkbuf_1 _07409_ (.A(_03269_),
    .X(_03273_));
 sky130_fd_sc_hd__a22o_1 _07410_ (.A1(_03273_),
    .A2(\u_spi2wb.reg_addr[10] ),
    .B1(wbm_adr_i[10]),
    .B2(_03265_),
    .X(_03274_));
 sky130_fd_sc_hd__a21o_1 _07411_ (.A1(\u_uart2wb.reg_addr[10] ),
    .A2(_03264_),
    .B1(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__clkbuf_2 _07412_ (.A(_03244_),
    .X(_03276_));
 sky130_fd_sc_hd__mux2_1 _07413_ (.A0(_03275_),
    .A1(\u_async_wb.u_cmd_if.mem[3][47] ),
    .S(_03276_),
    .X(_03277_));
 sky130_fd_sc_hd__clkbuf_1 _07414_ (.A(_03277_),
    .X(_00495_));
 sky130_fd_sc_hd__a22o_1 _07415_ (.A1(_03273_),
    .A2(\u_spi2wb.reg_addr[11] ),
    .B1(wbm_adr_i[11]),
    .B2(_03265_),
    .X(_03278_));
 sky130_fd_sc_hd__a21o_1 _07416_ (.A1(\u_uart2wb.reg_addr[11] ),
    .A2(_03264_),
    .B1(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__mux2_1 _07417_ (.A0(_03279_),
    .A1(\u_async_wb.u_cmd_if.mem[3][48] ),
    .S(_03276_),
    .X(_03280_));
 sky130_fd_sc_hd__clkbuf_1 _07418_ (.A(_03280_),
    .X(_00496_));
 sky130_fd_sc_hd__clkbuf_1 _07419_ (.A(_03263_),
    .X(_03281_));
 sky130_fd_sc_hd__a22o_1 _07420_ (.A1(_03273_),
    .A2(\u_spi2wb.reg_addr[12] ),
    .B1(wbm_adr_i[12]),
    .B2(_03265_),
    .X(_03282_));
 sky130_fd_sc_hd__a21o_1 _07421_ (.A1(\u_uart2wb.reg_addr[12] ),
    .A2(_03281_),
    .B1(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__mux2_1 _07422_ (.A0(_03283_),
    .A1(\u_async_wb.u_cmd_if.mem[3][49] ),
    .S(_03276_),
    .X(_03284_));
 sky130_fd_sc_hd__clkbuf_1 _07423_ (.A(_03284_),
    .X(_00497_));
 sky130_fd_sc_hd__clkbuf_1 _07424_ (.A(_01736_),
    .X(_03285_));
 sky130_fd_sc_hd__a22o_1 _07425_ (.A1(_03273_),
    .A2(\u_spi2wb.reg_addr[13] ),
    .B1(wbm_adr_i[13]),
    .B2(_03285_),
    .X(_03286_));
 sky130_fd_sc_hd__a21o_2 _07426_ (.A1(\u_uart2wb.reg_addr[13] ),
    .A2(_03281_),
    .B1(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__mux2_1 _07427_ (.A0(_03287_),
    .A1(\u_async_wb.u_cmd_if.mem[3][50] ),
    .S(_03276_),
    .X(_03288_));
 sky130_fd_sc_hd__clkbuf_1 _07428_ (.A(_03288_),
    .X(_00498_));
 sky130_fd_sc_hd__and2_1 _07429_ (.A(_03269_),
    .B(\u_spi2wb.reg_addr[14] ),
    .X(_03289_));
 sky130_fd_sc_hd__a221o_2 _07430_ (.A1(wbm_adr_i[14]),
    .A2(_01741_),
    .B1(_03263_),
    .B2(\u_uart2wb.reg_addr[14] ),
    .C1(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__clkbuf_2 _07431_ (.A(_03244_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _07432_ (.A0(_03290_),
    .A1(\u_async_wb.u_cmd_if.mem[3][51] ),
    .S(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__clkbuf_1 _07433_ (.A(_03292_),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_1 _07434_ (.A1(_03235_),
    .A2(\u_spi2wb.reg_addr[15] ),
    .B1(wbm_adr_i[15]),
    .B2(_03285_),
    .X(_03293_));
 sky130_fd_sc_hd__a21o_2 _07435_ (.A1(\u_uart2wb.reg_addr[15] ),
    .A2(_03281_),
    .B1(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__mux2_1 _07436_ (.A0(_03294_),
    .A1(\u_async_wb.u_cmd_if.mem[3][52] ),
    .S(_03291_),
    .X(_03295_));
 sky130_fd_sc_hd__clkbuf_1 _07437_ (.A(_03295_),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _07438_ (.A1(_03235_),
    .A2(\u_spi2wb.reg_addr[16] ),
    .B1(wbm_adr_i[16]),
    .B2(_03285_),
    .X(_03296_));
 sky130_fd_sc_hd__a21o_2 _07439_ (.A1(\u_uart2wb.reg_addr[16] ),
    .A2(_03281_),
    .B1(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__mux2_1 _07440_ (.A0(_03297_),
    .A1(\u_async_wb.u_cmd_if.mem[3][53] ),
    .S(_03291_),
    .X(_03298_));
 sky130_fd_sc_hd__clkbuf_1 _07441_ (.A(_03298_),
    .X(_00501_));
 sky130_fd_sc_hd__and2_1 _07442_ (.A(_03269_),
    .B(\u_spi2wb.reg_addr[17] ),
    .X(_03299_));
 sky130_fd_sc_hd__a221o_2 _07443_ (.A1(wbm_adr_i[17]),
    .A2(_01741_),
    .B1(_03263_),
    .B2(\u_uart2wb.reg_addr[17] ),
    .C1(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__mux2_1 _07444_ (.A0(_03300_),
    .A1(\u_async_wb.u_cmd_if.mem[3][54] ),
    .S(_03291_),
    .X(_03301_));
 sky130_fd_sc_hd__clkbuf_1 _07445_ (.A(_03301_),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _07446_ (.A1(_03235_),
    .A2(\u_spi2wb.reg_addr[18] ),
    .B1(wbm_adr_i[18]),
    .B2(_03285_),
    .X(_03302_));
 sky130_fd_sc_hd__a21o_2 _07447_ (.A1(\u_uart2wb.reg_addr[18] ),
    .A2(_03234_),
    .B1(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07448_ (.A(_03191_),
    .X(_03304_));
 sky130_fd_sc_hd__mux2_1 _07449_ (.A0(_03303_),
    .A1(\u_async_wb.u_cmd_if.mem[3][55] ),
    .S(_03304_),
    .X(_03305_));
 sky130_fd_sc_hd__clkbuf_1 _07450_ (.A(_03305_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _07451_ (.A0(_02249_),
    .A1(\u_async_wb.u_cmd_if.mem[3][56] ),
    .S(_03304_),
    .X(_03306_));
 sky130_fd_sc_hd__clkbuf_1 _07452_ (.A(_03306_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _07453_ (.A0(_02241_),
    .A1(\u_async_wb.u_cmd_if.mem[3][57] ),
    .S(_03304_),
    .X(_03307_));
 sky130_fd_sc_hd__clkbuf_1 _07454_ (.A(_03307_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _07455_ (.A0(_02235_),
    .A1(\u_async_wb.u_cmd_if.mem[3][58] ),
    .S(_03304_),
    .X(_03308_));
 sky130_fd_sc_hd__clkbuf_1 _07456_ (.A(_03308_),
    .X(_00506_));
 sky130_fd_sc_hd__clkbuf_2 _07457_ (.A(_03191_),
    .X(_03309_));
 sky130_fd_sc_hd__mux2_1 _07458_ (.A0(_02230_),
    .A1(\u_async_wb.u_cmd_if.mem[3][59] ),
    .S(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__clkbuf_1 _07459_ (.A(_03310_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _07460_ (.A0(_02224_),
    .A1(\u_async_wb.u_cmd_if.mem[3][60] ),
    .S(_03309_),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_1 _07461_ (.A(_03311_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _07462_ (.A0(_02218_),
    .A1(\u_async_wb.u_cmd_if.mem[3][61] ),
    .S(_03309_),
    .X(_03312_));
 sky130_fd_sc_hd__clkbuf_1 _07463_ (.A(_03312_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _07464_ (.A0(_02410_),
    .A1(\u_async_wb.u_cmd_if.mem[3][62] ),
    .S(_03309_),
    .X(_03313_));
 sky130_fd_sc_hd__clkbuf_1 _07465_ (.A(_03313_),
    .X(_00510_));
 sky130_fd_sc_hd__clkbuf_2 _07466_ (.A(_03191_),
    .X(_03314_));
 sky130_fd_sc_hd__mux2_1 _07467_ (.A0(_02280_),
    .A1(\u_async_wb.u_cmd_if.mem[3][63] ),
    .S(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__clkbuf_1 _07468_ (.A(_03315_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _07469_ (.A0(_02277_),
    .A1(\u_async_wb.u_cmd_if.mem[3][64] ),
    .S(_03314_),
    .X(_03316_));
 sky130_fd_sc_hd__clkbuf_1 _07470_ (.A(_03316_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _07471_ (.A0(_02275_),
    .A1(\u_async_wb.u_cmd_if.mem[3][65] ),
    .S(_03314_),
    .X(_03317_));
 sky130_fd_sc_hd__clkbuf_1 _07472_ (.A(_03317_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _07473_ (.A0(_02273_),
    .A1(\u_async_wb.u_cmd_if.mem[3][66] ),
    .S(_03314_),
    .X(_03318_));
 sky130_fd_sc_hd__clkbuf_1 _07474_ (.A(_03318_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _07475_ (.A0(_02271_),
    .A1(\u_async_wb.u_cmd_if.mem[3][67] ),
    .S(_02808_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_1 _07476_ (.A(_03319_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _07477_ (.A0(_02268_),
    .A1(\u_async_wb.u_cmd_if.mem[3][68] ),
    .S(_02808_),
    .X(_03320_));
 sky130_fd_sc_hd__clkbuf_1 _07478_ (.A(_03320_),
    .X(_00516_));
 sky130_fd_sc_hd__and3b_1 _07479_ (.A_N(_01489_),
    .B(_02798_),
    .C(_01501_),
    .X(_03321_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07480_ (.A(_03321_),
    .X(_03322_));
 sky130_fd_sc_hd__clkbuf_2 _07481_ (.A(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__mux2_1 _07482_ (.A0(\u_async_wb.u_cmd_if.mem[2][0] ),
    .A1(_03179_),
    .S(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__clkbuf_1 _07483_ (.A(_03324_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _07484_ (.A0(\u_async_wb.u_cmd_if.mem[2][1] ),
    .A1(_03181_),
    .S(_03323_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_1 _07485_ (.A(_03325_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _07486_ (.A0(\u_async_wb.u_cmd_if.mem[2][2] ),
    .A1(_03183_),
    .S(_03323_),
    .X(_03326_));
 sky130_fd_sc_hd__clkbuf_1 _07487_ (.A(_03326_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _07488_ (.A0(\u_async_wb.u_cmd_if.mem[2][3] ),
    .A1(_03185_),
    .S(_03323_),
    .X(_03327_));
 sky130_fd_sc_hd__clkbuf_1 _07489_ (.A(_03327_),
    .X(_00520_));
 sky130_fd_sc_hd__clkbuf_2 _07490_ (.A(_03322_),
    .X(_03328_));
 sky130_fd_sc_hd__mux2_1 _07491_ (.A0(\u_async_wb.u_cmd_if.mem[2][4] ),
    .A1(_02285_),
    .S(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__clkbuf_1 _07492_ (.A(_03329_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _07493_ (.A0(\u_async_wb.u_cmd_if.mem[2][5] ),
    .A1(_02265_),
    .S(_03328_),
    .X(_03330_));
 sky130_fd_sc_hd__clkbuf_1 _07494_ (.A(_03330_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _07495_ (.A0(\u_async_wb.u_cmd_if.mem[2][6] ),
    .A1(_02258_),
    .S(_03328_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_1 _07496_ (.A(_03331_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _07497_ (.A0(\u_async_wb.u_cmd_if.mem[2][7] ),
    .A1(_02253_),
    .S(_03328_),
    .X(_03332_));
 sky130_fd_sc_hd__clkbuf_1 _07498_ (.A(_03332_),
    .X(_00524_));
 sky130_fd_sc_hd__clkbuf_2 _07499_ (.A(_03322_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _07500_ (.A0(\u_async_wb.u_cmd_if.mem[2][8] ),
    .A1(_02245_),
    .S(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__clkbuf_1 _07501_ (.A(_03334_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _07502_ (.A0(\u_async_wb.u_cmd_if.mem[2][9] ),
    .A1(_02239_),
    .S(_03333_),
    .X(_03335_));
 sky130_fd_sc_hd__clkbuf_1 _07503_ (.A(_03335_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _07504_ (.A0(\u_async_wb.u_cmd_if.mem[2][10] ),
    .A1(_02233_),
    .S(_03333_),
    .X(_03336_));
 sky130_fd_sc_hd__clkbuf_1 _07505_ (.A(_03336_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _07506_ (.A0(\u_async_wb.u_cmd_if.mem[2][11] ),
    .A1(_02227_),
    .S(_03333_),
    .X(_03337_));
 sky130_fd_sc_hd__clkbuf_1 _07507_ (.A(_03337_),
    .X(_00528_));
 sky130_fd_sc_hd__clkbuf_2 _07508_ (.A(_03321_),
    .X(_03338_));
 sky130_fd_sc_hd__clkbuf_2 _07509_ (.A(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__clkbuf_2 _07510_ (.A(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__mux2_1 _07511_ (.A0(\u_async_wb.u_cmd_if.mem[2][12] ),
    .A1(_02154_),
    .S(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__clkbuf_1 _07512_ (.A(_03341_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _07513_ (.A0(\u_async_wb.u_cmd_if.mem[2][13] ),
    .A1(_02180_),
    .S(_03340_),
    .X(_03342_));
 sky130_fd_sc_hd__clkbuf_1 _07514_ (.A(_03342_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _07515_ (.A0(\u_async_wb.u_cmd_if.mem[2][14] ),
    .A1(_02186_),
    .S(_03340_),
    .X(_03343_));
 sky130_fd_sc_hd__clkbuf_1 _07516_ (.A(_03343_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _07517_ (.A0(\u_async_wb.u_cmd_if.mem[2][15] ),
    .A1(_02191_),
    .S(_03340_),
    .X(_03344_));
 sky130_fd_sc_hd__clkbuf_1 _07518_ (.A(_03344_),
    .X(_00532_));
 sky130_fd_sc_hd__clkbuf_2 _07519_ (.A(_03339_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _07520_ (.A0(\u_async_wb.u_cmd_if.mem[2][16] ),
    .A1(_02199_),
    .S(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__clkbuf_1 _07521_ (.A(_03346_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _07522_ (.A0(\u_async_wb.u_cmd_if.mem[2][17] ),
    .A1(_02205_),
    .S(_03345_),
    .X(_03347_));
 sky130_fd_sc_hd__clkbuf_1 _07523_ (.A(_03347_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _07524_ (.A0(\u_async_wb.u_cmd_if.mem[2][18] ),
    .A1(_02210_),
    .S(_03345_),
    .X(_03348_));
 sky130_fd_sc_hd__clkbuf_1 _07525_ (.A(_03348_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _07526_ (.A0(\u_async_wb.u_cmd_if.mem[2][19] ),
    .A1(_02216_),
    .S(_03345_),
    .X(_03349_));
 sky130_fd_sc_hd__clkbuf_1 _07527_ (.A(_03349_),
    .X(_00536_));
 sky130_fd_sc_hd__clkbuf_2 _07528_ (.A(_03339_),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_1 _07529_ (.A0(\u_async_wb.u_cmd_if.mem[2][20] ),
    .A1(_02412_),
    .S(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_1 _07530_ (.A(_03351_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _07531_ (.A0(\u_async_wb.u_cmd_if.mem[2][21] ),
    .A1(_02423_),
    .S(_03350_),
    .X(_03352_));
 sky130_fd_sc_hd__clkbuf_1 _07532_ (.A(_03352_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _07533_ (.A0(\u_async_wb.u_cmd_if.mem[2][22] ),
    .A1(_02426_),
    .S(_03350_),
    .X(_03353_));
 sky130_fd_sc_hd__clkbuf_1 _07534_ (.A(_03353_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _07535_ (.A0(\u_async_wb.u_cmd_if.mem[2][23] ),
    .A1(_02429_),
    .S(_03350_),
    .X(_03354_));
 sky130_fd_sc_hd__clkbuf_1 _07536_ (.A(_03354_),
    .X(_00540_));
 sky130_fd_sc_hd__clkbuf_2 _07537_ (.A(_03339_),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_1 _07538_ (.A0(\u_async_wb.u_cmd_if.mem[2][24] ),
    .A1(_02432_),
    .S(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_1 _07539_ (.A(_03356_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _07540_ (.A0(\u_async_wb.u_cmd_if.mem[2][25] ),
    .A1(_02438_),
    .S(_03355_),
    .X(_03357_));
 sky130_fd_sc_hd__clkbuf_1 _07541_ (.A(_03357_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _07542_ (.A0(\u_async_wb.u_cmd_if.mem[2][26] ),
    .A1(_02441_),
    .S(_03355_),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_1 _07543_ (.A(_03358_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _07544_ (.A0(\u_async_wb.u_cmd_if.mem[2][27] ),
    .A1(_02444_),
    .S(_03355_),
    .X(_03359_));
 sky130_fd_sc_hd__clkbuf_1 _07545_ (.A(_03359_),
    .X(_00544_));
 sky130_fd_sc_hd__clkbuf_2 _07546_ (.A(_03338_),
    .X(_03360_));
 sky130_fd_sc_hd__clkbuf_2 _07547_ (.A(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__mux2_1 _07548_ (.A0(\u_async_wb.u_cmd_if.mem[2][28] ),
    .A1(_02374_),
    .S(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__clkbuf_1 _07549_ (.A(_03362_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _07550_ (.A0(\u_async_wb.u_cmd_if.mem[2][29] ),
    .A1(_02380_),
    .S(_03361_),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_1 _07551_ (.A(_03363_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _07552_ (.A0(\u_async_wb.u_cmd_if.mem[2][30] ),
    .A1(_02385_),
    .S(_03361_),
    .X(_03364_));
 sky130_fd_sc_hd__clkbuf_1 _07553_ (.A(_03364_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _07554_ (.A0(\u_async_wb.u_cmd_if.mem[2][31] ),
    .A1(_02733_),
    .S(_03361_),
    .X(_03365_));
 sky130_fd_sc_hd__clkbuf_1 _07555_ (.A(_03365_),
    .X(_00548_));
 sky130_fd_sc_hd__clkbuf_2 _07556_ (.A(_03360_),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_1 _07557_ (.A0(\u_async_wb.u_cmd_if.mem[2][32] ),
    .A1(_02394_),
    .S(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_1 _07558_ (.A(_03367_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _07559_ (.A0(\u_async_wb.u_cmd_if.mem[2][33] ),
    .A1(_03227_),
    .S(_03366_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_1 _07560_ (.A(_03368_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _07561_ (.A0(\u_async_wb.u_cmd_if.mem[2][34] ),
    .A1(_02403_),
    .S(_03366_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_1 _07562_ (.A(_03369_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _07563_ (.A0(\u_async_wb.u_cmd_if.mem[2][35] ),
    .A1(_02407_),
    .S(_03366_),
    .X(_03370_));
 sky130_fd_sc_hd__clkbuf_1 _07564_ (.A(_03370_),
    .X(_00552_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07565_ (.A(_03360_),
    .X(_03371_));
 sky130_fd_sc_hd__mux2_1 _07566_ (.A0(\u_async_wb.u_cmd_if.mem[2][36] ),
    .A1(_03232_),
    .S(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__clkbuf_1 _07567_ (.A(_03372_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _07568_ (.A0(\u_async_wb.u_cmd_if.mem[2][37] ),
    .A1(_03237_),
    .S(_03371_),
    .X(_03373_));
 sky130_fd_sc_hd__clkbuf_1 _07569_ (.A(_03373_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _07570_ (.A0(\u_async_wb.u_cmd_if.mem[2][38] ),
    .A1(_03241_),
    .S(_03371_),
    .X(_03374_));
 sky130_fd_sc_hd__clkbuf_1 _07571_ (.A(_03374_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _07572_ (.A0(\u_async_wb.u_cmd_if.mem[2][39] ),
    .A1(_03243_),
    .S(_03371_),
    .X(_03375_));
 sky130_fd_sc_hd__clkbuf_1 _07573_ (.A(_03375_),
    .X(_00556_));
 sky130_fd_sc_hd__clkbuf_2 _07574_ (.A(_03360_),
    .X(_03376_));
 sky130_fd_sc_hd__mux2_1 _07575_ (.A0(\u_async_wb.u_cmd_if.mem[2][40] ),
    .A1(_03247_),
    .S(_03376_),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_1 _07576_ (.A(_03377_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _07577_ (.A0(\u_async_wb.u_cmd_if.mem[2][41] ),
    .A1(_03249_),
    .S(_03376_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_1 _07578_ (.A(_03378_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _07579_ (.A0(\u_async_wb.u_cmd_if.mem[2][42] ),
    .A1(_03254_),
    .S(_03376_),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_1 _07580_ (.A(_03379_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _07581_ (.A0(\u_async_wb.u_cmd_if.mem[2][43] ),
    .A1(_03257_),
    .S(_03376_),
    .X(_03380_));
 sky130_fd_sc_hd__clkbuf_1 _07582_ (.A(_03380_),
    .X(_00560_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07583_ (.A(_03321_),
    .X(_03381_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07584_ (.A(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__mux2_1 _07585_ (.A0(\u_async_wb.u_cmd_if.mem[2][44] ),
    .A1(_03261_),
    .S(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_1 _07586_ (.A(_03383_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _07587_ (.A0(\u_async_wb.u_cmd_if.mem[2][45] ),
    .A1(_03267_),
    .S(_03382_),
    .X(_03384_));
 sky130_fd_sc_hd__clkbuf_1 _07588_ (.A(_03384_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _07589_ (.A0(\u_async_wb.u_cmd_if.mem[2][46] ),
    .A1(_03271_),
    .S(_03382_),
    .X(_03385_));
 sky130_fd_sc_hd__clkbuf_1 _07590_ (.A(_03385_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _07591_ (.A0(\u_async_wb.u_cmd_if.mem[2][47] ),
    .A1(_03275_),
    .S(_03382_),
    .X(_03386_));
 sky130_fd_sc_hd__clkbuf_1 _07592_ (.A(_03386_),
    .X(_00564_));
 sky130_fd_sc_hd__clkbuf_2 _07593_ (.A(_03381_),
    .X(_03387_));
 sky130_fd_sc_hd__mux2_1 _07594_ (.A0(\u_async_wb.u_cmd_if.mem[2][48] ),
    .A1(_03279_),
    .S(_03387_),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_1 _07595_ (.A(_03388_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _07596_ (.A0(\u_async_wb.u_cmd_if.mem[2][49] ),
    .A1(_03283_),
    .S(_03387_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_1 _07597_ (.A(_03389_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _07598_ (.A0(\u_async_wb.u_cmd_if.mem[2][50] ),
    .A1(_03287_),
    .S(_03387_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _07599_ (.A(_03390_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _07600_ (.A0(\u_async_wb.u_cmd_if.mem[2][51] ),
    .A1(_03290_),
    .S(_03387_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_1 _07601_ (.A(_03391_),
    .X(_00568_));
 sky130_fd_sc_hd__clkbuf_2 _07602_ (.A(_03381_),
    .X(_03392_));
 sky130_fd_sc_hd__mux2_1 _07603_ (.A0(\u_async_wb.u_cmd_if.mem[2][52] ),
    .A1(_03294_),
    .S(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_1 _07604_ (.A(_03393_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _07605_ (.A0(\u_async_wb.u_cmd_if.mem[2][53] ),
    .A1(_03297_),
    .S(_03392_),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_1 _07606_ (.A(_03394_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _07607_ (.A0(\u_async_wb.u_cmd_if.mem[2][54] ),
    .A1(_03300_),
    .S(_03392_),
    .X(_03395_));
 sky130_fd_sc_hd__clkbuf_1 _07608_ (.A(_03395_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _07609_ (.A0(\u_async_wb.u_cmd_if.mem[2][55] ),
    .A1(_03303_),
    .S(_03392_),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_1 _07610_ (.A(_03396_),
    .X(_00572_));
 sky130_fd_sc_hd__clkbuf_2 _07611_ (.A(_03381_),
    .X(_03397_));
 sky130_fd_sc_hd__mux2_1 _07612_ (.A0(\u_async_wb.u_cmd_if.mem[2][56] ),
    .A1(_02249_),
    .S(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__clkbuf_1 _07613_ (.A(_03398_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _07614_ (.A0(\u_async_wb.u_cmd_if.mem[2][57] ),
    .A1(_02241_),
    .S(_03397_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_1 _07615_ (.A(_03399_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _07616_ (.A0(\u_async_wb.u_cmd_if.mem[2][58] ),
    .A1(_02235_),
    .S(_03397_),
    .X(_03400_));
 sky130_fd_sc_hd__clkbuf_1 _07617_ (.A(_03400_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _07618_ (.A0(\u_async_wb.u_cmd_if.mem[2][59] ),
    .A1(_02230_),
    .S(_03397_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_1 _07619_ (.A(_03401_),
    .X(_00576_));
 sky130_fd_sc_hd__clkbuf_2 _07620_ (.A(_03338_),
    .X(_03402_));
 sky130_fd_sc_hd__mux2_1 _07621_ (.A0(\u_async_wb.u_cmd_if.mem[2][60] ),
    .A1(_02224_),
    .S(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__clkbuf_1 _07622_ (.A(_03403_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _07623_ (.A0(\u_async_wb.u_cmd_if.mem[2][61] ),
    .A1(_02218_),
    .S(_03402_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_1 _07624_ (.A(_03404_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _07625_ (.A0(\u_async_wb.u_cmd_if.mem[2][62] ),
    .A1(_02410_),
    .S(_03402_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_1 _07626_ (.A(_03405_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _07627_ (.A0(\u_async_wb.u_cmd_if.mem[2][63] ),
    .A1(_02280_),
    .S(_03402_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_1 _07628_ (.A(_03406_),
    .X(_00580_));
 sky130_fd_sc_hd__clkbuf_2 _07629_ (.A(_03338_),
    .X(_03407_));
 sky130_fd_sc_hd__mux2_1 _07630_ (.A0(\u_async_wb.u_cmd_if.mem[2][64] ),
    .A1(_02277_),
    .S(_03407_),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _07631_ (.A(_03408_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _07632_ (.A0(\u_async_wb.u_cmd_if.mem[2][65] ),
    .A1(_02275_),
    .S(_03407_),
    .X(_03409_));
 sky130_fd_sc_hd__clkbuf_1 _07633_ (.A(_03409_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _07634_ (.A0(\u_async_wb.u_cmd_if.mem[2][66] ),
    .A1(_02273_),
    .S(_03407_),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_1 _07635_ (.A(_03410_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _07636_ (.A0(\u_async_wb.u_cmd_if.mem[2][67] ),
    .A1(_02271_),
    .S(_03407_),
    .X(_03411_));
 sky130_fd_sc_hd__clkbuf_1 _07637_ (.A(_03411_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _07638_ (.A0(\u_async_wb.u_cmd_if.mem[2][68] ),
    .A1(_02268_),
    .S(_03322_),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_1 _07639_ (.A(_03412_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _07640_ (.A0(_03179_),
    .A1(\u_async_wb.u_cmd_if.mem[1][0] ),
    .S(_02801_),
    .X(_03413_));
 sky130_fd_sc_hd__clkbuf_1 _07641_ (.A(_03413_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _07642_ (.A0(_03181_),
    .A1(\u_async_wb.u_cmd_if.mem[1][1] ),
    .S(_02801_),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _07643_ (.A(_03414_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _07644_ (.A0(_03183_),
    .A1(\u_async_wb.u_cmd_if.mem[1][2] ),
    .S(_02801_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_1 _07645_ (.A(_03415_),
    .X(_00588_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07646_ (.A(_02799_),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_2 _07647_ (.A(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_1 _07648_ (.A0(_03185_),
    .A1(\u_async_wb.u_cmd_if.mem[1][3] ),
    .S(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _07649_ (.A(_03418_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _07650_ (.A0(_02286_),
    .A1(\u_async_wb.u_cmd_if.mem[1][4] ),
    .S(_03417_),
    .X(_03419_));
 sky130_fd_sc_hd__clkbuf_1 _07651_ (.A(_03419_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _07652_ (.A0(_02266_),
    .A1(\u_async_wb.u_cmd_if.mem[1][5] ),
    .S(_03417_),
    .X(_03420_));
 sky130_fd_sc_hd__clkbuf_1 _07653_ (.A(_03420_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _07654_ (.A0(_02259_),
    .A1(\u_async_wb.u_cmd_if.mem[1][6] ),
    .S(_03417_),
    .X(_03421_));
 sky130_fd_sc_hd__clkbuf_1 _07655_ (.A(_03421_),
    .X(_00592_));
 sky130_fd_sc_hd__clkbuf_2 _07656_ (.A(_03416_),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_1 _07657_ (.A0(_02254_),
    .A1(\u_async_wb.u_cmd_if.mem[1][7] ),
    .S(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__clkbuf_1 _07658_ (.A(_03423_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _07659_ (.A0(_02246_),
    .A1(\u_async_wb.u_cmd_if.mem[1][8] ),
    .S(_03422_),
    .X(_03424_));
 sky130_fd_sc_hd__clkbuf_1 _07660_ (.A(_03424_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _07661_ (.A0(_02239_),
    .A1(\u_async_wb.u_cmd_if.mem[1][9] ),
    .S(_03422_),
    .X(_03425_));
 sky130_fd_sc_hd__clkbuf_1 _07662_ (.A(_03425_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _07663_ (.A0(_02473_),
    .A1(\u_async_wb.u_cmd_if.mem[1][10] ),
    .S(_03422_),
    .X(_03426_));
 sky130_fd_sc_hd__clkbuf_1 _07664_ (.A(_03426_),
    .X(_00596_));
 sky130_fd_sc_hd__clkbuf_2 _07665_ (.A(_02800_),
    .X(_03427_));
 sky130_fd_sc_hd__clkbuf_2 _07666_ (.A(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__mux2_1 _07667_ (.A0(_02228_),
    .A1(\u_async_wb.u_cmd_if.mem[1][11] ),
    .S(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__clkbuf_1 _07668_ (.A(_03429_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _07669_ (.A0(_02477_),
    .A1(\u_async_wb.u_cmd_if.mem[1][12] ),
    .S(_03428_),
    .X(_03430_));
 sky130_fd_sc_hd__clkbuf_1 _07670_ (.A(_03430_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _07671_ (.A0(_02181_),
    .A1(\u_async_wb.u_cmd_if.mem[1][13] ),
    .S(_03428_),
    .X(_03431_));
 sky130_fd_sc_hd__clkbuf_1 _07672_ (.A(_03431_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _07673_ (.A0(_02187_),
    .A1(\u_async_wb.u_cmd_if.mem[1][14] ),
    .S(_03428_),
    .X(_03432_));
 sky130_fd_sc_hd__clkbuf_1 _07674_ (.A(_03432_),
    .X(_00600_));
 sky130_fd_sc_hd__clkbuf_2 _07675_ (.A(_03427_),
    .X(_03433_));
 sky130_fd_sc_hd__mux2_1 _07676_ (.A0(_02485_),
    .A1(\u_async_wb.u_cmd_if.mem[1][15] ),
    .S(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__clkbuf_1 _07677_ (.A(_03434_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _07678_ (.A0(_02200_),
    .A1(\u_async_wb.u_cmd_if.mem[1][16] ),
    .S(_03433_),
    .X(_03435_));
 sky130_fd_sc_hd__clkbuf_1 _07679_ (.A(_03435_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _07680_ (.A0(_02206_),
    .A1(\u_async_wb.u_cmd_if.mem[1][17] ),
    .S(_03433_),
    .X(_03436_));
 sky130_fd_sc_hd__clkbuf_1 _07681_ (.A(_03436_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _07682_ (.A0(_02211_),
    .A1(\u_async_wb.u_cmd_if.mem[1][18] ),
    .S(_03433_),
    .X(_03437_));
 sky130_fd_sc_hd__clkbuf_1 _07683_ (.A(_03437_),
    .X(_00604_));
 sky130_fd_sc_hd__clkbuf_2 _07684_ (.A(_03427_),
    .X(_03438_));
 sky130_fd_sc_hd__mux2_1 _07685_ (.A0(_02493_),
    .A1(\u_async_wb.u_cmd_if.mem[1][19] ),
    .S(_03438_),
    .X(_03439_));
 sky130_fd_sc_hd__clkbuf_1 _07686_ (.A(_03439_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _07687_ (.A0(_02412_),
    .A1(\u_async_wb.u_cmd_if.mem[1][20] ),
    .S(_03438_),
    .X(_03440_));
 sky130_fd_sc_hd__clkbuf_1 _07688_ (.A(_03440_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _07689_ (.A0(_02423_),
    .A1(\u_async_wb.u_cmd_if.mem[1][21] ),
    .S(_03438_),
    .X(_03441_));
 sky130_fd_sc_hd__clkbuf_1 _07690_ (.A(_03441_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _07691_ (.A0(_02426_),
    .A1(\u_async_wb.u_cmd_if.mem[1][22] ),
    .S(_03438_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_1 _07692_ (.A(_03442_),
    .X(_00608_));
 sky130_fd_sc_hd__clkbuf_2 _07693_ (.A(_03427_),
    .X(_03443_));
 sky130_fd_sc_hd__mux2_1 _07694_ (.A0(_02430_),
    .A1(\u_async_wb.u_cmd_if.mem[1][23] ),
    .S(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__clkbuf_1 _07695_ (.A(_03444_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _07696_ (.A0(_02432_),
    .A1(\u_async_wb.u_cmd_if.mem[1][24] ),
    .S(_03443_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_1 _07697_ (.A(_03445_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _07698_ (.A0(_02438_),
    .A1(\u_async_wb.u_cmd_if.mem[1][25] ),
    .S(_03443_),
    .X(_03446_));
 sky130_fd_sc_hd__clkbuf_1 _07699_ (.A(_03446_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _07700_ (.A0(_02441_),
    .A1(\u_async_wb.u_cmd_if.mem[1][26] ),
    .S(_03443_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_1 _07701_ (.A(_03447_),
    .X(_00612_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07702_ (.A(_02799_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_2 _07703_ (.A(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__mux2_1 _07704_ (.A0(_02445_),
    .A1(\u_async_wb.u_cmd_if.mem[1][27] ),
    .S(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_1 _07705_ (.A(_03450_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _07706_ (.A0(_02513_),
    .A1(\u_async_wb.u_cmd_if.mem[1][28] ),
    .S(_03449_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_1 _07707_ (.A(_03451_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _07708_ (.A0(_02515_),
    .A1(\u_async_wb.u_cmd_if.mem[1][29] ),
    .S(_03449_),
    .X(_03452_));
 sky130_fd_sc_hd__clkbuf_1 _07709_ (.A(_03452_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _07710_ (.A0(_02521_),
    .A1(\u_async_wb.u_cmd_if.mem[1][30] ),
    .S(_03449_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_1 _07711_ (.A(_03453_),
    .X(_00616_));
 sky130_fd_sc_hd__clkbuf_2 _07712_ (.A(_03448_),
    .X(_03454_));
 sky130_fd_sc_hd__mux2_1 _07713_ (.A0(_02733_),
    .A1(\u_async_wb.u_cmd_if.mem[1][31] ),
    .S(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_1 _07714_ (.A(_03455_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _07715_ (.A0(_02525_),
    .A1(\u_async_wb.u_cmd_if.mem[1][32] ),
    .S(_03454_),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_1 _07716_ (.A(_03456_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _07717_ (.A0(_03227_),
    .A1(\u_async_wb.u_cmd_if.mem[1][33] ),
    .S(_03454_),
    .X(_03457_));
 sky130_fd_sc_hd__clkbuf_1 _07718_ (.A(_03457_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _07719_ (.A0(_02529_),
    .A1(\u_async_wb.u_cmd_if.mem[1][34] ),
    .S(_03454_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_1 _07720_ (.A(_03458_),
    .X(_00620_));
 sky130_fd_sc_hd__clkbuf_2 _07721_ (.A(_03448_),
    .X(_03459_));
 sky130_fd_sc_hd__mux2_1 _07722_ (.A0(_02531_),
    .A1(\u_async_wb.u_cmd_if.mem[1][35] ),
    .S(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_1 _07723_ (.A(_03460_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _07724_ (.A0(_03232_),
    .A1(\u_async_wb.u_cmd_if.mem[1][36] ),
    .S(_03459_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_1 _07725_ (.A(_03461_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _07726_ (.A0(_03237_),
    .A1(\u_async_wb.u_cmd_if.mem[1][37] ),
    .S(_03459_),
    .X(_03462_));
 sky130_fd_sc_hd__clkbuf_1 _07727_ (.A(_03462_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _07728_ (.A0(_03241_),
    .A1(\u_async_wb.u_cmd_if.mem[1][38] ),
    .S(_03459_),
    .X(_03463_));
 sky130_fd_sc_hd__clkbuf_1 _07729_ (.A(_03463_),
    .X(_00624_));
 sky130_fd_sc_hd__clkbuf_2 _07730_ (.A(_03448_),
    .X(_03464_));
 sky130_fd_sc_hd__mux2_1 _07731_ (.A0(_03243_),
    .A1(\u_async_wb.u_cmd_if.mem[1][39] ),
    .S(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_1 _07732_ (.A(_03465_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _07733_ (.A0(_03247_),
    .A1(\u_async_wb.u_cmd_if.mem[1][40] ),
    .S(_03464_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_1 _07734_ (.A(_03466_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _07735_ (.A0(_03249_),
    .A1(\u_async_wb.u_cmd_if.mem[1][41] ),
    .S(_03464_),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_1 _07736_ (.A(_03467_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _07737_ (.A0(_03254_),
    .A1(\u_async_wb.u_cmd_if.mem[1][42] ),
    .S(_03464_),
    .X(_03468_));
 sky130_fd_sc_hd__clkbuf_1 _07738_ (.A(_03468_),
    .X(_00628_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07739_ (.A(_02799_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_2 _07740_ (.A(_03469_),
    .X(_03470_));
 sky130_fd_sc_hd__mux2_1 _07741_ (.A0(_03257_),
    .A1(\u_async_wb.u_cmd_if.mem[1][43] ),
    .S(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_1 _07742_ (.A(_03471_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _07743_ (.A0(_03261_),
    .A1(\u_async_wb.u_cmd_if.mem[1][44] ),
    .S(_03470_),
    .X(_03472_));
 sky130_fd_sc_hd__clkbuf_1 _07744_ (.A(_03472_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _07745_ (.A0(_03267_),
    .A1(\u_async_wb.u_cmd_if.mem[1][45] ),
    .S(_03470_),
    .X(_03473_));
 sky130_fd_sc_hd__clkbuf_1 _07746_ (.A(_03473_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _07747_ (.A0(_03271_),
    .A1(\u_async_wb.u_cmd_if.mem[1][46] ),
    .S(_03470_),
    .X(_03474_));
 sky130_fd_sc_hd__clkbuf_1 _07748_ (.A(_03474_),
    .X(_00632_));
 sky130_fd_sc_hd__clkbuf_2 _07749_ (.A(_03469_),
    .X(_03475_));
 sky130_fd_sc_hd__mux2_1 _07750_ (.A0(_03275_),
    .A1(\u_async_wb.u_cmd_if.mem[1][47] ),
    .S(_03475_),
    .X(_03476_));
 sky130_fd_sc_hd__clkbuf_1 _07751_ (.A(_03476_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _07752_ (.A0(_03279_),
    .A1(\u_async_wb.u_cmd_if.mem[1][48] ),
    .S(_03475_),
    .X(_03477_));
 sky130_fd_sc_hd__clkbuf_1 _07753_ (.A(_03477_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _07754_ (.A0(_03283_),
    .A1(\u_async_wb.u_cmd_if.mem[1][49] ),
    .S(_03475_),
    .X(_03478_));
 sky130_fd_sc_hd__clkbuf_1 _07755_ (.A(_03478_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _07756_ (.A0(_03287_),
    .A1(\u_async_wb.u_cmd_if.mem[1][50] ),
    .S(_03475_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_1 _07757_ (.A(_03479_),
    .X(_00636_));
 sky130_fd_sc_hd__clkbuf_2 _07758_ (.A(_03469_),
    .X(_03480_));
 sky130_fd_sc_hd__mux2_1 _07759_ (.A0(_03290_),
    .A1(\u_async_wb.u_cmd_if.mem[1][51] ),
    .S(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__clkbuf_1 _07760_ (.A(_03481_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _07761_ (.A0(_03294_),
    .A1(\u_async_wb.u_cmd_if.mem[1][52] ),
    .S(_03480_),
    .X(_03482_));
 sky130_fd_sc_hd__clkbuf_1 _07762_ (.A(_03482_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _07763_ (.A0(_03297_),
    .A1(\u_async_wb.u_cmd_if.mem[1][53] ),
    .S(_03480_),
    .X(_03483_));
 sky130_fd_sc_hd__clkbuf_1 _07764_ (.A(_03483_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _07765_ (.A0(_03300_),
    .A1(\u_async_wb.u_cmd_if.mem[1][54] ),
    .S(_03480_),
    .X(_03484_));
 sky130_fd_sc_hd__clkbuf_1 _07766_ (.A(_03484_),
    .X(_00640_));
 sky130_fd_sc_hd__clkbuf_2 _07767_ (.A(_03469_),
    .X(_03485_));
 sky130_fd_sc_hd__mux2_1 _07768_ (.A0(_03303_),
    .A1(\u_async_wb.u_cmd_if.mem[1][55] ),
    .S(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__clkbuf_1 _07769_ (.A(_03486_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _07770_ (.A0(_02249_),
    .A1(\u_async_wb.u_cmd_if.mem[1][56] ),
    .S(_03485_),
    .X(_03487_));
 sky130_fd_sc_hd__clkbuf_1 _07771_ (.A(_03487_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _07772_ (.A0(_02241_),
    .A1(\u_async_wb.u_cmd_if.mem[1][57] ),
    .S(_03485_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_1 _07773_ (.A(_03488_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _07774_ (.A0(_02235_),
    .A1(\u_async_wb.u_cmd_if.mem[1][58] ),
    .S(_03485_),
    .X(_03489_));
 sky130_fd_sc_hd__clkbuf_1 _07775_ (.A(_03489_),
    .X(_00644_));
 sky130_fd_sc_hd__clkbuf_2 _07776_ (.A(_02800_),
    .X(_03490_));
 sky130_fd_sc_hd__mux2_1 _07777_ (.A0(_02230_),
    .A1(\u_async_wb.u_cmd_if.mem[1][59] ),
    .S(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__clkbuf_1 _07778_ (.A(_03491_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _07779_ (.A0(_02224_),
    .A1(\u_async_wb.u_cmd_if.mem[1][60] ),
    .S(_03490_),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_1 _07780_ (.A(_03492_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _07781_ (.A0(_02218_),
    .A1(\u_async_wb.u_cmd_if.mem[1][61] ),
    .S(_03490_),
    .X(_03493_));
 sky130_fd_sc_hd__clkbuf_1 _07782_ (.A(_03493_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _07783_ (.A0(_02410_),
    .A1(\u_async_wb.u_cmd_if.mem[1][62] ),
    .S(_03490_),
    .X(_03494_));
 sky130_fd_sc_hd__clkbuf_1 _07784_ (.A(_03494_),
    .X(_00648_));
 sky130_fd_sc_hd__clkbuf_2 _07785_ (.A(_02800_),
    .X(_03495_));
 sky130_fd_sc_hd__mux2_1 _07786_ (.A0(_02280_),
    .A1(\u_async_wb.u_cmd_if.mem[1][63] ),
    .S(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__clkbuf_1 _07787_ (.A(_03496_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _07788_ (.A0(_02277_),
    .A1(\u_async_wb.u_cmd_if.mem[1][64] ),
    .S(_03495_),
    .X(_03497_));
 sky130_fd_sc_hd__clkbuf_1 _07789_ (.A(_03497_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _07790_ (.A0(_02275_),
    .A1(\u_async_wb.u_cmd_if.mem[1][65] ),
    .S(_03495_),
    .X(_03498_));
 sky130_fd_sc_hd__clkbuf_1 _07791_ (.A(_03498_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _07792_ (.A0(_02273_),
    .A1(\u_async_wb.u_cmd_if.mem[1][66] ),
    .S(_03495_),
    .X(_03499_));
 sky130_fd_sc_hd__clkbuf_1 _07793_ (.A(_03499_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _07794_ (.A0(_02271_),
    .A1(\u_async_wb.u_cmd_if.mem[1][67] ),
    .S(_03416_),
    .X(_03500_));
 sky130_fd_sc_hd__clkbuf_1 _07795_ (.A(_03500_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _07796_ (.A0(_02268_),
    .A1(\u_async_wb.u_cmd_if.mem[1][68] ),
    .S(_03416_),
    .X(_03501_));
 sky130_fd_sc_hd__clkbuf_1 _07797_ (.A(_03501_),
    .X(_00654_));
 sky130_fd_sc_hd__and2_1 _07798_ (.A(_01491_),
    .B(_01501_),
    .X(_03502_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07799_ (.A(_03502_),
    .X(_03503_));
 sky130_fd_sc_hd__clkbuf_2 _07800_ (.A(_03503_),
    .X(_03504_));
 sky130_fd_sc_hd__mux2_1 _07801_ (.A0(\u_async_wb.u_cmd_if.mem[0][0] ),
    .A1(_03179_),
    .S(_03504_),
    .X(_03505_));
 sky130_fd_sc_hd__clkbuf_1 _07802_ (.A(_03505_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _07803_ (.A0(\u_async_wb.u_cmd_if.mem[0][1] ),
    .A1(_03181_),
    .S(_03504_),
    .X(_03506_));
 sky130_fd_sc_hd__clkbuf_1 _07804_ (.A(_03506_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _07805_ (.A0(\u_async_wb.u_cmd_if.mem[0][2] ),
    .A1(_03183_),
    .S(_03504_),
    .X(_03507_));
 sky130_fd_sc_hd__clkbuf_1 _07806_ (.A(_03507_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _07807_ (.A0(\u_async_wb.u_cmd_if.mem[0][3] ),
    .A1(_03185_),
    .S(_03504_),
    .X(_03508_));
 sky130_fd_sc_hd__clkbuf_1 _07808_ (.A(_03508_),
    .X(_00658_));
 sky130_fd_sc_hd__clkbuf_2 _07809_ (.A(_03503_),
    .X(_03509_));
 sky130_fd_sc_hd__mux2_1 _07810_ (.A0(\u_async_wb.u_cmd_if.mem[0][4] ),
    .A1(_02285_),
    .S(_03509_),
    .X(_03510_));
 sky130_fd_sc_hd__clkbuf_1 _07811_ (.A(_03510_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _07812_ (.A0(\u_async_wb.u_cmd_if.mem[0][5] ),
    .A1(_02265_),
    .S(_03509_),
    .X(_03511_));
 sky130_fd_sc_hd__clkbuf_1 _07813_ (.A(_03511_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _07814_ (.A0(\u_async_wb.u_cmd_if.mem[0][6] ),
    .A1(_02258_),
    .S(_03509_),
    .X(_03512_));
 sky130_fd_sc_hd__clkbuf_1 _07815_ (.A(_03512_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _07816_ (.A0(\u_async_wb.u_cmd_if.mem[0][7] ),
    .A1(_02253_),
    .S(_03509_),
    .X(_03513_));
 sky130_fd_sc_hd__clkbuf_1 _07817_ (.A(_03513_),
    .X(_00662_));
 sky130_fd_sc_hd__clkbuf_2 _07818_ (.A(_03503_),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_1 _07819_ (.A0(\u_async_wb.u_cmd_if.mem[0][8] ),
    .A1(_02245_),
    .S(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__clkbuf_1 _07820_ (.A(_03515_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _07821_ (.A0(\u_async_wb.u_cmd_if.mem[0][9] ),
    .A1(_02238_),
    .S(_03514_),
    .X(_03516_));
 sky130_fd_sc_hd__clkbuf_1 _07822_ (.A(_03516_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _07823_ (.A0(\u_async_wb.u_cmd_if.mem[0][10] ),
    .A1(_02233_),
    .S(_03514_),
    .X(_03517_));
 sky130_fd_sc_hd__clkbuf_1 _07824_ (.A(_03517_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _07825_ (.A0(\u_async_wb.u_cmd_if.mem[0][11] ),
    .A1(_02227_),
    .S(_03514_),
    .X(_03518_));
 sky130_fd_sc_hd__clkbuf_1 _07826_ (.A(_03518_),
    .X(_00666_));
 sky130_fd_sc_hd__clkbuf_2 _07827_ (.A(_03502_),
    .X(_03519_));
 sky130_fd_sc_hd__clkbuf_2 _07828_ (.A(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__clkbuf_2 _07829_ (.A(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__mux2_1 _07830_ (.A0(\u_async_wb.u_cmd_if.mem[0][12] ),
    .A1(_02154_),
    .S(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__clkbuf_1 _07831_ (.A(_03522_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _07832_ (.A0(\u_async_wb.u_cmd_if.mem[0][13] ),
    .A1(_02180_),
    .S(_03521_),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_1 _07833_ (.A(_03523_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _07834_ (.A0(\u_async_wb.u_cmd_if.mem[0][14] ),
    .A1(_02186_),
    .S(_03521_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_1 _07835_ (.A(_03524_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _07836_ (.A0(\u_async_wb.u_cmd_if.mem[0][15] ),
    .A1(_02191_),
    .S(_03521_),
    .X(_03525_));
 sky130_fd_sc_hd__clkbuf_1 _07837_ (.A(_03525_),
    .X(_00670_));
 sky130_fd_sc_hd__clkbuf_2 _07838_ (.A(_03520_),
    .X(_03526_));
 sky130_fd_sc_hd__mux2_1 _07839_ (.A0(\u_async_wb.u_cmd_if.mem[0][16] ),
    .A1(_02199_),
    .S(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__clkbuf_1 _07840_ (.A(_03527_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _07841_ (.A0(\u_async_wb.u_cmd_if.mem[0][17] ),
    .A1(_02205_),
    .S(_03526_),
    .X(_03528_));
 sky130_fd_sc_hd__clkbuf_1 _07842_ (.A(_03528_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _07843_ (.A0(\u_async_wb.u_cmd_if.mem[0][18] ),
    .A1(_02210_),
    .S(_03526_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_1 _07844_ (.A(_03529_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _07845_ (.A0(\u_async_wb.u_cmd_if.mem[0][19] ),
    .A1(_02216_),
    .S(_03526_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_1 _07846_ (.A(_03530_),
    .X(_00674_));
 sky130_fd_sc_hd__clkbuf_2 _07847_ (.A(_03520_),
    .X(_03531_));
 sky130_fd_sc_hd__mux2_1 _07848_ (.A0(\u_async_wb.u_cmd_if.mem[0][20] ),
    .A1(_02412_),
    .S(_03531_),
    .X(_03532_));
 sky130_fd_sc_hd__clkbuf_1 _07849_ (.A(_03532_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _07850_ (.A0(\u_async_wb.u_cmd_if.mem[0][21] ),
    .A1(_02423_),
    .S(_03531_),
    .X(_03533_));
 sky130_fd_sc_hd__clkbuf_1 _07851_ (.A(_03533_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _07852_ (.A0(\u_async_wb.u_cmd_if.mem[0][22] ),
    .A1(_02426_),
    .S(_03531_),
    .X(_03534_));
 sky130_fd_sc_hd__clkbuf_1 _07853_ (.A(_03534_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _07854_ (.A0(\u_async_wb.u_cmd_if.mem[0][23] ),
    .A1(_02429_),
    .S(_03531_),
    .X(_03535_));
 sky130_fd_sc_hd__clkbuf_1 _07855_ (.A(_03535_),
    .X(_00678_));
 sky130_fd_sc_hd__clkbuf_2 _07856_ (.A(_03520_),
    .X(_03536_));
 sky130_fd_sc_hd__mux2_1 _07857_ (.A0(\u_async_wb.u_cmd_if.mem[0][24] ),
    .A1(_02432_),
    .S(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__clkbuf_1 _07858_ (.A(_03537_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _07859_ (.A0(\u_async_wb.u_cmd_if.mem[0][25] ),
    .A1(_02438_),
    .S(_03536_),
    .X(_03538_));
 sky130_fd_sc_hd__clkbuf_1 _07860_ (.A(_03538_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _07861_ (.A0(\u_async_wb.u_cmd_if.mem[0][26] ),
    .A1(_02441_),
    .S(_03536_),
    .X(_03539_));
 sky130_fd_sc_hd__clkbuf_1 _07862_ (.A(_03539_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _07863_ (.A0(\u_async_wb.u_cmd_if.mem[0][27] ),
    .A1(_02444_),
    .S(_03536_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_1 _07864_ (.A(_03540_),
    .X(_00682_));
 sky130_fd_sc_hd__clkbuf_2 _07865_ (.A(_03519_),
    .X(_03541_));
 sky130_fd_sc_hd__clkbuf_2 _07866_ (.A(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__mux2_1 _07867_ (.A0(\u_async_wb.u_cmd_if.mem[0][28] ),
    .A1(_02374_),
    .S(_03542_),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_1 _07868_ (.A(_03543_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _07869_ (.A0(\u_async_wb.u_cmd_if.mem[0][29] ),
    .A1(_02380_),
    .S(_03542_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _07870_ (.A(_03544_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _07871_ (.A0(\u_async_wb.u_cmd_if.mem[0][30] ),
    .A1(_02385_),
    .S(_03542_),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _07872_ (.A(_03545_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _07873_ (.A0(\u_async_wb.u_cmd_if.mem[0][31] ),
    .A1(_02390_),
    .S(_03542_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _07874_ (.A(_03546_),
    .X(_00686_));
 sky130_fd_sc_hd__clkbuf_2 _07875_ (.A(_03541_),
    .X(_03547_));
 sky130_fd_sc_hd__mux2_1 _07876_ (.A0(\u_async_wb.u_cmd_if.mem[0][32] ),
    .A1(_02394_),
    .S(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__clkbuf_1 _07877_ (.A(_03548_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _07878_ (.A0(\u_async_wb.u_cmd_if.mem[0][33] ),
    .A1(_02399_),
    .S(_03547_),
    .X(_03549_));
 sky130_fd_sc_hd__clkbuf_1 _07879_ (.A(_03549_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _07880_ (.A0(\u_async_wb.u_cmd_if.mem[0][34] ),
    .A1(_02403_),
    .S(_03547_),
    .X(_03550_));
 sky130_fd_sc_hd__clkbuf_1 _07881_ (.A(_03550_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _07882_ (.A0(\u_async_wb.u_cmd_if.mem[0][35] ),
    .A1(_02407_),
    .S(_03547_),
    .X(_03551_));
 sky130_fd_sc_hd__clkbuf_1 _07883_ (.A(_03551_),
    .X(_00690_));
 sky130_fd_sc_hd__clkbuf_2 _07884_ (.A(_03541_),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_1 _07885_ (.A0(\u_async_wb.u_cmd_if.mem[0][36] ),
    .A1(_03232_),
    .S(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _07886_ (.A(_03553_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _07887_ (.A0(\u_async_wb.u_cmd_if.mem[0][37] ),
    .A1(_03237_),
    .S(_03552_),
    .X(_03554_));
 sky130_fd_sc_hd__clkbuf_1 _07888_ (.A(_03554_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _07889_ (.A0(\u_async_wb.u_cmd_if.mem[0][38] ),
    .A1(_03241_),
    .S(_03552_),
    .X(_03555_));
 sky130_fd_sc_hd__clkbuf_1 _07890_ (.A(_03555_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _07891_ (.A0(\u_async_wb.u_cmd_if.mem[0][39] ),
    .A1(_03243_),
    .S(_03552_),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_1 _07892_ (.A(_03556_),
    .X(_00694_));
 sky130_fd_sc_hd__clkbuf_2 _07893_ (.A(_03541_),
    .X(_03557_));
 sky130_fd_sc_hd__mux2_1 _07894_ (.A0(\u_async_wb.u_cmd_if.mem[0][40] ),
    .A1(_03247_),
    .S(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__clkbuf_1 _07895_ (.A(_03558_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _07896_ (.A0(\u_async_wb.u_cmd_if.mem[0][41] ),
    .A1(_03249_),
    .S(_03557_),
    .X(_03559_));
 sky130_fd_sc_hd__clkbuf_1 _07897_ (.A(_03559_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _07898_ (.A0(\u_async_wb.u_cmd_if.mem[0][42] ),
    .A1(_03254_),
    .S(_03557_),
    .X(_03560_));
 sky130_fd_sc_hd__clkbuf_1 _07899_ (.A(_03560_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _07900_ (.A0(\u_async_wb.u_cmd_if.mem[0][43] ),
    .A1(_03257_),
    .S(_03557_),
    .X(_03561_));
 sky130_fd_sc_hd__clkbuf_1 _07901_ (.A(_03561_),
    .X(_00698_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07902_ (.A(_03502_),
    .X(_03562_));
 sky130_fd_sc_hd__clkbuf_2 _07903_ (.A(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_1 _07904_ (.A0(\u_async_wb.u_cmd_if.mem[0][44] ),
    .A1(_03261_),
    .S(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_1 _07905_ (.A(_03564_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _07906_ (.A0(\u_async_wb.u_cmd_if.mem[0][45] ),
    .A1(_03267_),
    .S(_03563_),
    .X(_03565_));
 sky130_fd_sc_hd__clkbuf_1 _07907_ (.A(_03565_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _07908_ (.A0(\u_async_wb.u_cmd_if.mem[0][46] ),
    .A1(_03271_),
    .S(_03563_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_1 _07909_ (.A(_03566_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _07910_ (.A0(\u_async_wb.u_cmd_if.mem[0][47] ),
    .A1(_03275_),
    .S(_03563_),
    .X(_03567_));
 sky130_fd_sc_hd__clkbuf_1 _07911_ (.A(_03567_),
    .X(_00702_));
 sky130_fd_sc_hd__clkbuf_2 _07912_ (.A(_03562_),
    .X(_03568_));
 sky130_fd_sc_hd__mux2_1 _07913_ (.A0(\u_async_wb.u_cmd_if.mem[0][48] ),
    .A1(_03279_),
    .S(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__clkbuf_1 _07914_ (.A(_03569_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _07915_ (.A0(\u_async_wb.u_cmd_if.mem[0][49] ),
    .A1(_03283_),
    .S(_03568_),
    .X(_03570_));
 sky130_fd_sc_hd__clkbuf_1 _07916_ (.A(_03570_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _07917_ (.A0(\u_async_wb.u_cmd_if.mem[0][50] ),
    .A1(_03287_),
    .S(_03568_),
    .X(_03571_));
 sky130_fd_sc_hd__clkbuf_1 _07918_ (.A(_03571_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _07919_ (.A0(\u_async_wb.u_cmd_if.mem[0][51] ),
    .A1(_03290_),
    .S(_03568_),
    .X(_03572_));
 sky130_fd_sc_hd__clkbuf_1 _07920_ (.A(_03572_),
    .X(_00706_));
 sky130_fd_sc_hd__clkbuf_2 _07921_ (.A(_03562_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_1 _07922_ (.A0(\u_async_wb.u_cmd_if.mem[0][52] ),
    .A1(_03294_),
    .S(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__clkbuf_1 _07923_ (.A(_03574_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _07924_ (.A0(\u_async_wb.u_cmd_if.mem[0][53] ),
    .A1(_03297_),
    .S(_03573_),
    .X(_03575_));
 sky130_fd_sc_hd__clkbuf_1 _07925_ (.A(_03575_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _07926_ (.A0(\u_async_wb.u_cmd_if.mem[0][54] ),
    .A1(_03300_),
    .S(_03573_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_1 _07927_ (.A(_03576_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _07928_ (.A0(\u_async_wb.u_cmd_if.mem[0][55] ),
    .A1(_03303_),
    .S(_03573_),
    .X(_03577_));
 sky130_fd_sc_hd__clkbuf_1 _07929_ (.A(_03577_),
    .X(_00710_));
 sky130_fd_sc_hd__clkbuf_2 _07930_ (.A(_03562_),
    .X(_03578_));
 sky130_fd_sc_hd__mux2_1 _07931_ (.A0(\u_async_wb.u_cmd_if.mem[0][56] ),
    .A1(\u_async_wb.m_cmd_wr_data[56] ),
    .S(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__clkbuf_1 _07932_ (.A(_03579_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _07933_ (.A0(\u_async_wb.u_cmd_if.mem[0][57] ),
    .A1(\u_async_wb.m_cmd_wr_data[57] ),
    .S(_03578_),
    .X(_03580_));
 sky130_fd_sc_hd__clkbuf_1 _07934_ (.A(_03580_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _07935_ (.A0(\u_async_wb.u_cmd_if.mem[0][58] ),
    .A1(\u_async_wb.m_cmd_wr_data[58] ),
    .S(_03578_),
    .X(_03581_));
 sky130_fd_sc_hd__clkbuf_1 _07936_ (.A(_03581_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _07937_ (.A0(\u_async_wb.u_cmd_if.mem[0][59] ),
    .A1(\u_async_wb.m_cmd_wr_data[59] ),
    .S(_03578_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_1 _07938_ (.A(_03582_),
    .X(_00714_));
 sky130_fd_sc_hd__clkbuf_2 _07939_ (.A(_03519_),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_1 _07940_ (.A0(\u_async_wb.u_cmd_if.mem[0][60] ),
    .A1(\u_async_wb.m_cmd_wr_data[60] ),
    .S(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _07941_ (.A(_03584_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _07942_ (.A0(\u_async_wb.u_cmd_if.mem[0][61] ),
    .A1(\u_async_wb.m_cmd_wr_data[61] ),
    .S(_03583_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_1 _07943_ (.A(_03585_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _07944_ (.A0(\u_async_wb.u_cmd_if.mem[0][62] ),
    .A1(\u_async_wb.m_cmd_wr_data[62] ),
    .S(_03583_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_1 _07945_ (.A(_03586_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _07946_ (.A0(\u_async_wb.u_cmd_if.mem[0][63] ),
    .A1(\u_async_wb.m_cmd_wr_data[63] ),
    .S(_03583_),
    .X(_03587_));
 sky130_fd_sc_hd__clkbuf_1 _07947_ (.A(_03587_),
    .X(_00718_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07948_ (.A(_03519_),
    .X(_03588_));
 sky130_fd_sc_hd__mux2_1 _07949_ (.A0(\u_async_wb.u_cmd_if.mem[0][64] ),
    .A1(\u_async_wb.m_cmd_wr_data[64] ),
    .S(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__clkbuf_1 _07950_ (.A(_03589_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _07951_ (.A0(\u_async_wb.u_cmd_if.mem[0][65] ),
    .A1(\u_async_wb.m_cmd_wr_data[65] ),
    .S(_03588_),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _07952_ (.A(_03590_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _07953_ (.A0(\u_async_wb.u_cmd_if.mem[0][66] ),
    .A1(\u_async_wb.m_cmd_wr_data[66] ),
    .S(_03588_),
    .X(_03591_));
 sky130_fd_sc_hd__clkbuf_1 _07954_ (.A(_03591_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _07955_ (.A0(\u_async_wb.u_cmd_if.mem[0][67] ),
    .A1(\u_async_wb.m_cmd_wr_data[67] ),
    .S(_03588_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _07956_ (.A(_03592_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _07957_ (.A0(\u_async_wb.u_cmd_if.mem[0][68] ),
    .A1(\u_async_wb.m_cmd_wr_data[68] ),
    .S(_03503_),
    .X(_03593_));
 sky130_fd_sc_hd__clkbuf_1 _07958_ (.A(_03593_),
    .X(_00723_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07959_ (.A(_02694_),
    .X(_03594_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07960_ (.A(_02725_),
    .X(_03595_));
 sky130_fd_sc_hd__a22o_1 _07961_ (.A1(net1),
    .A2(_03594_),
    .B1(_03595_),
    .B2(_02286_),
    .X(_00724_));
 sky130_fd_sc_hd__clkbuf_2 _07962_ (.A(_02712_),
    .X(_03596_));
 sky130_fd_sc_hd__clkbuf_2 _07963_ (.A(_02714_),
    .X(_03597_));
 sky130_fd_sc_hd__o22a_1 _07964_ (.A1(net27),
    .A2(_03596_),
    .B1(_03597_),
    .B2(_02246_),
    .X(_00725_));
 sky130_fd_sc_hd__a22o_1 _07965_ (.A1(net31),
    .A2(_03594_),
    .B1(_03595_),
    .B2(_02477_),
    .X(_00726_));
 sky130_fd_sc_hd__o22a_1 _07966_ (.A1(net4),
    .A2(_03596_),
    .B1(_03597_),
    .B2(_02200_),
    .X(_00727_));
 sky130_fd_sc_hd__a22o_1 _07967_ (.A1(net8),
    .A2(_03594_),
    .B1(_03595_),
    .B2(_02413_),
    .X(_00728_));
 sky130_fd_sc_hd__o22a_1 _07968_ (.A1(net13),
    .A2(_03596_),
    .B1(_03597_),
    .B2(_02433_),
    .X(_00729_));
 sky130_fd_sc_hd__a22o_1 _07969_ (.A1(net17),
    .A2(_03594_),
    .B1(_03595_),
    .B2(_02513_),
    .X(_00730_));
 sky130_fd_sc_hd__or2_1 _07970_ (.A(\u_spi2wb.u_if.adr_phase ),
    .B(\u_spi2wb.u_if.wr_phase ),
    .X(_03598_));
 sky130_fd_sc_hd__or3_1 _07971_ (.A(\u_spi2wb.u_if.cmd_phase ),
    .B(\u_spi2wb.u_if.spi_if_st[1] ),
    .C(\u_spi2wb.u_if.spi_if_st[5] ),
    .X(_03599_));
 sky130_fd_sc_hd__or3_1 _07972_ (.A(\u_spi2wb.u_if.rd_phase ),
    .B(_03598_),
    .C(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__and3_1 _07973_ (.A(_01110_),
    .B(_01130_),
    .C(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__mux2_1 _07974_ (.A0(_01111_),
    .A1(_01130_),
    .S(_03600_),
    .X(_03602_));
 sky130_fd_sc_hd__nor2_1 _07975_ (.A(_01459_),
    .B(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__clkbuf_1 _07976_ (.A(\u_spi2wb.u_if.bitcnt[0] ),
    .X(_03604_));
 sky130_fd_sc_hd__mux2_1 _07977_ (.A0(_03601_),
    .A1(_03603_),
    .S(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__clkbuf_1 _07978_ (.A(_03605_),
    .X(_00731_));
 sky130_fd_sc_hd__clkbuf_1 _07979_ (.A(\u_spi2wb.u_if.bitcnt[1] ),
    .X(_03606_));
 sky130_fd_sc_hd__nand2_1 _07980_ (.A(_03606_),
    .B(_03604_),
    .Y(_03607_));
 sky130_fd_sc_hd__clkbuf_1 _07981_ (.A(_03601_),
    .X(_03608_));
 sky130_fd_sc_hd__or2_1 _07982_ (.A(_03606_),
    .B(_03604_),
    .X(_03609_));
 sky130_fd_sc_hd__clkbuf_1 _07983_ (.A(_03603_),
    .X(_03610_));
 sky130_fd_sc_hd__a32o_1 _07984_ (.A1(_03607_),
    .A2(_03608_),
    .A3(_03609_),
    .B1(_03610_),
    .B2(_03606_),
    .X(_00732_));
 sky130_fd_sc_hd__a21o_1 _07985_ (.A1(_03606_),
    .A2(_03604_),
    .B1(\u_spi2wb.u_if.bitcnt[2] ),
    .X(_03611_));
 sky130_fd_sc_hd__a32o_1 _07986_ (.A1(_01115_),
    .A2(_03608_),
    .A3(_03611_),
    .B1(_03610_),
    .B2(\u_spi2wb.u_if.bitcnt[2] ),
    .X(_00733_));
 sky130_fd_sc_hd__o32a_1 _07987_ (.A1(_01120_),
    .A2(_01116_),
    .A3(_03598_),
    .B1(_01114_),
    .B2(\u_spi2wb.u_if.bitcnt[3] ),
    .X(_03612_));
 sky130_fd_sc_hd__nand2_1 _07988_ (.A(_03601_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__a2bb2o_1 _07989_ (.A1_N(_01125_),
    .A2_N(_03613_),
    .B1(_03610_),
    .B2(\u_spi2wb.u_if.bitcnt[3] ),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _07990_ (.A(\u_spi2wb.u_if.bitcnt[4] ),
    .B(_01125_),
    .X(_03614_));
 sky130_fd_sc_hd__a32o_1 _07991_ (.A1(_01127_),
    .A2(_03608_),
    .A3(_03614_),
    .B1(_03603_),
    .B2(\u_spi2wb.u_if.bitcnt[4] ),
    .X(_00735_));
 sky130_fd_sc_hd__or3b_1 _07992_ (.A(_01128_),
    .B(_01127_),
    .C_N(_03599_),
    .X(_03615_));
 sky130_fd_sc_hd__a21bo_1 _07993_ (.A1(_01128_),
    .A2(_01127_),
    .B1_N(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__a22o_1 _07994_ (.A1(_01128_),
    .A2(_03610_),
    .B1(_03616_),
    .B2(_03608_),
    .X(_00736_));
 sky130_fd_sc_hd__and2b_1 _07995_ (.A_N(\u_uart2wb.u_async_reg_bus.in_state[1] ),
    .B(\u_uart2wb.u_async_reg_bus.in_state[0] ),
    .X(_03617_));
 sky130_fd_sc_hd__and3_1 _07996_ (.A(\u_uart2wb.u_async_reg_bus.out_flag_ss ),
    .B(_01739_),
    .C(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__clkbuf_1 _07997_ (.A(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__clkbuf_1 _07998_ (.A(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _07999_ (.A(\u_uart2wb.u_async_reg_bus.in_state[1] ),
    .X(_03621_));
 sky130_fd_sc_hd__and4_1 _08000_ (.A(\u_uart2wb.u_async_reg_bus.in_timer[1] ),
    .B(\u_uart2wb.u_async_reg_bus.in_timer[0] ),
    .C(\u_uart2wb.u_async_reg_bus.in_timer[3] ),
    .D(\u_uart2wb.u_async_reg_bus.in_timer[2] ),
    .X(_03622_));
 sky130_fd_sc_hd__and3_1 _08001_ (.A(\u_uart2wb.u_async_reg_bus.in_timer[5] ),
    .B(\u_uart2wb.u_async_reg_bus.in_timer[4] ),
    .C(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__and2_1 _08002_ (.A(\u_uart2wb.u_async_reg_bus.in_timer[6] ),
    .B(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__a31o_1 _08003_ (.A1(\u_uart2wb.u_async_reg_bus.in_timer[7] ),
    .A2(\u_uart2wb.u_async_reg_bus.in_timer[8] ),
    .A3(_03624_),
    .B1(\u_uart2wb.u_async_reg_bus.out_flag_ss ),
    .X(_03625_));
 sky130_fd_sc_hd__clkbuf_1 _08004_ (.A(\u_uart2wb.u_async_reg_bus.in_state[0] ),
    .X(_03626_));
 sky130_fd_sc_hd__o21ai_1 _08005_ (.A1(_03621_),
    .A2(_03625_),
    .B1(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08006_ (.A(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__a22o_1 _08007_ (.A1(\wb_dat_o[0] ),
    .A2(_03620_),
    .B1(_03628_),
    .B2(\u_uart2wb.reg_rdata[0] ),
    .X(_00737_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08008_ (.A(\u_uart2wb.reg_rdata[1] ),
    .X(_03629_));
 sky130_fd_sc_hd__a22o_1 _08009_ (.A1(\wb_dat_o[1] ),
    .A2(_03620_),
    .B1(_03628_),
    .B2(_03629_),
    .X(_00738_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08010_ (.A(\u_uart2wb.reg_rdata[2] ),
    .X(_03630_));
 sky130_fd_sc_hd__a22o_1 _08011_ (.A1(\wb_dat_o[2] ),
    .A2(_03620_),
    .B1(_03628_),
    .B2(_03630_),
    .X(_00739_));
 sky130_fd_sc_hd__clkbuf_2 _08012_ (.A(_03627_),
    .X(_03631_));
 sky130_fd_sc_hd__clkbuf_1 _08013_ (.A(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__a22o_1 _08014_ (.A1(\wb_dat_o[3] ),
    .A2(_03620_),
    .B1(_03632_),
    .B2(\u_uart2wb.reg_rdata[3] ),
    .X(_00740_));
 sky130_fd_sc_hd__clkbuf_1 _08015_ (.A(_03619_),
    .X(_03633_));
 sky130_fd_sc_hd__a22o_1 _08016_ (.A1(\wb_dat_o[4] ),
    .A2(_03633_),
    .B1(_03632_),
    .B2(\u_uart2wb.reg_rdata[4] ),
    .X(_00741_));
 sky130_fd_sc_hd__a22o_1 _08017_ (.A1(\wb_dat_o[5] ),
    .A2(_03633_),
    .B1(_03632_),
    .B2(_03032_),
    .X(_00742_));
 sky130_fd_sc_hd__a22o_1 _08018_ (.A1(\wb_dat_o[6] ),
    .A2(_03633_),
    .B1(_03632_),
    .B2(_03031_),
    .X(_00743_));
 sky130_fd_sc_hd__clkbuf_1 _08019_ (.A(_03631_),
    .X(_03634_));
 sky130_fd_sc_hd__a22o_1 _08020_ (.A1(\wb_dat_o[7] ),
    .A2(_03633_),
    .B1(_03634_),
    .B2(\u_uart2wb.reg_rdata[7] ),
    .X(_00744_));
 sky130_fd_sc_hd__clkbuf_1 _08021_ (.A(_03619_),
    .X(_03635_));
 sky130_fd_sc_hd__a22o_1 _08022_ (.A1(\wb_dat_o[8] ),
    .A2(_03635_),
    .B1(_03634_),
    .B2(\u_uart2wb.reg_rdata[8] ),
    .X(_00745_));
 sky130_fd_sc_hd__a22o_1 _08023_ (.A1(\wb_dat_o[9] ),
    .A2(_03635_),
    .B1(_03634_),
    .B2(_03068_),
    .X(_00746_));
 sky130_fd_sc_hd__a22o_1 _08024_ (.A1(\wb_dat_o[10] ),
    .A2(_03635_),
    .B1(_03634_),
    .B2(_03066_),
    .X(_00747_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08025_ (.A(_03631_),
    .X(_03636_));
 sky130_fd_sc_hd__a22o_1 _08026_ (.A1(\wb_dat_o[11] ),
    .A2(_03635_),
    .B1(_03636_),
    .B2(\u_uart2wb.reg_rdata[11] ),
    .X(_00748_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08027_ (.A(_03619_),
    .X(_03637_));
 sky130_fd_sc_hd__a22o_1 _08028_ (.A1(\wb_dat_o[12] ),
    .A2(_03637_),
    .B1(_03636_),
    .B2(\u_uart2wb.reg_rdata[12] ),
    .X(_00749_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08029_ (.A(\u_uart2wb.reg_rdata[13] ),
    .X(_03638_));
 sky130_fd_sc_hd__a22o_1 _08030_ (.A1(\wb_dat_o[13] ),
    .A2(_03637_),
    .B1(_03636_),
    .B2(_03638_),
    .X(_00750_));
 sky130_fd_sc_hd__a22o_1 _08031_ (.A1(\wb_dat_o[14] ),
    .A2(_03637_),
    .B1(_03636_),
    .B2(\u_uart2wb.reg_rdata[14] ),
    .X(_00751_));
 sky130_fd_sc_hd__clkbuf_2 _08032_ (.A(_03627_),
    .X(_03639_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08033_ (.A(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__a22o_1 _08034_ (.A1(\wb_dat_o[15] ),
    .A2(_03637_),
    .B1(_03640_),
    .B2(\u_uart2wb.reg_rdata[15] ),
    .X(_00752_));
 sky130_fd_sc_hd__clkbuf_2 _08035_ (.A(_03618_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _08036_ (.A(_03641_),
    .X(_03642_));
 sky130_fd_sc_hd__a22o_1 _08037_ (.A1(\wb_dat_o[16] ),
    .A2(_03642_),
    .B1(_03640_),
    .B2(\u_uart2wb.reg_rdata[16] ),
    .X(_00753_));
 sky130_fd_sc_hd__a22o_1 _08038_ (.A1(\wb_dat_o[17] ),
    .A2(_03642_),
    .B1(_03640_),
    .B2(_03100_),
    .X(_00754_));
 sky130_fd_sc_hd__a22o_1 _08039_ (.A1(\wb_dat_o[18] ),
    .A2(_03642_),
    .B1(_03640_),
    .B2(_03099_),
    .X(_00755_));
 sky130_fd_sc_hd__clkbuf_1 _08040_ (.A(_03639_),
    .X(_03643_));
 sky130_fd_sc_hd__a22o_1 _08041_ (.A1(\wb_dat_o[19] ),
    .A2(_03642_),
    .B1(_03643_),
    .B2(\u_uart2wb.reg_rdata[19] ),
    .X(_00756_));
 sky130_fd_sc_hd__clkbuf_1 _08042_ (.A(_03641_),
    .X(_03644_));
 sky130_fd_sc_hd__a22o_1 _08043_ (.A1(\wb_dat_o[20] ),
    .A2(_03644_),
    .B1(_03643_),
    .B2(\u_uart2wb.reg_rdata[20] ),
    .X(_00757_));
 sky130_fd_sc_hd__a22o_1 _08044_ (.A1(\wb_dat_o[21] ),
    .A2(_03644_),
    .B1(_03643_),
    .B2(_03129_),
    .X(_00758_));
 sky130_fd_sc_hd__a22o_1 _08045_ (.A1(\wb_dat_o[22] ),
    .A2(_03644_),
    .B1(_03643_),
    .B2(_03128_),
    .X(_00759_));
 sky130_fd_sc_hd__clkbuf_1 _08046_ (.A(_03639_),
    .X(_03645_));
 sky130_fd_sc_hd__a22o_1 _08047_ (.A1(\wb_dat_o[23] ),
    .A2(_03644_),
    .B1(_03645_),
    .B2(\u_uart2wb.reg_rdata[23] ),
    .X(_00760_));
 sky130_fd_sc_hd__clkbuf_1 _08048_ (.A(_03641_),
    .X(_03646_));
 sky130_fd_sc_hd__a22o_1 _08049_ (.A1(\wb_dat_o[24] ),
    .A2(_03646_),
    .B1(_03645_),
    .B2(\u_uart2wb.reg_rdata[24] ),
    .X(_00761_));
 sky130_fd_sc_hd__a22o_1 _08050_ (.A1(\wb_dat_o[25] ),
    .A2(_03646_),
    .B1(_03645_),
    .B2(_03158_),
    .X(_00762_));
 sky130_fd_sc_hd__a22o_1 _08051_ (.A1(\wb_dat_o[26] ),
    .A2(_03646_),
    .B1(_03645_),
    .B2(_03157_),
    .X(_00763_));
 sky130_fd_sc_hd__clkbuf_1 _08052_ (.A(_03639_),
    .X(_03647_));
 sky130_fd_sc_hd__a22o_1 _08053_ (.A1(\wb_dat_o[27] ),
    .A2(_03646_),
    .B1(_03647_),
    .B2(\u_uart2wb.reg_rdata[27] ),
    .X(_00764_));
 sky130_fd_sc_hd__clkbuf_1 _08054_ (.A(_03641_),
    .X(_03648_));
 sky130_fd_sc_hd__a22o_1 _08055_ (.A1(\wb_dat_o[28] ),
    .A2(_03648_),
    .B1(_03647_),
    .B2(\u_uart2wb.reg_rdata[28] ),
    .X(_00765_));
 sky130_fd_sc_hd__a22o_1 _08056_ (.A1(\wb_dat_o[29] ),
    .A2(_03648_),
    .B1(_03647_),
    .B2(_03000_),
    .X(_00766_));
 sky130_fd_sc_hd__a22o_1 _08057_ (.A1(\wb_dat_o[30] ),
    .A2(_03648_),
    .B1(_03647_),
    .B2(\u_uart2wb.reg_rdata[30] ),
    .X(_00767_));
 sky130_fd_sc_hd__a22o_1 _08058_ (.A1(\wb_dat_o[31] ),
    .A2(_03648_),
    .B1(_03631_),
    .B2(_02985_),
    .X(_00768_));
 sky130_fd_sc_hd__and2_1 _08059_ (.A(_03617_),
    .B(_03625_),
    .X(_03649_));
 sky130_fd_sc_hd__o21a_1 _08060_ (.A1(\u_uart2wb.reg_ack ),
    .A2(_03649_),
    .B1(_03626_),
    .X(_00769_));
 sky130_fd_sc_hd__or2b_1 _08061_ (.A(_03621_),
    .B_N(_03626_),
    .X(_03650_));
 sky130_fd_sc_hd__clkbuf_1 _08062_ (.A(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__or3b_1 _08063_ (.A(_03626_),
    .B(_03621_),
    .C_N(\u_uart2wb.reg_req ),
    .X(_03652_));
 sky130_fd_sc_hd__o21ai_1 _08064_ (.A1(_03651_),
    .A2(_03625_),
    .B1(_03652_),
    .Y(_00770_));
 sky130_fd_sc_hd__and2b_1 _08065_ (.A_N(\u_uart2wb.u_async_reg_bus.in_state[0] ),
    .B(_03621_),
    .X(_03653_));
 sky130_fd_sc_hd__o21a_1 _08066_ (.A1(_03617_),
    .A2(_03653_),
    .B1(\u_uart2wb.u_async_reg_bus.out_flag_ss ),
    .X(_00771_));
 sky130_fd_sc_hd__clkbuf_1 _08067_ (.A(\u_uart2wb.u_async_reg_bus.in_timer[0] ),
    .X(_03654_));
 sky130_fd_sc_hd__nor2_1 _08068_ (.A(_03650_),
    .B(_03625_),
    .Y(_03655_));
 sky130_fd_sc_hd__nor2_1 _08069_ (.A(_03649_),
    .B(_03653_),
    .Y(_03656_));
 sky130_fd_sc_hd__clkbuf_1 _08070_ (.A(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__clkbuf_1 _08071_ (.A(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__nand2_1 _08072_ (.A(_03654_),
    .B(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__o21a_1 _08073_ (.A1(_03654_),
    .A2(_03655_),
    .B1(_03659_),
    .X(_00772_));
 sky130_fd_sc_hd__clkbuf_1 _08074_ (.A(\u_uart2wb.u_async_reg_bus.in_timer[1] ),
    .X(_03660_));
 sky130_fd_sc_hd__inv_2 _08075_ (.A(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__a21o_1 _08076_ (.A1(_03660_),
    .A2(\u_uart2wb.u_async_reg_bus.in_timer[0] ),
    .B1(_03650_),
    .X(_03662_));
 sky130_fd_sc_hd__nand2_1 _08077_ (.A(_03657_),
    .B(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__a21boi_1 _08078_ (.A1(_03661_),
    .A2(_03659_),
    .B1_N(_03663_),
    .Y(_00773_));
 sky130_fd_sc_hd__and3_1 _08079_ (.A(_03660_),
    .B(_03654_),
    .C(_03655_),
    .X(_03664_));
 sky130_fd_sc_hd__mux2_1 _08080_ (.A0(_03664_),
    .A1(_03663_),
    .S(\u_uart2wb.u_async_reg_bus.in_timer[2] ),
    .X(_03665_));
 sky130_fd_sc_hd__clkbuf_1 _08081_ (.A(_03665_),
    .X(_00774_));
 sky130_fd_sc_hd__a41o_1 _08082_ (.A1(_03660_),
    .A2(_03654_),
    .A3(\u_uart2wb.u_async_reg_bus.in_timer[2] ),
    .A4(_03656_),
    .B1(\u_uart2wb.u_async_reg_bus.in_timer[3] ),
    .X(_03666_));
 sky130_fd_sc_hd__o21ai_1 _08083_ (.A1(_03651_),
    .A2(_03622_),
    .B1(_03657_),
    .Y(_03667_));
 sky130_fd_sc_hd__and2_1 _08084_ (.A(_03666_),
    .B(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__clkbuf_1 _08085_ (.A(_03668_),
    .X(_00775_));
 sky130_fd_sc_hd__and2_1 _08086_ (.A(_03622_),
    .B(_03655_),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_1 _08087_ (.A0(_03669_),
    .A1(_03667_),
    .S(\u_uart2wb.u_async_reg_bus.in_timer[4] ),
    .X(_03670_));
 sky130_fd_sc_hd__clkbuf_1 _08088_ (.A(_03670_),
    .X(_00776_));
 sky130_fd_sc_hd__o21ai_1 _08089_ (.A1(_03651_),
    .A2(_03623_),
    .B1(_03657_),
    .Y(_03671_));
 sky130_fd_sc_hd__a31o_1 _08090_ (.A1(\u_uart2wb.u_async_reg_bus.in_timer[4] ),
    .A2(_03622_),
    .A3(_03656_),
    .B1(\u_uart2wb.u_async_reg_bus.in_timer[5] ),
    .X(_03672_));
 sky130_fd_sc_hd__and2_1 _08091_ (.A(_03671_),
    .B(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__clkbuf_1 _08092_ (.A(_03673_),
    .X(_00777_));
 sky130_fd_sc_hd__and2_1 _08093_ (.A(_03623_),
    .B(_03655_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _08094_ (.A0(_03674_),
    .A1(_03671_),
    .S(\u_uart2wb.u_async_reg_bus.in_timer[6] ),
    .X(_03675_));
 sky130_fd_sc_hd__clkbuf_1 _08095_ (.A(_03675_),
    .X(_00778_));
 sky130_fd_sc_hd__a31o_1 _08096_ (.A1(\u_uart2wb.u_async_reg_bus.in_timer[7] ),
    .A2(\u_uart2wb.u_async_reg_bus.in_timer[6] ),
    .A3(_03623_),
    .B1(_03651_),
    .X(_03676_));
 sky130_fd_sc_hd__a21oi_1 _08097_ (.A1(_03624_),
    .A2(_03658_),
    .B1(\u_uart2wb.u_async_reg_bus.in_timer[7] ),
    .Y(_03677_));
 sky130_fd_sc_hd__a21oi_1 _08098_ (.A1(_03658_),
    .A2(_03676_),
    .B1(_03677_),
    .Y(_00779_));
 sky130_fd_sc_hd__a31o_1 _08099_ (.A1(\u_uart2wb.u_async_reg_bus.in_timer[7] ),
    .A2(_03624_),
    .A3(_03658_),
    .B1(\u_uart2wb.u_async_reg_bus.in_timer[8] ),
    .X(_03678_));
 sky130_fd_sc_hd__o21a_1 _08100_ (.A1(_03617_),
    .A2(_03653_),
    .B1(_03678_),
    .X(_00780_));
 sky130_fd_sc_hd__a21bo_1 _08101_ (.A1(\u_uart2wb.u_async_reg_bus.in_flag ),
    .A2(_03628_),
    .B1_N(_03652_),
    .X(_00781_));
 sky130_fd_sc_hd__inv_2 _08102_ (.A(\u_uart2wb.u_async_reg_bus.out_state[0] ),
    .Y(_03679_));
 sky130_fd_sc_hd__a21oi_1 _08103_ (.A1(_01511_),
    .A2(_03264_),
    .B1(\u_uart2wb.u_async_reg_bus.out_state[1] ),
    .Y(_03680_));
 sky130_fd_sc_hd__or3b_1 _08104_ (.A(\u_uart2wb.u_async_reg_bus.out_state[0] ),
    .B(\u_uart2wb.u_async_reg_bus.out_state[1] ),
    .C_N(\u_uart2wb.u_async_reg_bus.in_flag_ss ),
    .X(_03681_));
 sky130_fd_sc_hd__or2b_1 _08105_ (.A(\u_uart2wb.u_async_reg_bus.out_reg_cs ),
    .B_N(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__o21a_1 _08106_ (.A1(_03679_),
    .A2(_03680_),
    .B1(_03682_),
    .X(_00782_));
 sky130_fd_sc_hd__a21bo_1 _08107_ (.A1(\u_uart2wb.u_async_reg_bus.out_state[0] ),
    .A2(_03680_),
    .B1_N(_03681_),
    .X(_00783_));
 sky130_fd_sc_hd__nor2_1 _08108_ (.A(_03679_),
    .B(\u_uart2wb.u_async_reg_bus.out_state[1] ),
    .Y(_03683_));
 sky130_fd_sc_hd__and3_1 _08109_ (.A(_01511_),
    .B(_03234_),
    .C(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__and3_1 _08110_ (.A(_03679_),
    .B(\u_uart2wb.u_async_reg_bus.out_state[1] ),
    .C(\u_uart2wb.u_async_reg_bus.in_flag_ss ),
    .X(_03685_));
 sky130_fd_sc_hd__or2_1 _08111_ (.A(_03684_),
    .B(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__clkbuf_1 _08112_ (.A(_03686_),
    .X(_00784_));
 sky130_fd_sc_hd__or2_1 _08113_ (.A(\u_uart2wb.auto_rx_enb ),
    .B(\u_uart2wb.u_aut_det.state[7] ),
    .X(_03687_));
 sky130_fd_sc_hd__clkbuf_1 _08114_ (.A(_03687_),
    .X(_00785_));
 sky130_fd_sc_hd__clkbuf_1 _08115_ (.A(\u_uart2wb.u_aut_det.clk_cnt[0] ),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _08116_ (.A0(\u_uart2wb.u_aut_det.ref1_cnt[0] ),
    .A1(_03688_),
    .S(_01180_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_1 _08117_ (.A(_03689_),
    .X(_00786_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08118_ (.A(\u_uart2wb.u_aut_det.clk_cnt[1] ),
    .X(_03690_));
 sky130_fd_sc_hd__mux2_1 _08119_ (.A0(_01193_),
    .A1(_03690_),
    .S(_01180_),
    .X(_03691_));
 sky130_fd_sc_hd__clkbuf_1 _08120_ (.A(_03691_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _08121_ (.A0(\u_uart2wb.u_aut_det.ref1_cnt[2] ),
    .A1(\u_uart2wb.u_aut_det.clk_cnt[2] ),
    .S(_01180_),
    .X(_03692_));
 sky130_fd_sc_hd__clkbuf_1 _08122_ (.A(_03692_),
    .X(_00788_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08123_ (.A(\u_uart2wb.u_aut_det.clk_cnt[3] ),
    .X(_03693_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08124_ (.A(_01179_),
    .X(_03694_));
 sky130_fd_sc_hd__clkbuf_2 _08125_ (.A(_03694_),
    .X(_03695_));
 sky130_fd_sc_hd__mux2_1 _08126_ (.A0(_01200_),
    .A1(_03693_),
    .S(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__clkbuf_1 _08127_ (.A(_03696_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _08128_ (.A0(_01222_),
    .A1(\u_uart2wb.u_aut_det.clk_cnt[4] ),
    .S(_03695_),
    .X(_03697_));
 sky130_fd_sc_hd__clkbuf_1 _08129_ (.A(_03697_),
    .X(_00790_));
 sky130_fd_sc_hd__clkbuf_1 _08130_ (.A(\u_uart2wb.u_aut_det.clk_cnt[5] ),
    .X(_03698_));
 sky130_fd_sc_hd__mux2_1 _08131_ (.A0(_01219_),
    .A1(_03698_),
    .S(_03695_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_1 _08132_ (.A(_03699_),
    .X(_00791_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08133_ (.A(\u_uart2wb.u_aut_det.clk_cnt[6] ),
    .X(_03700_));
 sky130_fd_sc_hd__mux2_1 _08134_ (.A0(_01229_),
    .A1(_03700_),
    .S(_03695_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_1 _08135_ (.A(_03701_),
    .X(_00792_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08136_ (.A(\u_uart2wb.u_aut_det.clk_cnt[7] ),
    .X(_03702_));
 sky130_fd_sc_hd__buf_2 _08137_ (.A(_03694_),
    .X(_03703_));
 sky130_fd_sc_hd__mux2_1 _08138_ (.A0(\u_uart2wb.u_aut_det.ref1_cnt[7] ),
    .A1(_03702_),
    .S(_03703_),
    .X(_03704_));
 sky130_fd_sc_hd__clkbuf_1 _08139_ (.A(_03704_),
    .X(_00793_));
 sky130_fd_sc_hd__clkbuf_2 _08140_ (.A(\u_uart2wb.u_aut_det.clk_cnt[8] ),
    .X(_03705_));
 sky130_fd_sc_hd__mux2_1 _08141_ (.A0(_01332_),
    .A1(_03705_),
    .S(_03703_),
    .X(_03706_));
 sky130_fd_sc_hd__clkbuf_1 _08142_ (.A(_03706_),
    .X(_00794_));
 sky130_fd_sc_hd__clkbuf_2 _08143_ (.A(\u_uart2wb.u_aut_det.clk_cnt[9] ),
    .X(_03707_));
 sky130_fd_sc_hd__mux2_1 _08144_ (.A0(_01246_),
    .A1(_03707_),
    .S(_03703_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_1 _08145_ (.A(_03708_),
    .X(_00795_));
 sky130_fd_sc_hd__clkbuf_2 _08146_ (.A(\u_uart2wb.u_aut_det.clk_cnt[10] ),
    .X(_03709_));
 sky130_fd_sc_hd__mux2_1 _08147_ (.A0(\u_uart2wb.u_aut_det.ref1_cnt[10] ),
    .A1(_03709_),
    .S(_03703_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_1 _08148_ (.A(_03710_),
    .X(_00796_));
 sky130_fd_sc_hd__clkbuf_2 _08149_ (.A(\u_uart2wb.u_aut_det.clk_cnt[11] ),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_2 _08150_ (.A(_03694_),
    .X(_03712_));
 sky130_fd_sc_hd__mux2_1 _08151_ (.A0(\u_uart2wb.u_aut_det.ref1_cnt[11] ),
    .A1(_03711_),
    .S(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_1 _08152_ (.A(_03713_),
    .X(_00797_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08153_ (.A(\u_uart2wb.u_aut_det.clk_cnt[12] ),
    .X(_03714_));
 sky130_fd_sc_hd__mux2_1 _08154_ (.A0(_01235_),
    .A1(_03714_),
    .S(_03712_),
    .X(_03715_));
 sky130_fd_sc_hd__clkbuf_1 _08155_ (.A(_03715_),
    .X(_00798_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08156_ (.A(\u_uart2wb.u_aut_det.clk_cnt[13] ),
    .X(_03716_));
 sky130_fd_sc_hd__mux2_1 _08157_ (.A0(_01273_),
    .A1(_03716_),
    .S(_03712_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_1 _08158_ (.A(_03717_),
    .X(_00799_));
 sky130_fd_sc_hd__clkbuf_1 _08159_ (.A(\u_uart2wb.u_aut_det.clk_cnt[14] ),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_2 _08160_ (.A(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__mux2_1 _08161_ (.A0(\u_uart2wb.u_aut_det.ref1_cnt[14] ),
    .A1(_03719_),
    .S(_03712_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _08162_ (.A(_03720_),
    .X(_00800_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08163_ (.A(\u_uart2wb.u_aut_det.clk_cnt[15] ),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_2 _08164_ (.A(_01179_),
    .X(_03722_));
 sky130_fd_sc_hd__mux2_1 _08165_ (.A0(_01269_),
    .A1(_03721_),
    .S(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_1 _08166_ (.A(_03723_),
    .X(_00801_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08167_ (.A(\u_uart2wb.u_aut_det.clk_cnt[16] ),
    .X(_03724_));
 sky130_fd_sc_hd__mux2_1 _08168_ (.A0(_01340_),
    .A1(_03724_),
    .S(_03722_),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_1 _08169_ (.A(_03725_),
    .X(_00802_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08170_ (.A(\u_uart2wb.u_aut_det.clk_cnt[17] ),
    .X(_03726_));
 sky130_fd_sc_hd__mux2_1 _08171_ (.A0(\u_uart2wb.u_aut_det.ref1_cnt[17] ),
    .A1(_03726_),
    .S(_03722_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_1 _08172_ (.A(_03727_),
    .X(_00803_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08173_ (.A(\u_uart2wb.u_aut_det.clk_cnt[18] ),
    .X(_03728_));
 sky130_fd_sc_hd__mux2_1 _08174_ (.A0(_01283_),
    .A1(_03728_),
    .S(_03722_),
    .X(_03729_));
 sky130_fd_sc_hd__clkbuf_1 _08175_ (.A(_03729_),
    .X(_00804_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08176_ (.A(\u_uart2wb.u_aut_det.clk_cnt[19] ),
    .X(_03730_));
 sky130_fd_sc_hd__mux2_1 _08177_ (.A0(\u_uart2wb.u_aut_det.ref1_cnt[19] ),
    .A1(_03730_),
    .S(_03694_),
    .X(_03731_));
 sky130_fd_sc_hd__clkbuf_1 _08178_ (.A(_03731_),
    .X(_00805_));
 sky130_fd_sc_hd__o22a_1 _08179_ (.A1(\u_uart2wb.u_async_reg_bus.out_flag ),
    .A2(_03684_),
    .B1(_03685_),
    .B2(_03683_),
    .X(_00806_));
 sky130_fd_sc_hd__or3_1 _08180_ (.A(\u_uart2wb.u_aut_det.state[0] ),
    .B(_01443_),
    .C(_01445_),
    .X(_03732_));
 sky130_fd_sc_hd__or3b_1 _08181_ (.A(_01182_),
    .B(_01447_),
    .C_N(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__nor2_1 _08182_ (.A(_01441_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08183_ (.A(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__or2_1 _08184_ (.A(\u_uart2wb.u_aut_det.clk_cnt[0] ),
    .B(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__clkbuf_1 _08185_ (.A(_03733_),
    .X(_03737_));
 sky130_fd_sc_hd__a221o_1 _08186_ (.A1(_01439_),
    .A2(_01443_),
    .B1(_01444_),
    .B2(_01165_),
    .C1(\u_uart2wb.u_aut_det.state[3] ),
    .X(_03738_));
 sky130_fd_sc_hd__or2_1 _08187_ (.A(_03737_),
    .B(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08188_ (.A(_03734_),
    .X(_03740_));
 sky130_fd_sc_hd__nand2_1 _08189_ (.A(_03688_),
    .B(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__and3_1 _08190_ (.A(_03736_),
    .B(_03739_),
    .C(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__clkbuf_1 _08191_ (.A(_03742_),
    .X(_00807_));
 sky130_fd_sc_hd__inv_2 _08192_ (.A(_03690_),
    .Y(_03743_));
 sky130_fd_sc_hd__nor3b_1 _08193_ (.A(_01182_),
    .B(_01447_),
    .C_N(_03732_),
    .Y(_03744_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08194_ (.A(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08195_ (.A(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__a21o_1 _08196_ (.A1(_03688_),
    .A2(_03746_),
    .B1(_03690_),
    .X(_03747_));
 sky130_fd_sc_hd__clkbuf_1 _08197_ (.A(_03739_),
    .X(_03748_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08198_ (.A(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__o211a_1 _08199_ (.A1(_03743_),
    .A2(_03741_),
    .B1(_03747_),
    .C1(_03749_),
    .X(_00808_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08200_ (.A(_03739_),
    .X(_03750_));
 sky130_fd_sc_hd__a31o_1 _08201_ (.A1(\u_uart2wb.u_aut_det.clk_cnt[1] ),
    .A2(\u_uart2wb.u_aut_det.clk_cnt[0] ),
    .A3(_03735_),
    .B1(\u_uart2wb.u_aut_det.clk_cnt[2] ),
    .X(_03751_));
 sky130_fd_sc_hd__nand2_1 _08202_ (.A(_01168_),
    .B(_03740_),
    .Y(_03752_));
 sky130_fd_sc_hd__and3_1 _08203_ (.A(_03750_),
    .B(_03751_),
    .C(_03752_),
    .X(_03753_));
 sky130_fd_sc_hd__clkbuf_1 _08204_ (.A(_03753_),
    .X(_00809_));
 sky130_fd_sc_hd__inv_2 _08205_ (.A(_03693_),
    .Y(_03754_));
 sky130_fd_sc_hd__a21o_1 _08206_ (.A1(_01168_),
    .A2(_03746_),
    .B1(_03693_),
    .X(_03755_));
 sky130_fd_sc_hd__o211a_1 _08207_ (.A1(_03754_),
    .A2(_03752_),
    .B1(_03755_),
    .C1(_03749_),
    .X(_00810_));
 sky130_fd_sc_hd__a31o_1 _08208_ (.A1(\u_uart2wb.u_aut_det.clk_cnt[3] ),
    .A2(_01168_),
    .A3(_03735_),
    .B1(\u_uart2wb.u_aut_det.clk_cnt[4] ),
    .X(_03756_));
 sky130_fd_sc_hd__clkbuf_1 _08209_ (.A(_01169_),
    .X(_03757_));
 sky130_fd_sc_hd__nand2_1 _08210_ (.A(_03757_),
    .B(_03740_),
    .Y(_03758_));
 sky130_fd_sc_hd__and3_1 _08211_ (.A(_03748_),
    .B(_03756_),
    .C(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_1 _08212_ (.A(_03759_),
    .X(_00811_));
 sky130_fd_sc_hd__nand3_1 _08213_ (.A(_03698_),
    .B(_03757_),
    .C(_03735_),
    .Y(_03760_));
 sky130_fd_sc_hd__a21o_1 _08214_ (.A1(_03757_),
    .A2(_03745_),
    .B1(\u_uart2wb.u_aut_det.clk_cnt[5] ),
    .X(_03761_));
 sky130_fd_sc_hd__and3_1 _08215_ (.A(_03748_),
    .B(_03760_),
    .C(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_1 _08216_ (.A(_03762_),
    .X(_00812_));
 sky130_fd_sc_hd__inv_2 _08217_ (.A(_03700_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand2_1 _08218_ (.A(_03763_),
    .B(_03760_),
    .Y(_03764_));
 sky130_fd_sc_hd__o211a_1 _08219_ (.A1(_03763_),
    .A2(_03760_),
    .B1(_03764_),
    .C1(_03749_),
    .X(_00813_));
 sky130_fd_sc_hd__clkbuf_1 _08220_ (.A(_01170_),
    .X(_03765_));
 sky130_fd_sc_hd__nand2_1 _08221_ (.A(_03765_),
    .B(_01440_),
    .Y(_03766_));
 sky130_fd_sc_hd__and2_1 _08222_ (.A(_03744_),
    .B(_03738_),
    .X(_03767_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08223_ (.A(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__a31o_1 _08224_ (.A1(_03698_),
    .A2(_03700_),
    .A3(_03757_),
    .B1(_03702_),
    .X(_03769_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08225_ (.A(_03737_),
    .X(_03770_));
 sky130_fd_sc_hd__a32o_1 _08226_ (.A1(_03766_),
    .A2(_03768_),
    .A3(_03769_),
    .B1(_03770_),
    .B2(_03702_),
    .X(_00814_));
 sky130_fd_sc_hd__nand2_1 _08227_ (.A(_03705_),
    .B(_03765_),
    .Y(_03771_));
 sky130_fd_sc_hd__a31o_1 _08228_ (.A1(_03765_),
    .A2(_01176_),
    .A3(_03746_),
    .B1(\u_uart2wb.u_aut_det.clk_cnt[8] ),
    .X(_03772_));
 sky130_fd_sc_hd__o311a_1 _08229_ (.A1(_03771_),
    .A2(_01442_),
    .A3(_03737_),
    .B1(_03750_),
    .C1(_03772_),
    .X(_00815_));
 sky130_fd_sc_hd__a21o_1 _08230_ (.A1(_03705_),
    .A2(_03765_),
    .B1(_03707_),
    .X(_03773_));
 sky130_fd_sc_hd__clkbuf_1 _08231_ (.A(_01171_),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_1 _08232_ (.A(_03767_),
    .X(_03775_));
 sky130_fd_sc_hd__a21boi_1 _08233_ (.A1(_03774_),
    .A2(_01440_),
    .B1_N(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__a22o_1 _08234_ (.A1(_03707_),
    .A2(_03770_),
    .B1(_03773_),
    .B2(_03776_),
    .X(_00816_));
 sky130_fd_sc_hd__inv_2 _08235_ (.A(\u_uart2wb.u_aut_det.clk_cnt[10] ),
    .Y(_03777_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08236_ (.A(_03737_),
    .X(_03778_));
 sky130_fd_sc_hd__a31o_1 _08237_ (.A1(_03774_),
    .A2(_01176_),
    .A3(_03775_),
    .B1(_03709_),
    .X(_03779_));
 sky130_fd_sc_hd__o31a_1 _08238_ (.A1(_03777_),
    .A2(_03778_),
    .A3(_03776_),
    .B1(_03779_),
    .X(_00817_));
 sky130_fd_sc_hd__and4_1 _08239_ (.A(_03711_),
    .B(\u_uart2wb.u_aut_det.clk_cnt[10] ),
    .C(_01171_),
    .D(_03744_),
    .X(_03780_));
 sky130_fd_sc_hd__inv_2 _08240_ (.A(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__a31o_1 _08241_ (.A1(_03709_),
    .A2(_03774_),
    .A3(_03746_),
    .B1(_03711_),
    .X(_03782_));
 sky130_fd_sc_hd__o211a_1 _08242_ (.A1(_01442_),
    .A2(_03781_),
    .B1(_03782_),
    .C1(_03749_),
    .X(_00818_));
 sky130_fd_sc_hd__or3_1 _08243_ (.A(_03714_),
    .B(_01441_),
    .C(_03781_),
    .X(_03783_));
 sky130_fd_sc_hd__o21ai_1 _08244_ (.A1(_01442_),
    .A2(_03781_),
    .B1(_03714_),
    .Y(_03784_));
 sky130_fd_sc_hd__a21boi_1 _08245_ (.A1(_03783_),
    .A2(_03784_),
    .B1_N(_03750_),
    .Y(_00819_));
 sky130_fd_sc_hd__a21o_1 _08246_ (.A1(_03774_),
    .A2(_01172_),
    .B1(_03716_),
    .X(_03785_));
 sky130_fd_sc_hd__clkbuf_1 _08247_ (.A(_01173_),
    .X(_03786_));
 sky130_fd_sc_hd__a21boi_1 _08248_ (.A1(_03786_),
    .A2(_01440_),
    .B1_N(_03775_),
    .Y(_03787_));
 sky130_fd_sc_hd__a22o_1 _08249_ (.A1(_03716_),
    .A2(_03770_),
    .B1(_03785_),
    .B2(_03787_),
    .X(_00820_));
 sky130_fd_sc_hd__inv_2 _08250_ (.A(_03719_),
    .Y(_03788_));
 sky130_fd_sc_hd__a31o_1 _08251_ (.A1(_03786_),
    .A2(_01176_),
    .A3(_03775_),
    .B1(_03719_),
    .X(_03789_));
 sky130_fd_sc_hd__o31a_1 _08252_ (.A1(_03788_),
    .A2(_03778_),
    .A3(_03787_),
    .B1(_03789_),
    .X(_00821_));
 sky130_fd_sc_hd__nand4_1 _08253_ (.A(_03721_),
    .B(_03718_),
    .C(_03786_),
    .D(_03740_),
    .Y(_03790_));
 sky130_fd_sc_hd__a31o_1 _08254_ (.A1(_03718_),
    .A2(_01173_),
    .A3(_03745_),
    .B1(\u_uart2wb.u_aut_det.clk_cnt[15] ),
    .X(_03791_));
 sky130_fd_sc_hd__and3_1 _08255_ (.A(_03748_),
    .B(_03790_),
    .C(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__clkbuf_1 _08256_ (.A(_03792_),
    .X(_00822_));
 sky130_fd_sc_hd__clkbuf_1 _08257_ (.A(\u_uart2wb.u_aut_det.clk_cnt[17] ),
    .X(_03793_));
 sky130_fd_sc_hd__clkbuf_1 _08258_ (.A(_01174_),
    .X(_03794_));
 sky130_fd_sc_hd__a21bo_1 _08259_ (.A1(_03793_),
    .A2(_01167_),
    .B1_N(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__a31o_1 _08260_ (.A1(_03721_),
    .A2(_03718_),
    .A3(_03786_),
    .B1(_03724_),
    .X(_03796_));
 sky130_fd_sc_hd__a32o_1 _08261_ (.A1(_03768_),
    .A2(_03795_),
    .A3(_03796_),
    .B1(_03770_),
    .B2(_03724_),
    .X(_00823_));
 sky130_fd_sc_hd__nand2_1 _08262_ (.A(_03793_),
    .B(_01174_),
    .Y(_03797_));
 sky130_fd_sc_hd__or2_1 _08263_ (.A(_01167_),
    .B(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__or2_1 _08264_ (.A(_03793_),
    .B(_03794_),
    .X(_03799_));
 sky130_fd_sc_hd__a32o_1 _08265_ (.A1(_03768_),
    .A2(_03798_),
    .A3(_03799_),
    .B1(_03778_),
    .B2(_03726_),
    .X(_00824_));
 sky130_fd_sc_hd__a21o_1 _08266_ (.A1(_03726_),
    .A2(_03794_),
    .B1(_03728_),
    .X(_03800_));
 sky130_fd_sc_hd__or3b_1 _08267_ (.A(_03730_),
    .B(_03797_),
    .C_N(\u_uart2wb.u_aut_det.clk_cnt[18] ),
    .X(_03801_));
 sky130_fd_sc_hd__a32o_1 _08268_ (.A1(_03768_),
    .A2(_03800_),
    .A3(_03801_),
    .B1(_03778_),
    .B2(_03728_),
    .X(_00825_));
 sky130_fd_sc_hd__a41o_1 _08269_ (.A1(_03793_),
    .A2(\u_uart2wb.u_aut_det.clk_cnt[18] ),
    .A3(_03794_),
    .A4(_03745_),
    .B1(_03730_),
    .X(_03802_));
 sky130_fd_sc_hd__and2_1 _08270_ (.A(_03750_),
    .B(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__clkbuf_1 _08271_ (.A(_03803_),
    .X(_00826_));
 sky130_fd_sc_hd__nand2_1 _08272_ (.A(\u_uart2wb.u_aut_det.state[5] ),
    .B(_01433_),
    .Y(_03804_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08273_ (.A(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__and3_1 _08274_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[4] ),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[4] ),
    .C(_01216_),
    .X(_03806_));
 sky130_fd_sc_hd__a21oi_1 _08275_ (.A1(_01220_),
    .A2(_01219_),
    .B1(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__a22o_1 _08276_ (.A1(\u_uart2wb.u_aut_det.ref2_cnt[1] ),
    .A2(\u_uart2wb.u_aut_det.ref1_cnt[1] ),
    .B1(\u_uart2wb.u_aut_det.ref2_cnt[0] ),
    .B2(\u_uart2wb.u_aut_det.ref1_cnt[0] ),
    .X(_03808_));
 sky130_fd_sc_hd__o2111ai_2 _08277_ (.A1(_01194_),
    .A2(_01193_),
    .B1(_01190_),
    .C1(_01191_),
    .D1(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__and2_1 _08278_ (.A(_01201_),
    .B(_01200_),
    .X(_03810_));
 sky130_fd_sc_hd__a31oi_2 _08279_ (.A1(_01198_),
    .A2(\u_uart2wb.u_aut_det.ref1_cnt[2] ),
    .A3(_01190_),
    .B1(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__a211o_1 _08280_ (.A1(_03809_),
    .A2(_03811_),
    .B1(_01396_),
    .C1(_01188_),
    .X(_03812_));
 sky130_fd_sc_hd__a211o_1 _08281_ (.A1(_03807_),
    .A2(_03812_),
    .B1(_01212_),
    .C1(_01213_),
    .X(_03813_));
 sky130_fd_sc_hd__clkbuf_1 _08282_ (.A(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__and3b_1 _08283_ (.A_N(_01212_),
    .B(_01229_),
    .C(\u_uart2wb.u_aut_det.ref2_cnt[6] ),
    .X(_03815_));
 sky130_fd_sc_hd__a21oi_2 _08284_ (.A1(\u_uart2wb.u_aut_det.ref2_cnt[7] ),
    .A2(\u_uart2wb.u_aut_det.ref1_cnt[7] ),
    .B1(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__a211o_1 _08285_ (.A1(_03814_),
    .A2(_03816_),
    .B1(_01346_),
    .C1(_01247_),
    .X(_03817_));
 sky130_fd_sc_hd__or2_1 _08286_ (.A(_01241_),
    .B(_01376_),
    .X(_03818_));
 sky130_fd_sc_hd__nand3_1 _08287_ (.A(_01331_),
    .B(_01332_),
    .C(_01324_),
    .Y(_03819_));
 sky130_fd_sc_hd__a21boi_1 _08288_ (.A1(_01245_),
    .A2(_01246_),
    .B1_N(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__nand2_1 _08289_ (.A(_01335_),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[10] ),
    .Y(_03821_));
 sky130_fd_sc_hd__o21a_1 _08290_ (.A1(_01376_),
    .A2(_03820_),
    .B1(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__nand2_1 _08291_ (.A(_01256_),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[11] ),
    .Y(_03823_));
 sky130_fd_sc_hd__o221a_2 _08292_ (.A1(_03817_),
    .A2(_03818_),
    .B1(_03822_),
    .B2(_01423_),
    .C1(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__nand2_1 _08293_ (.A(_01251_),
    .B(_01234_),
    .Y(_03825_));
 sky130_fd_sc_hd__or4_1 _08294_ (.A(_01321_),
    .B(_01411_),
    .C(_03824_),
    .D(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__nand2_1 _08295_ (.A(_01268_),
    .B(_01269_),
    .Y(_03827_));
 sky130_fd_sc_hd__nand2_1 _08296_ (.A(_01359_),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[14] ),
    .Y(_03828_));
 sky130_fd_sc_hd__nand2_1 _08297_ (.A(_01355_),
    .B(_01235_),
    .Y(_03829_));
 sky130_fd_sc_hd__nand2_1 _08298_ (.A(_01274_),
    .B(_01273_),
    .Y(_03830_));
 sky130_fd_sc_hd__o21ai_1 _08299_ (.A1(_01254_),
    .A2(_03829_),
    .B1(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand2_1 _08300_ (.A(_01251_),
    .B(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__a21o_1 _08301_ (.A1(_03828_),
    .A2(_03832_),
    .B1(_01271_),
    .X(_03833_));
 sky130_fd_sc_hd__and3_1 _08302_ (.A(_03826_),
    .B(_03827_),
    .C(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__xnor2_1 _08303_ (.A(_01342_),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__inv_2 _08304_ (.A(_03831_),
    .Y(_03836_));
 sky130_fd_sc_hd__o31a_1 _08305_ (.A1(_01321_),
    .A2(_01411_),
    .A3(_03824_),
    .B1(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__xnor2_1 _08306_ (.A(_01415_),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__a21o_1 _08307_ (.A1(_03817_),
    .A2(_03820_),
    .B1(_01377_),
    .X(_03839_));
 sky130_fd_sc_hd__clkbuf_1 _08308_ (.A(_03839_),
    .X(_03840_));
 sky130_fd_sc_hd__a21boi_1 _08309_ (.A1(_03821_),
    .A2(_03840_),
    .B1_N(_01423_),
    .Y(_03841_));
 sky130_fd_sc_hd__and3b_1 _08310_ (.A_N(_01423_),
    .B(_03821_),
    .C(_03839_),
    .X(_03842_));
 sky130_fd_sc_hd__o21a_1 _08311_ (.A1(_01321_),
    .A2(_03824_),
    .B1(_03829_),
    .X(_03843_));
 sky130_fd_sc_hd__xnor2_1 _08312_ (.A(_01238_),
    .B(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand3_1 _08313_ (.A(_01377_),
    .B(_03817_),
    .C(_03820_),
    .Y(_03845_));
 sky130_fd_sc_hd__a21oi_1 _08314_ (.A1(_03814_),
    .A2(_03816_),
    .B1(_01346_),
    .Y(_03846_));
 sky130_fd_sc_hd__a21o_1 _08315_ (.A1(_01331_),
    .A2(_01332_),
    .B1(_01324_),
    .X(_03847_));
 sky130_fd_sc_hd__o211a_1 _08316_ (.A1(_03846_),
    .A2(_03847_),
    .B1(_03819_),
    .C1(_03817_),
    .X(_03848_));
 sky130_fd_sc_hd__a21o_1 _08317_ (.A1(_03814_),
    .A2(_03816_),
    .B1(_01346_),
    .X(_03849_));
 sky130_fd_sc_hd__nand3_1 _08318_ (.A(_01347_),
    .B(_03814_),
    .C(_03816_),
    .Y(_03850_));
 sky130_fd_sc_hd__and2_1 _08319_ (.A(_03849_),
    .B(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__a21oi_1 _08320_ (.A1(_03807_),
    .A2(_03812_),
    .B1(_01313_),
    .Y(_03852_));
 sky130_fd_sc_hd__o21ai_1 _08321_ (.A1(_01317_),
    .A2(_01230_),
    .B1(_01225_),
    .Y(_03853_));
 sky130_fd_sc_hd__inv_2 _08322_ (.A(_03815_),
    .Y(_03854_));
 sky130_fd_sc_hd__o211a_1 _08323_ (.A1(_03852_),
    .A2(_03853_),
    .B1(_03813_),
    .C1(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__o21a_1 _08324_ (.A1(_01282_),
    .A2(_01283_),
    .B1(_01395_),
    .X(_03856_));
 sky130_fd_sc_hd__and3_1 _08325_ (.A(_01313_),
    .B(_03807_),
    .C(_03812_),
    .X(_03857_));
 sky130_fd_sc_hd__nor2_1 _08326_ (.A(_03852_),
    .B(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__or3_1 _08327_ (.A(\u_uart2wb.u_aut_det.ref2_cnt[16] ),
    .B(_01289_),
    .C(_01291_),
    .X(_03859_));
 sky130_fd_sc_hd__o21ai_1 _08328_ (.A1(_01288_),
    .A2(_01289_),
    .B1(_01292_),
    .Y(_03860_));
 sky130_fd_sc_hd__o311a_1 _08329_ (.A1(_01282_),
    .A2(_01283_),
    .A3(_01395_),
    .B1(_03859_),
    .C1(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__or4b_1 _08330_ (.A(_03855_),
    .B(_03856_),
    .C(_03858_),
    .D_N(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__or3_1 _08331_ (.A(_03848_),
    .B(_03851_),
    .C(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__xnor2_2 _08332_ (.A(_01236_),
    .B(_03824_),
    .Y(_03864_));
 sky130_fd_sc_hd__a211o_1 _08333_ (.A1(_03840_),
    .A2(_03845_),
    .B1(_03863_),
    .C1(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__or4_1 _08334_ (.A(_03841_),
    .B(_03842_),
    .C(_03844_),
    .D(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__o21a_1 _08335_ (.A1(_01429_),
    .A2(_03837_),
    .B1(_03828_),
    .X(_03867_));
 sky130_fd_sc_hd__xnor2_1 _08336_ (.A(_01234_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__or4_1 _08337_ (.A(_03835_),
    .B(_03838_),
    .C(_03866_),
    .D(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__nand2_1 _08338_ (.A(_01296_),
    .B(\u_uart2wb.u_aut_det.ref1_cnt[17] ),
    .Y(_03870_));
 sky130_fd_sc_hd__a31o_1 _08339_ (.A1(_03826_),
    .A2(_03827_),
    .A3(_03833_),
    .B1(_01290_),
    .X(_03871_));
 sky130_fd_sc_hd__nand2_1 _08340_ (.A(_01343_),
    .B(_01340_),
    .Y(_03872_));
 sky130_fd_sc_hd__a21o_1 _08341_ (.A1(_03871_),
    .A2(_03872_),
    .B1(_01292_),
    .X(_03873_));
 sky130_fd_sc_hd__and3_1 _08342_ (.A(_01389_),
    .B(_03870_),
    .C(_03873_),
    .X(_03874_));
 sky130_fd_sc_hd__a21oi_1 _08343_ (.A1(_03870_),
    .A2(_03873_),
    .B1(_01389_),
    .Y(_03875_));
 sky130_fd_sc_hd__o311a_1 _08344_ (.A1(_03869_),
    .A2(_03874_),
    .A3(_03875_),
    .B1(_01433_),
    .C1(\u_uart2wb.u_aut_det.state[5] ),
    .X(_03876_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08345_ (.A(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__a21oi_1 _08346_ (.A1(_03809_),
    .A2(_03811_),
    .B1(_01189_),
    .Y(_03878_));
 sky130_fd_sc_hd__a211o_1 _08347_ (.A1(_01223_),
    .A2(_01222_),
    .B1(_01216_),
    .C1(_03878_),
    .X(_03879_));
 sky130_fd_sc_hd__and3b_1 _08348_ (.A_N(_03806_),
    .B(_03812_),
    .C(_03879_),
    .X(_03880_));
 sky130_fd_sc_hd__clkbuf_1 _08349_ (.A(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__inv_2 _08350_ (.A(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__a22o_1 _08351_ (.A1(\u_uart2wb.auto_baud_16x[0] ),
    .A2(_03805_),
    .B1(_03877_),
    .B2(_03882_),
    .X(_00827_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08352_ (.A(_03858_),
    .X(_03883_));
 sky130_fd_sc_hd__or2_1 _08353_ (.A(_03883_),
    .B(_03881_),
    .X(_03884_));
 sky130_fd_sc_hd__nand2_1 _08354_ (.A(_03883_),
    .B(_03881_),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_1 _08355_ (.A(_03884_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__a22o_1 _08356_ (.A1(\u_uart2wb.auto_baud_16x[1] ),
    .A2(_03805_),
    .B1(_03877_),
    .B2(_03886_),
    .X(_00828_));
 sky130_fd_sc_hd__xnor2_1 _08357_ (.A(_03855_),
    .B(_03884_),
    .Y(_03887_));
 sky130_fd_sc_hd__a22o_1 _08358_ (.A1(\u_uart2wb.auto_baud_16x[2] ),
    .A2(_03805_),
    .B1(_03877_),
    .B2(_03887_),
    .X(_00829_));
 sky130_fd_sc_hd__a2111o_1 _08359_ (.A1(_03849_),
    .A2(_03850_),
    .B1(_03855_),
    .C1(_03883_),
    .D1(_03880_),
    .X(_03888_));
 sky130_fd_sc_hd__o31ai_1 _08360_ (.A1(_03855_),
    .A2(_03883_),
    .A3(_03881_),
    .B1(_03851_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_1 _08361_ (.A(_03888_),
    .B(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__a22o_1 _08362_ (.A1(\u_uart2wb.auto_baud_16x[3] ),
    .A2(_03805_),
    .B1(_03877_),
    .B2(_03890_),
    .X(_00830_));
 sky130_fd_sc_hd__clkbuf_1 _08363_ (.A(_03804_),
    .X(_03891_));
 sky130_fd_sc_hd__clkbuf_1 _08364_ (.A(_03876_),
    .X(_03892_));
 sky130_fd_sc_hd__xnor2_1 _08365_ (.A(_03848_),
    .B(_03888_),
    .Y(_03893_));
 sky130_fd_sc_hd__a22o_1 _08366_ (.A1(\u_uart2wb.auto_baud_16x[4] ),
    .A2(_03891_),
    .B1(_03892_),
    .B2(_03893_),
    .X(_00831_));
 sky130_fd_sc_hd__a211o_1 _08367_ (.A1(_03840_),
    .A2(_03845_),
    .B1(_03888_),
    .C1(_03848_),
    .X(_03894_));
 sky130_fd_sc_hd__o211ai_1 _08368_ (.A1(_03848_),
    .A2(_03888_),
    .B1(_03845_),
    .C1(_03840_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand2_1 _08369_ (.A(_03894_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__a22o_1 _08370_ (.A1(\u_uart2wb.auto_baud_16x[5] ),
    .A2(_03891_),
    .B1(_03892_),
    .B2(_03896_),
    .X(_00832_));
 sky130_fd_sc_hd__or3_1 _08371_ (.A(_03841_),
    .B(_03842_),
    .C(_03894_),
    .X(_03897_));
 sky130_fd_sc_hd__o21ai_1 _08372_ (.A1(_03841_),
    .A2(_03842_),
    .B1(_03894_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand2_1 _08373_ (.A(_03897_),
    .B(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__a22o_1 _08374_ (.A1(\u_uart2wb.auto_baud_16x[6] ),
    .A2(_03891_),
    .B1(_03892_),
    .B2(_03899_),
    .X(_00833_));
 sky130_fd_sc_hd__nor2_1 _08375_ (.A(_03864_),
    .B(_03897_),
    .Y(_03900_));
 sky130_fd_sc_hd__nand2_1 _08376_ (.A(_03864_),
    .B(_03897_),
    .Y(_03901_));
 sky130_fd_sc_hd__or2b_1 _08377_ (.A(_03900_),
    .B_N(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__a22o_1 _08378_ (.A1(\u_uart2wb.auto_baud_16x[7] ),
    .A2(_03891_),
    .B1(_03892_),
    .B2(_03902_),
    .X(_00834_));
 sky130_fd_sc_hd__clkbuf_1 _08379_ (.A(_03804_),
    .X(_03903_));
 sky130_fd_sc_hd__clkbuf_1 _08380_ (.A(_03876_),
    .X(_03904_));
 sky130_fd_sc_hd__xnor2_1 _08381_ (.A(_01411_),
    .B(_03843_),
    .Y(_03905_));
 sky130_fd_sc_hd__xnor2_1 _08382_ (.A(_03905_),
    .B(_03900_),
    .Y(_03906_));
 sky130_fd_sc_hd__a22o_1 _08383_ (.A1(\u_uart2wb.auto_baud_16x[8] ),
    .A2(_03903_),
    .B1(_03904_),
    .B2(_03906_),
    .X(_00835_));
 sky130_fd_sc_hd__a21bo_1 _08384_ (.A1(_03905_),
    .A2(_03900_),
    .B1_N(_03838_),
    .X(_03907_));
 sky130_fd_sc_hd__or4_1 _08385_ (.A(_03838_),
    .B(_03844_),
    .C(_03864_),
    .D(_03897_),
    .X(_03908_));
 sky130_fd_sc_hd__nand2_1 _08386_ (.A(_03907_),
    .B(_03908_),
    .Y(_03909_));
 sky130_fd_sc_hd__a22o_1 _08387_ (.A1(\u_uart2wb.auto_baud_16x[9] ),
    .A2(_03903_),
    .B1(_03904_),
    .B2(_03909_),
    .X(_00836_));
 sky130_fd_sc_hd__nor2_1 _08388_ (.A(_03868_),
    .B(_03908_),
    .Y(_03910_));
 sky130_fd_sc_hd__and2_1 _08389_ (.A(_03868_),
    .B(_03908_),
    .X(_03911_));
 sky130_fd_sc_hd__or2_1 _08390_ (.A(_03910_),
    .B(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__a22o_1 _08391_ (.A1(\u_uart2wb.auto_baud_16x[10] ),
    .A2(_03903_),
    .B1(_03904_),
    .B2(_03912_),
    .X(_00837_));
 sky130_fd_sc_hd__xor2_1 _08392_ (.A(_03835_),
    .B(_03910_),
    .X(_03913_));
 sky130_fd_sc_hd__a22o_1 _08393_ (.A1(\u_uart2wb.auto_baud_16x[11] ),
    .A2(_03903_),
    .B1(_03904_),
    .B2(_03913_),
    .X(_00838_));
 sky130_fd_sc_hd__inv_2 _08394_ (.A(\u_uart2wb.u_core.u_txfsm.cnt[0] ),
    .Y(_03914_));
 sky130_fd_sc_hd__o21ba_1 _08395_ (.A1(\u_uart2wb.u_core.u_txfsm.cnt[0] ),
    .A2(\u_uart2wb.u_core.u_txfsm.txdata[0] ),
    .B1_N(\u_uart2wb.u_core.u_txfsm.cnt[1] ),
    .X(_03915_));
 sky130_fd_sc_hd__o21a_1 _08396_ (.A1(_03914_),
    .A2(\u_uart2wb.u_core.u_txfsm.txdata[1] ),
    .B1(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__a31o_1 _08397_ (.A1(\u_uart2wb.u_core.u_txfsm.cnt[1] ),
    .A2(_01140_),
    .A3(\u_uart2wb.u_core.u_txfsm.txdata[3] ),
    .B1(\u_uart2wb.u_core.u_txfsm.cnt[2] ),
    .X(_03917_));
 sky130_fd_sc_hd__a311o_1 _08398_ (.A1(_01139_),
    .A2(_03914_),
    .A3(\u_uart2wb.u_core.u_txfsm.txdata[2] ),
    .B1(_03916_),
    .C1(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__mux2_1 _08399_ (.A0(\u_uart2wb.u_core.u_txfsm.txdata[4] ),
    .A1(\u_uart2wb.u_core.u_txfsm.txdata[5] ),
    .S(\u_uart2wb.u_core.u_txfsm.cnt[0] ),
    .X(_03919_));
 sky130_fd_sc_hd__inv_2 _08400_ (.A(_03919_),
    .Y(_03920_));
 sky130_fd_sc_hd__o21ai_1 _08401_ (.A1(\u_uart2wb.u_core.u_txfsm.cnt[1] ),
    .A2(_03920_),
    .B1(\u_uart2wb.u_core.u_txfsm.cnt[2] ),
    .Y(_03921_));
 sky130_fd_sc_hd__a31o_1 _08402_ (.A1(_01139_),
    .A2(_03914_),
    .A3(\u_uart2wb.u_core.u_txfsm.txdata[6] ),
    .B1(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__or3b_1 _08403_ (.A(_01156_),
    .B(la_data_in[16]),
    .C_N(la_data_in[17]),
    .X(_03923_));
 sky130_fd_sc_hd__xor2_1 _08404_ (.A(\u_uart2wb.u_core.u_txfsm.txdata[3] ),
    .B(\u_uart2wb.u_core.u_txfsm.txdata[2] ),
    .X(_03924_));
 sky130_fd_sc_hd__xnor2_1 _08405_ (.A(\u_uart2wb.u_core.u_txfsm.txdata[5] ),
    .B(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__xnor2_1 _08406_ (.A(\u_uart2wb.u_core.u_txfsm.txdata[1] ),
    .B(\u_uart2wb.u_core.u_txfsm.txdata[0] ),
    .Y(_03926_));
 sky130_fd_sc_hd__xnor2_1 _08407_ (.A(\u_uart2wb.u_core.u_txfsm.txdata[4] ),
    .B(\u_uart2wb.u_core.u_txfsm.txdata[6] ),
    .Y(_03927_));
 sky130_fd_sc_hd__xnor2_1 _08408_ (.A(_03926_),
    .B(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__xnor2_1 _08409_ (.A(_03925_),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__xnor2_1 _08410_ (.A(_03923_),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__a32o_1 _08411_ (.A1(\u_uart2wb.u_core.u_txfsm.txstate[3] ),
    .A2(_03918_),
    .A3(_03922_),
    .B1(_03930_),
    .B2(\u_uart2wb.u_core.u_txfsm.txstate[2] ),
    .X(_03931_));
 sky130_fd_sc_hd__or3_1 _08412_ (.A(\u_uart2wb.u_core.u_txfsm.txstate[4] ),
    .B(\u_uart2wb.u_core.u_txfsm.txstate[1] ),
    .C(_03931_),
    .X(_03932_));
 sky130_fd_sc_hd__nor2_1 _08413_ (.A(_01138_),
    .B(_01185_),
    .Y(_03933_));
 sky130_fd_sc_hd__o41a_1 _08414_ (.A1(\u_uart2wb.u_core.u_txfsm.txstate[2] ),
    .A2(\u_uart2wb.u_core.u_txfsm.txstate[3] ),
    .A3(\u_uart2wb.u_core.u_txfsm.txstate[0] ),
    .A4(_01186_),
    .B1(_03933_),
    .X(_03934_));
 sky130_fd_sc_hd__mux2_1 _08415_ (.A0(net105),
    .A1(_03932_),
    .S(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__clkbuf_1 _08416_ (.A(_03935_),
    .X(_00839_));
 sky130_fd_sc_hd__a31o_1 _08417_ (.A1(\u_uart2wb.tx_data_avail ),
    .A2(_01184_),
    .A3(_01159_),
    .B1(\u_uart2wb.tx_rd ),
    .X(_03936_));
 sky130_fd_sc_hd__o211a_1 _08418_ (.A1(_01151_),
    .A2(_01185_),
    .B1(_03936_),
    .C1(_01135_),
    .X(_00840_));
 sky130_fd_sc_hd__clkbuf_1 _08419_ (.A(\u_uart2wb.u_core.u_rxfsm.rxstate[0] ),
    .X(_03937_));
 sky130_fd_sc_hd__clkbuf_1 _08420_ (.A(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__clkbuf_1 _08421_ (.A(\u_uart2wb.u_core.u_rxfsm.rxstate[1] ),
    .X(_03939_));
 sky130_fd_sc_hd__or2_1 _08422_ (.A(_03939_),
    .B(\u_uart2wb.u_core.u_rxfsm.rxstate[2] ),
    .X(_03940_));
 sky130_fd_sc_hd__nor2_1 _08423_ (.A(_03937_),
    .B(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__nor2_1 _08424_ (.A(_03937_),
    .B(_03939_),
    .Y(_03942_));
 sky130_fd_sc_hd__clkbuf_1 _08425_ (.A(\u_uart2wb.u_core.u_rxfsm.rxstate[2] ),
    .X(_03943_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08426_ (.A(\u_uart2wb.u_core.si_ss ),
    .X(_03944_));
 sky130_fd_sc_hd__and4b_1 _08427_ (.A_N(_01163_),
    .B(_03942_),
    .C(_03943_),
    .D(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__or3b_1 _08428_ (.A(\u_uart2wb.u_core.u_rxfsm.rxstate[0] ),
    .B(\u_uart2wb.u_core.u_rxfsm.rxstate[2] ),
    .C_N(\u_uart2wb.u_core.u_rxfsm.rxstate[1] ),
    .X(_03946_));
 sky130_fd_sc_hd__nor2_1 _08429_ (.A(_01149_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__or3_1 _08430_ (.A(_03941_),
    .B(_03945_),
    .C(_03947_),
    .X(_03948_));
 sky130_fd_sc_hd__xor2_1 _08431_ (.A(\u_uart2wb.u_core.u_rxfsm.offset[3] ),
    .B(\u_uart2wb.u_core.u_rxfsm.rxpos[3] ),
    .X(_03949_));
 sky130_fd_sc_hd__xor2_1 _08432_ (.A(\u_uart2wb.u_core.u_rxfsm.offset[0] ),
    .B(\u_uart2wb.u_core.u_rxfsm.rxpos[0] ),
    .X(_03950_));
 sky130_fd_sc_hd__xor2_1 _08433_ (.A(\u_uart2wb.u_core.u_rxfsm.rxpos[1] ),
    .B(\u_uart2wb.u_core.u_rxfsm.offset[1] ),
    .X(_03951_));
 sky130_fd_sc_hd__xor2_1 _08434_ (.A(\u_uart2wb.u_core.u_rxfsm.rxpos[2] ),
    .B(\u_uart2wb.u_core.u_rxfsm.offset[2] ),
    .X(_03952_));
 sky130_fd_sc_hd__or4_2 _08435_ (.A(_03949_),
    .B(_03950_),
    .C(_03951_),
    .D(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__inv_2 _08436_ (.A(\u_uart2wb.u_core.u_rxfsm.cnt[2] ),
    .Y(_03954_));
 sky130_fd_sc_hd__nand2_1 _08437_ (.A(\u_uart2wb.u_core.u_rxfsm.cnt[1] ),
    .B(\u_uart2wb.u_core.u_rxfsm.cnt[0] ),
    .Y(_03955_));
 sky130_fd_sc_hd__or2_1 _08438_ (.A(_03954_),
    .B(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__clkbuf_1 _08439_ (.A(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__nor2_1 _08440_ (.A(_03953_),
    .B(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__clkbuf_1 _08441_ (.A(_03939_),
    .X(_03959_));
 sky130_fd_sc_hd__inv_2 _08442_ (.A(_03943_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand4_1 _08443_ (.A(_03937_),
    .B(_03959_),
    .C(_03960_),
    .D(_03953_),
    .Y(_03961_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(_03943_),
    .B(_03953_),
    .Y(_03962_));
 sky130_fd_sc_hd__inv_2 _08445_ (.A(la_data_in[2]),
    .Y(_03963_));
 sky130_fd_sc_hd__inv_2 _08446_ (.A(\u_uart2wb.auto_rx_enb ),
    .Y(_03964_));
 sky130_fd_sc_hd__a221o_1 _08447_ (.A1(_03963_),
    .A2(_01146_),
    .B1(_01435_),
    .B2(_03964_),
    .C1(\u_uart2wb.u_core.si_ss ),
    .X(_03965_));
 sky130_fd_sc_hd__nand2_1 _08448_ (.A(_03965_),
    .B(_03941_),
    .Y(_03966_));
 sky130_fd_sc_hd__or3b_1 _08449_ (.A(\u_uart2wb.u_core.u_rxfsm.rxstate[1] ),
    .B(\u_uart2wb.u_core.u_rxfsm.rxstate[2] ),
    .C_N(\u_uart2wb.u_core.u_rxfsm.rxstate[0] ),
    .X(_03967_));
 sky130_fd_sc_hd__a21oi_1 _08450_ (.A1(\u_uart2wb.u_core.si_ss ),
    .A2(_03956_),
    .B1(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__o21ai_1 _08451_ (.A1(\u_uart2wb.u_core.si_ss ),
    .A2(_03956_),
    .B1(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__o211a_1 _08452_ (.A1(_03939_),
    .A2(_03962_),
    .B1(_03966_),
    .C1(_03969_),
    .X(_03970_));
 sky130_fd_sc_hd__o211a_1 _08453_ (.A1(_03946_),
    .A2(_03958_),
    .B1(_03961_),
    .C1(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__mux2_1 _08454_ (.A0(_03938_),
    .A1(_03948_),
    .S(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__clkbuf_1 _08455_ (.A(_03972_),
    .X(_00841_));
 sky130_fd_sc_hd__inv_2 _08456_ (.A(_03971_),
    .Y(_03973_));
 sky130_fd_sc_hd__o31a_1 _08457_ (.A1(_03968_),
    .A2(_03973_),
    .A3(_03947_),
    .B1(_03970_),
    .X(_00842_));
 sky130_fd_sc_hd__or2_1 _08458_ (.A(_03938_),
    .B(_01149_),
    .X(_03974_));
 sky130_fd_sc_hd__a31o_1 _08459_ (.A1(_03959_),
    .A2(_03960_),
    .A3(_03974_),
    .B1(_03945_),
    .X(_03975_));
 sky130_fd_sc_hd__a2bb2o_1 _08460_ (.A1_N(_03959_),
    .A2_N(_03962_),
    .B1(_03971_),
    .B2(_03975_),
    .X(_00843_));
 sky130_fd_sc_hd__or3_2 _08461_ (.A(_03938_),
    .B(_03965_),
    .C(_03940_),
    .X(_03976_));
 sky130_fd_sc_hd__mux2_1 _08462_ (.A0(_01108_),
    .A1(\u_uart2wb.u_core.u_rxfsm.rxpos[0] ),
    .S(_03976_),
    .X(_03977_));
 sky130_fd_sc_hd__clkbuf_1 _08463_ (.A(_03977_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _08464_ (.A0(_01810_),
    .A1(\u_uart2wb.u_core.u_rxfsm.rxpos[1] ),
    .S(_03976_),
    .X(_03978_));
 sky130_fd_sc_hd__clkbuf_1 _08465_ (.A(_03978_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _08466_ (.A0(\u_uart2wb.u_core.u_rxfsm.offset[2] ),
    .A1(\u_uart2wb.u_core.u_rxfsm.rxpos[2] ),
    .S(_03976_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_1 _08467_ (.A(_03979_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _08468_ (.A0(_01813_),
    .A1(\u_uart2wb.u_core.u_rxfsm.rxpos[3] ),
    .S(_03976_),
    .X(_03980_));
 sky130_fd_sc_hd__clkbuf_1 _08469_ (.A(_03980_),
    .X(_00847_));
 sky130_fd_sc_hd__nor2_1 _08470_ (.A(_03959_),
    .B(_03945_),
    .Y(_03981_));
 sky130_fd_sc_hd__nand3b_1 _08471_ (.A_N(_03938_),
    .B(_03962_),
    .C(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__clkbuf_1 _08472_ (.A(\u_uart2wb.rx_wr ),
    .X(_03983_));
 sky130_fd_sc_hd__clkbuf_2 _08473_ (.A(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__a32o_1 _08474_ (.A1(_03943_),
    .A2(_03962_),
    .A3(_03981_),
    .B1(_03982_),
    .B2(_03984_),
    .X(_00848_));
 sky130_fd_sc_hd__clkbuf_1 _08475_ (.A(\u_uart2wb.u_core.u_rxfsm.cnt[0] ),
    .X(_03985_));
 sky130_fd_sc_hd__clkbuf_1 _08476_ (.A(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__nor2_1 _08477_ (.A(_03986_),
    .B(_03942_),
    .Y(_03987_));
 sky130_fd_sc_hd__inv_2 _08478_ (.A(_03967_),
    .Y(_03988_));
 sky130_fd_sc_hd__or2_1 _08479_ (.A(_03953_),
    .B(_03946_),
    .X(_03989_));
 sky130_fd_sc_hd__a21bo_1 _08480_ (.A1(_03940_),
    .A2(_03989_),
    .B1_N(_03966_),
    .X(_03990_));
 sky130_fd_sc_hd__a31o_1 _08481_ (.A1(_03944_),
    .A2(_03957_),
    .A3(_03988_),
    .B1(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__mux2_1 _08482_ (.A0(_03987_),
    .A1(_03986_),
    .S(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__clkbuf_1 _08483_ (.A(_03992_),
    .X(_00849_));
 sky130_fd_sc_hd__or2_1 _08484_ (.A(\u_uart2wb.u_core.u_rxfsm.cnt[1] ),
    .B(_03985_),
    .X(_03993_));
 sky130_fd_sc_hd__nand2_1 _08485_ (.A(_03946_),
    .B(_03967_),
    .Y(_03994_));
 sky130_fd_sc_hd__and3_1 _08486_ (.A(_03955_),
    .B(_03993_),
    .C(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__clkbuf_1 _08487_ (.A(\u_uart2wb.u_core.u_rxfsm.cnt[1] ),
    .X(_03996_));
 sky130_fd_sc_hd__mux2_1 _08488_ (.A0(_03995_),
    .A1(_03996_),
    .S(_03991_),
    .X(_03997_));
 sky130_fd_sc_hd__clkbuf_1 _08489_ (.A(_03997_),
    .X(_00850_));
 sky130_fd_sc_hd__or2_1 _08490_ (.A(_03955_),
    .B(_03991_),
    .X(_03998_));
 sky130_fd_sc_hd__a21oi_1 _08491_ (.A1(_03957_),
    .A2(_03994_),
    .B1(_03991_),
    .Y(_03999_));
 sky130_fd_sc_hd__a21oi_1 _08492_ (.A1(_03954_),
    .A2(_03998_),
    .B1(_03999_),
    .Y(_00851_));
 sky130_fd_sc_hd__clkbuf_1 _08493_ (.A(_03944_),
    .X(_04000_));
 sky130_fd_sc_hd__clkbuf_1 _08494_ (.A(\u_uart2wb.rx_data[0] ),
    .X(_04001_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08495_ (.A(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__or2_1 _08496_ (.A(\u_uart2wb.u_core.u_rxfsm.cnt[2] ),
    .B(_03989_),
    .X(_04003_));
 sky130_fd_sc_hd__or2_1 _08497_ (.A(_03993_),
    .B(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__mux2_1 _08498_ (.A0(_04000_),
    .A1(_04002_),
    .S(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__clkbuf_1 _08499_ (.A(_04005_),
    .X(_00852_));
 sky130_fd_sc_hd__clkbuf_1 _08500_ (.A(\u_uart2wb.rx_data[1] ),
    .X(_04006_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08501_ (.A(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__or3b_1 _08502_ (.A(_04003_),
    .B(_03996_),
    .C_N(_03986_),
    .X(_04008_));
 sky130_fd_sc_hd__mux2_1 _08503_ (.A0(_04000_),
    .A1(_04007_),
    .S(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__clkbuf_1 _08504_ (.A(_04009_),
    .X(_00853_));
 sky130_fd_sc_hd__clkbuf_1 _08505_ (.A(\u_uart2wb.rx_data[2] ),
    .X(_04010_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08506_ (.A(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__or3b_1 _08507_ (.A(_03985_),
    .B(_04003_),
    .C_N(_03996_),
    .X(_04012_));
 sky130_fd_sc_hd__mux2_1 _08508_ (.A0(_04000_),
    .A1(_04011_),
    .S(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__clkbuf_1 _08509_ (.A(_04013_),
    .X(_00854_));
 sky130_fd_sc_hd__clkbuf_1 _08510_ (.A(\u_uart2wb.rx_data[3] ),
    .X(_04014_));
 sky130_fd_sc_hd__clkbuf_1 _08511_ (.A(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__clkbuf_1 _08512_ (.A(_03944_),
    .X(_04016_));
 sky130_fd_sc_hd__nor2_1 _08513_ (.A(_03955_),
    .B(_04003_),
    .Y(_04017_));
 sky130_fd_sc_hd__mux2_1 _08514_ (.A0(_04015_),
    .A1(_04016_),
    .S(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__clkbuf_1 _08515_ (.A(_04018_),
    .X(_00855_));
 sky130_fd_sc_hd__clkbuf_1 _08516_ (.A(\u_uart2wb.rx_data[4] ),
    .X(_04019_));
 sky130_fd_sc_hd__or2_1 _08517_ (.A(_03954_),
    .B(_03989_),
    .X(_04020_));
 sky130_fd_sc_hd__or2_1 _08518_ (.A(_03993_),
    .B(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__mux2_1 _08519_ (.A0(_04000_),
    .A1(_04019_),
    .S(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__clkbuf_1 _08520_ (.A(_04022_),
    .X(_00856_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08521_ (.A(\u_uart2wb.rx_data[5] ),
    .X(_04023_));
 sky130_fd_sc_hd__or3b_1 _08522_ (.A(_04020_),
    .B(\u_uart2wb.u_core.u_rxfsm.cnt[1] ),
    .C_N(_03986_),
    .X(_04024_));
 sky130_fd_sc_hd__mux2_1 _08523_ (.A0(_04016_),
    .A1(_04023_),
    .S(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__clkbuf_1 _08524_ (.A(_04025_),
    .X(_00857_));
 sky130_fd_sc_hd__clkbuf_1 _08525_ (.A(\u_uart2wb.rx_data[6] ),
    .X(_04026_));
 sky130_fd_sc_hd__or3b_1 _08526_ (.A(_03985_),
    .B(_04020_),
    .C_N(_03996_),
    .X(_04027_));
 sky130_fd_sc_hd__mux2_1 _08527_ (.A0(_04016_),
    .A1(_04026_),
    .S(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__clkbuf_1 _08528_ (.A(_04028_),
    .X(_00858_));
 sky130_fd_sc_hd__clkbuf_1 _08529_ (.A(\u_uart2wb.rx_data[7] ),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_1 _08530_ (.A(_03957_),
    .B(_03989_),
    .Y(_04030_));
 sky130_fd_sc_hd__mux2_1 _08531_ (.A0(_04029_),
    .A1(_04016_),
    .S(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__clkbuf_1 _08532_ (.A(_04031_),
    .X(_00859_));
 sky130_fd_sc_hd__clkbuf_1 _08533_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[0] ),
    .X(_04032_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08534_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[11] ),
    .X(_04033_));
 sky130_fd_sc_hd__nor3_2 _08535_ (.A(_04033_),
    .B(\u_uart2wb.u_core.u_clk_ctl.low_count[10] ),
    .C(_01822_),
    .Y(_04034_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08536_ (.A(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__a22o_1 _08537_ (.A1(la_data_in[5]),
    .A2(_01145_),
    .B1(_01434_),
    .B2(\u_uart2wb.auto_baud_16x[1] ),
    .X(_04036_));
 sky130_fd_sc_hd__clkbuf_1 _08538_ (.A(_04036_),
    .X(_04037_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08539_ (.A(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__a21oi_1 _08540_ (.A1(_04035_),
    .A2(_04038_),
    .B1(_04032_),
    .Y(_04039_));
 sky130_fd_sc_hd__mux2_1 _08541_ (.A0(_04032_),
    .A1(_04039_),
    .S(_01832_),
    .X(_04040_));
 sky130_fd_sc_hd__clkbuf_1 _08542_ (.A(_04040_),
    .X(_00860_));
 sky130_fd_sc_hd__xnor2_1 _08543_ (.A(_04032_),
    .B(\u_uart2wb.u_core.u_clk_ctl.low_count[1] ),
    .Y(_04041_));
 sky130_fd_sc_hd__inv_2 _08544_ (.A(strap_uartm[1]),
    .Y(_04042_));
 sky130_fd_sc_hd__clkbuf_1 _08545_ (.A(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__or2b_1 _08546_ (.A(la_data_in[6]),
    .B_N(_01144_),
    .X(_04044_));
 sky130_fd_sc_hd__a22o_1 _08547_ (.A1(_04043_),
    .A2(\u_uart2wb.auto_baud_16x[2] ),
    .B1(_04044_),
    .B2(_01153_),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_1 _08548_ (.A(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__nand2_1 _08549_ (.A(_04038_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__o21a_1 _08550_ (.A1(_04037_),
    .A2(_04046_),
    .B1(_04034_),
    .X(_04048_));
 sky130_fd_sc_hd__or2_1 _08551_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[11] ),
    .B(_01831_),
    .X(_04049_));
 sky130_fd_sc_hd__clkbuf_1 _08552_ (.A(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__a221o_1 _08553_ (.A1(_01825_),
    .A2(_04041_),
    .B1(_04047_),
    .B2(_04048_),
    .C1(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__o21a_1 _08554_ (.A1(\u_uart2wb.u_core.u_clk_ctl.low_count[1] ),
    .A2(_01834_),
    .B1(_04051_),
    .X(_00861_));
 sky130_fd_sc_hd__inv_2 _08555_ (.A(strap_uartm[0]),
    .Y(_04052_));
 sky130_fd_sc_hd__or2b_1 _08556_ (.A(la_data_in[7]),
    .B_N(_01153_),
    .X(_04053_));
 sky130_fd_sc_hd__a22o_1 _08557_ (.A1(_04052_),
    .A2(\u_uart2wb.auto_baud_16x[3] ),
    .B1(_04053_),
    .B2(_01155_),
    .X(_04054_));
 sky130_fd_sc_hd__and3_1 _08558_ (.A(_04036_),
    .B(_04045_),
    .C(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__a21oi_1 _08559_ (.A1(_04037_),
    .A2(_04046_),
    .B1(_04054_),
    .Y(_04056_));
 sky130_fd_sc_hd__o21ai_1 _08560_ (.A1(_04032_),
    .A2(\u_uart2wb.u_core.u_clk_ctl.low_count[1] ),
    .B1(\u_uart2wb.u_core.u_clk_ctl.low_count[2] ),
    .Y(_04057_));
 sky130_fd_sc_hd__a21o_1 _08561_ (.A1(_01816_),
    .A2(_04057_),
    .B1(_04034_),
    .X(_04058_));
 sky130_fd_sc_hd__o311a_1 _08562_ (.A1(_01824_),
    .A2(_04055_),
    .A3(_04056_),
    .B1(_04058_),
    .C1(_01833_),
    .X(_04059_));
 sky130_fd_sc_hd__o21ba_1 _08563_ (.A1(\u_uart2wb.u_core.u_clk_ctl.low_count[2] ),
    .A2(_01834_),
    .B1_N(_04059_),
    .X(_00862_));
 sky130_fd_sc_hd__clkbuf_1 _08564_ (.A(_04049_),
    .X(_04060_));
 sky130_fd_sc_hd__nor2_1 _08565_ (.A(_04060_),
    .B(_04034_),
    .Y(_04061_));
 sky130_fd_sc_hd__nand2_1 _08566_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[3] ),
    .B(_01816_),
    .Y(_04062_));
 sky130_fd_sc_hd__and3_1 _08567_ (.A(_01817_),
    .B(_04061_),
    .C(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__nor2_1 _08568_ (.A(_04049_),
    .B(_01823_),
    .Y(_04064_));
 sky130_fd_sc_hd__or2b_1 _08569_ (.A(la_data_in[8]),
    .B_N(strap_uartm[0]),
    .X(_04065_));
 sky130_fd_sc_hd__a22o_1 _08570_ (.A1(_04052_),
    .A2(\u_uart2wb.auto_baud_16x[4] ),
    .B1(_04065_),
    .B2(_01155_),
    .X(_04066_));
 sky130_fd_sc_hd__and4_1 _08571_ (.A(_04036_),
    .B(_04045_),
    .C(_04054_),
    .D(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__nor2_1 _08572_ (.A(_04055_),
    .B(_04066_),
    .Y(_04068_));
 sky130_fd_sc_hd__or2_1 _08573_ (.A(_04067_),
    .B(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__a2bb2o_1 _08574_ (.A1_N(\u_uart2wb.u_core.u_clk_ctl.low_count[3] ),
    .A2_N(_01833_),
    .B1(_04064_),
    .B2(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__nor2_1 _08575_ (.A(_04063_),
    .B(_04070_),
    .Y(_00863_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08576_ (.A(_04050_),
    .X(_04071_));
 sky130_fd_sc_hd__nand2_1 _08577_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[4] ),
    .B(_01817_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand2_1 _08578_ (.A(_01818_),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__a22o_1 _08579_ (.A1(la_data_in[9]),
    .A2(_01145_),
    .B1(_01434_),
    .B2(\u_uart2wb.auto_baud_16x[5] ),
    .X(_04074_));
 sky130_fd_sc_hd__nand2_1 _08580_ (.A(_04067_),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__or2_1 _08581_ (.A(_04067_),
    .B(_04074_),
    .X(_04076_));
 sky130_fd_sc_hd__and2_1 _08582_ (.A(_04075_),
    .B(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__o21a_1 _08583_ (.A1(_01825_),
    .A2(_04077_),
    .B1(_01833_),
    .X(_04078_));
 sky130_fd_sc_hd__a22o_1 _08584_ (.A1(\u_uart2wb.u_core.u_clk_ctl.low_count[4] ),
    .A2(_04071_),
    .B1(_04073_),
    .B2(_04078_),
    .X(_00864_));
 sky130_fd_sc_hd__inv_2 _08585_ (.A(_01819_),
    .Y(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _08586_ (.A(_04064_),
    .X(_04080_));
 sky130_fd_sc_hd__or2_1 _08587_ (.A(_04042_),
    .B(la_data_in[10]),
    .X(_04081_));
 sky130_fd_sc_hd__a22o_1 _08588_ (.A1(_04043_),
    .A2(\u_uart2wb.auto_baud_16x[6] ),
    .B1(_04081_),
    .B2(_01154_),
    .X(_04082_));
 sky130_fd_sc_hd__inv_2 _08589_ (.A(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__nor2_1 _08590_ (.A(_04075_),
    .B(_04083_),
    .Y(_04084_));
 sky130_fd_sc_hd__and2_1 _08591_ (.A(_04075_),
    .B(_04083_),
    .X(_04085_));
 sky130_fd_sc_hd__nor2_1 _08592_ (.A(_04084_),
    .B(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__o21a_1 _08593_ (.A1(_04060_),
    .A2(_01818_),
    .B1(\u_uart2wb.u_core.u_clk_ctl.low_count[5] ),
    .X(_04087_));
 sky130_fd_sc_hd__a221o_1 _08594_ (.A1(_04079_),
    .A2(_04061_),
    .B1(_04080_),
    .B2(_04086_),
    .C1(_04087_),
    .X(_00865_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08595_ (.A(_04060_),
    .X(_04088_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08596_ (.A(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__a22o_1 _08597_ (.A1(la_data_in[11]),
    .A2(_01145_),
    .B1(_01435_),
    .B2(\u_uart2wb.auto_baud_16x[7] ),
    .X(_04090_));
 sky130_fd_sc_hd__nand2_1 _08598_ (.A(_04084_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__or2_1 _08599_ (.A(_04084_),
    .B(_04090_),
    .X(_04092_));
 sky130_fd_sc_hd__nand2_1 _08600_ (.A(_04091_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__nand2_1 _08601_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[6] ),
    .B(_01819_),
    .Y(_04094_));
 sky130_fd_sc_hd__clkbuf_1 _08602_ (.A(_01820_),
    .X(_04095_));
 sky130_fd_sc_hd__a221o_1 _08603_ (.A1(_04035_),
    .A2(_04093_),
    .B1(_04094_),
    .B2(_04095_),
    .C1(_04050_),
    .X(_04096_));
 sky130_fd_sc_hd__a21bo_1 _08604_ (.A1(\u_uart2wb.u_core.u_clk_ctl.low_count[6] ),
    .A2(_04089_),
    .B1_N(_04096_),
    .X(_00866_));
 sky130_fd_sc_hd__nor2_1 _08605_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[7] ),
    .B(_04095_),
    .Y(_04097_));
 sky130_fd_sc_hd__a21o_1 _08606_ (.A1(_04043_),
    .A2(\u_uart2wb.auto_baud_16x[8] ),
    .B1(_01154_),
    .X(_04098_));
 sky130_fd_sc_hd__o21ai_1 _08607_ (.A1(_04043_),
    .A2(la_data_in[12]),
    .B1(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__nor2_1 _08608_ (.A(_04091_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _08609_ (.A(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__and2_1 _08610_ (.A(_04091_),
    .B(_04099_),
    .X(_04102_));
 sky130_fd_sc_hd__nor2_1 _08611_ (.A(_04101_),
    .B(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__o21a_1 _08612_ (.A1(_04060_),
    .A2(_04095_),
    .B1(\u_uart2wb.u_core.u_clk_ctl.low_count[7] ),
    .X(_04104_));
 sky130_fd_sc_hd__a221o_1 _08613_ (.A1(_04097_),
    .A2(_04061_),
    .B1(_04080_),
    .B2(_04103_),
    .C1(_04104_),
    .X(_00867_));
 sky130_fd_sc_hd__inv_2 _08614_ (.A(_01821_),
    .Y(_04105_));
 sky130_fd_sc_hd__clkbuf_1 _08615_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[10] ),
    .X(_04106_));
 sky130_fd_sc_hd__a22o_1 _08616_ (.A1(la_data_in[13]),
    .A2(_01146_),
    .B1(_01435_),
    .B2(\u_uart2wb.auto_baud_16x[9] ),
    .X(_04107_));
 sky130_fd_sc_hd__and2_1 _08617_ (.A(_04100_),
    .B(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__nor2_1 _08618_ (.A(_04101_),
    .B(_04107_),
    .Y(_04109_));
 sky130_fd_sc_hd__nor2_1 _08619_ (.A(_04108_),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__or4_1 _08620_ (.A(\u_uart2wb.u_core.u_clk_ctl.low_count[9] ),
    .B(_04033_),
    .C(_04106_),
    .D(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__o31a_1 _08621_ (.A1(\u_uart2wb.u_core.u_clk_ctl.low_count[7] ),
    .A2(_04050_),
    .A3(_04095_),
    .B1(\u_uart2wb.u_core.u_clk_ctl.low_count[8] ),
    .X(_04112_));
 sky130_fd_sc_hd__a31o_1 _08622_ (.A1(_01834_),
    .A2(_04105_),
    .A3(_04111_),
    .B1(_04112_),
    .X(_00868_));
 sky130_fd_sc_hd__or2_1 _08623_ (.A(_04049_),
    .B(_01822_),
    .X(_04113_));
 sky130_fd_sc_hd__o21ai_1 _08624_ (.A1(_04088_),
    .A2(_01821_),
    .B1(\u_uart2wb.u_core.u_clk_ctl.low_count[9] ),
    .Y(_04114_));
 sky130_fd_sc_hd__a22o_1 _08625_ (.A1(la_data_in[14]),
    .A2(_01146_),
    .B1(_01436_),
    .B2(\u_uart2wb.auto_baud_16x[10] ),
    .X(_04115_));
 sky130_fd_sc_hd__nand2_1 _08626_ (.A(_04108_),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _08627_ (.A(_04108_),
    .X(_04117_));
 sky130_fd_sc_hd__clkbuf_1 _08628_ (.A(_04115_),
    .X(_04118_));
 sky130_fd_sc_hd__or2_1 _08629_ (.A(_04117_),
    .B(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__nand2_1 _08630_ (.A(_04116_),
    .B(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08631_ (.A(_04080_),
    .X(_04121_));
 sky130_fd_sc_hd__a22oi_1 _08632_ (.A1(_04113_),
    .A2(_04114_),
    .B1(_04120_),
    .B2(_04121_),
    .Y(_00869_));
 sky130_fd_sc_hd__inv_2 _08633_ (.A(_04033_),
    .Y(_04122_));
 sky130_fd_sc_hd__a22o_1 _08634_ (.A1(la_data_in[15]),
    .A2(_01147_),
    .B1(_01436_),
    .B2(\u_uart2wb.auto_baud_16x[11] ),
    .X(_04123_));
 sky130_fd_sc_hd__xor2_1 _08635_ (.A(_04116_),
    .B(_04123_),
    .X(_04124_));
 sky130_fd_sc_hd__a211o_1 _08636_ (.A1(_04122_),
    .A2(_04124_),
    .B1(_04113_),
    .C1(_04106_),
    .X(_04125_));
 sky130_fd_sc_hd__a21bo_1 _08637_ (.A1(_04106_),
    .A2(_04113_),
    .B1_N(_04125_),
    .X(_00870_));
 sky130_fd_sc_hd__and3_1 _08638_ (.A(_04108_),
    .B(_04115_),
    .C(_04123_),
    .X(_04126_));
 sky130_fd_sc_hd__o21a_1 _08639_ (.A1(_04106_),
    .A2(_04113_),
    .B1(_04033_),
    .X(_04127_));
 sky130_fd_sc_hd__a21o_1 _08640_ (.A1(_04121_),
    .A2(_04126_),
    .B1(_04127_),
    .X(_00871_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08641_ (.A(_01832_),
    .X(_04128_));
 sky130_fd_sc_hd__a22o_1 _08642_ (.A1(la_data_in[4]),
    .A2(_01147_),
    .B1(_01436_),
    .B2(\u_uart2wb.auto_baud_16x[0] ),
    .X(_04129_));
 sky130_fd_sc_hd__clkbuf_2 _08643_ (.A(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__xnor2_1 _08644_ (.A(_04038_),
    .B(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__clkbuf_1 _08645_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[0] ),
    .X(_04132_));
 sky130_fd_sc_hd__a211oi_1 _08646_ (.A1(_04128_),
    .A2(_04131_),
    .B1(_04061_),
    .C1(_04132_),
    .Y(_00872_));
 sky130_fd_sc_hd__nor2_1 _08647_ (.A(_04132_),
    .B(\u_uart2wb.u_core.u_clk_ctl.high_count[1] ),
    .Y(_04133_));
 sky130_fd_sc_hd__and2_1 _08648_ (.A(_04132_),
    .B(\u_uart2wb.u_core.u_clk_ctl.high_count[1] ),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_1 _08649_ (.A(_04129_),
    .X(_04135_));
 sky130_fd_sc_hd__and3_1 _08650_ (.A(_04037_),
    .B(_04045_),
    .C(_04135_),
    .X(_04136_));
 sky130_fd_sc_hd__a21oi_1 _08651_ (.A1(_04038_),
    .A2(_04130_),
    .B1(_04046_),
    .Y(_04137_));
 sky130_fd_sc_hd__nor2_1 _08652_ (.A(_04136_),
    .B(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__nand2_1 _08653_ (.A(_04128_),
    .B(_01825_),
    .Y(_04139_));
 sky130_fd_sc_hd__o221a_1 _08654_ (.A1(_04133_),
    .A2(_04134_),
    .B1(_04138_),
    .B2(_04088_),
    .C1(_04139_),
    .X(_00873_));
 sky130_fd_sc_hd__and2b_1 _08655_ (.A_N(\u_uart2wb.u_core.u_clk_ctl.high_count[2] ),
    .B(_04133_),
    .X(_04140_));
 sky130_fd_sc_hd__o21a_1 _08656_ (.A1(_04132_),
    .A2(\u_uart2wb.u_core.u_clk_ctl.high_count[1] ),
    .B1(\u_uart2wb.u_core.u_clk_ctl.high_count[2] ),
    .X(_04141_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08657_ (.A(_04129_),
    .X(_04142_));
 sky130_fd_sc_hd__nand2_1 _08658_ (.A(_04055_),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__o211a_1 _08659_ (.A1(_04054_),
    .A2(_04136_),
    .B1(_04143_),
    .C1(_04035_),
    .X(_04144_));
 sky130_fd_sc_hd__o22a_1 _08660_ (.A1(_04140_),
    .A2(_04141_),
    .B1(_04144_),
    .B2(_04089_),
    .X(_00874_));
 sky130_fd_sc_hd__xnor2_1 _08661_ (.A(_04066_),
    .B(_04143_),
    .Y(_04145_));
 sky130_fd_sc_hd__xor2_1 _08662_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[3] ),
    .B(_04140_),
    .X(_04146_));
 sky130_fd_sc_hd__o211a_1 _08663_ (.A1(_04071_),
    .A2(_04145_),
    .B1(_04146_),
    .C1(_04139_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _08664_ (.A0(_04074_),
    .A1(_04077_),
    .S(_04142_),
    .X(_04147_));
 sky130_fd_sc_hd__xnor2_1 _08665_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[4] ),
    .B(_01826_),
    .Y(_04148_));
 sky130_fd_sc_hd__o211a_1 _08666_ (.A1(_04071_),
    .A2(_04147_),
    .B1(_04148_),
    .C1(_04139_),
    .X(_00876_));
 sky130_fd_sc_hd__o21ai_1 _08667_ (.A1(\u_uart2wb.u_core.u_clk_ctl.high_count[4] ),
    .A2(_01826_),
    .B1(\u_uart2wb.u_core.u_clk_ctl.high_count[5] ),
    .Y(_04149_));
 sky130_fd_sc_hd__nand2_1 _08668_ (.A(_01827_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__mux2_1 _08669_ (.A0(_04082_),
    .A1(_04086_),
    .S(_04130_),
    .X(_04151_));
 sky130_fd_sc_hd__a22o_1 _08670_ (.A1(_04089_),
    .A2(_04150_),
    .B1(_04151_),
    .B2(_04121_),
    .X(_00877_));
 sky130_fd_sc_hd__nand2_1 _08671_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[6] ),
    .B(_01827_),
    .Y(_04152_));
 sky130_fd_sc_hd__clkbuf_1 _08672_ (.A(_04135_),
    .X(_04153_));
 sky130_fd_sc_hd__nand2_1 _08673_ (.A(_04093_),
    .B(_04142_),
    .Y(_04154_));
 sky130_fd_sc_hd__o211a_1 _08674_ (.A1(_04090_),
    .A2(_04153_),
    .B1(_04154_),
    .C1(_04035_),
    .X(_04155_));
 sky130_fd_sc_hd__o2bb2a_1 _08675_ (.A1_N(_01828_),
    .A2_N(_04152_),
    .B1(_04155_),
    .B2(_04089_),
    .X(_00878_));
 sky130_fd_sc_hd__xnor2_1 _08676_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[7] ),
    .B(_01828_),
    .Y(_04156_));
 sky130_fd_sc_hd__clkinv_2 _08677_ (.A(_04099_),
    .Y(_04157_));
 sky130_fd_sc_hd__mux2_1 _08678_ (.A0(_04157_),
    .A1(_04103_),
    .S(_04130_),
    .X(_04158_));
 sky130_fd_sc_hd__a22o_1 _08679_ (.A1(_04071_),
    .A2(_04156_),
    .B1(_04158_),
    .B2(_04121_),
    .X(_00879_));
 sky130_fd_sc_hd__o21ai_1 _08680_ (.A1(\u_uart2wb.u_core.u_clk_ctl.high_count[7] ),
    .A2(_01828_),
    .B1(\u_uart2wb.u_core.u_clk_ctl.high_count[8] ),
    .Y(_04159_));
 sky130_fd_sc_hd__a21oi_1 _08681_ (.A1(_04101_),
    .A2(_04135_),
    .B1(_04107_),
    .Y(_04160_));
 sky130_fd_sc_hd__a211o_1 _08682_ (.A1(_04117_),
    .A2(_04153_),
    .B1(_04160_),
    .C1(_01824_),
    .X(_04161_));
 sky130_fd_sc_hd__a22oi_1 _08683_ (.A1(_01829_),
    .A2(_04159_),
    .B1(_04161_),
    .B2(_04128_),
    .Y(_00880_));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[9] ),
    .B(_01829_),
    .Y(_04162_));
 sky130_fd_sc_hd__a21oi_1 _08685_ (.A1(_04117_),
    .A2(_04135_),
    .B1(_04118_),
    .Y(_04163_));
 sky130_fd_sc_hd__a311o_1 _08686_ (.A1(_04117_),
    .A2(_04118_),
    .A3(_04142_),
    .B1(_04163_),
    .C1(_01824_),
    .X(_04164_));
 sky130_fd_sc_hd__a22oi_1 _08687_ (.A1(_01830_),
    .A2(_04162_),
    .B1(_04164_),
    .B2(_04128_),
    .Y(_00881_));
 sky130_fd_sc_hd__and4_1 _08688_ (.A(_04101_),
    .B(_04107_),
    .C(_04118_),
    .D(_04129_),
    .X(_04165_));
 sky130_fd_sc_hd__o2bb2a_1 _08689_ (.A1_N(_04126_),
    .A2_N(_04153_),
    .B1(_04165_),
    .B2(_04123_),
    .X(_04166_));
 sky130_fd_sc_hd__nand2_1 _08690_ (.A(\u_uart2wb.u_core.u_clk_ctl.high_count[10] ),
    .B(_01830_),
    .Y(_04167_));
 sky130_fd_sc_hd__nand2_1 _08691_ (.A(_01831_),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__o211a_1 _08692_ (.A1(_04088_),
    .A2(_04166_),
    .B1(_04168_),
    .C1(_04139_),
    .X(_00882_));
 sky130_fd_sc_hd__a32o_1 _08693_ (.A1(_04080_),
    .A2(_04126_),
    .A3(_04153_),
    .B1(_01831_),
    .B2(\u_uart2wb.u_core.u_clk_ctl.high_count[11] ),
    .X(_00883_));
 sky130_fd_sc_hd__and3_1 _08694_ (.A(\u_uart2wb.u_aut_det.state[1] ),
    .B(net280),
    .C(_01178_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_2 _08695_ (.A(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__clkbuf_2 _08696_ (.A(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__mux2_1 _08697_ (.A0(\u_uart2wb.u_aut_det.ref2_cnt[0] ),
    .A1(_03688_),
    .S(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _08698_ (.A(_04172_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _08699_ (.A0(_01194_),
    .A1(_03690_),
    .S(_04171_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _08700_ (.A(_04173_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _08701_ (.A0(_01198_),
    .A1(\u_uart2wb.u_aut_det.clk_cnt[2] ),
    .S(_04171_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _08702_ (.A(_04174_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _08703_ (.A0(_01201_),
    .A1(_03693_),
    .S(_04171_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _08704_ (.A(_04175_),
    .X(_00887_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08705_ (.A(_04170_),
    .X(_04176_));
 sky130_fd_sc_hd__mux2_1 _08706_ (.A0(_01223_),
    .A1(\u_uart2wb.u_aut_det.clk_cnt[4] ),
    .S(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _08707_ (.A(_04177_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _08708_ (.A0(_01220_),
    .A1(_03698_),
    .S(_04176_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _08709_ (.A(_04178_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _08710_ (.A0(_01228_),
    .A1(_03700_),
    .S(_04176_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _08711_ (.A(_04179_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _08712_ (.A0(\u_uart2wb.u_aut_det.ref2_cnt[7] ),
    .A1(_03702_),
    .S(_04176_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _08713_ (.A(_04180_),
    .X(_00891_));
 sky130_fd_sc_hd__clkbuf_2 _08714_ (.A(_04170_),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _08715_ (.A0(_01331_),
    .A1(_03705_),
    .S(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__clkbuf_1 _08716_ (.A(_04182_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _08717_ (.A0(_01245_),
    .A1(_03707_),
    .S(_04181_),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _08718_ (.A(_04183_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _08719_ (.A0(_01335_),
    .A1(_03709_),
    .S(_04181_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _08720_ (.A(_04184_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _08721_ (.A0(_01256_),
    .A1(_03711_),
    .S(_04181_),
    .X(_04185_));
 sky130_fd_sc_hd__clkbuf_1 _08722_ (.A(_04185_),
    .X(_00895_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08723_ (.A(_04170_),
    .X(_04186_));
 sky130_fd_sc_hd__mux2_1 _08724_ (.A0(_01355_),
    .A1(_03714_),
    .S(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _08725_ (.A(_04187_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _08726_ (.A0(_01274_),
    .A1(_03716_),
    .S(_04186_),
    .X(_04188_));
 sky130_fd_sc_hd__clkbuf_1 _08727_ (.A(_04188_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _08728_ (.A0(_01359_),
    .A1(_03719_),
    .S(_04186_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _08729_ (.A(_04189_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _08730_ (.A0(_01268_),
    .A1(_03721_),
    .S(_04186_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _08731_ (.A(_04190_),
    .X(_00899_));
 sky130_fd_sc_hd__clkbuf_2 _08732_ (.A(_04169_),
    .X(_04191_));
 sky130_fd_sc_hd__mux2_1 _08733_ (.A0(_01343_),
    .A1(_03724_),
    .S(_04191_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _08734_ (.A(_04192_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _08735_ (.A0(_01296_),
    .A1(_03726_),
    .S(_04191_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _08736_ (.A(_04193_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _08737_ (.A0(_01282_),
    .A1(_03728_),
    .S(_04191_),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _08738_ (.A(_04194_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _08739_ (.A0(\u_uart2wb.u_aut_det.ref2_cnt[19] ),
    .A1(_03730_),
    .S(_04191_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _08740_ (.A(_04195_),
    .X(_00903_));
 sky130_fd_sc_hd__inv_2 _08741_ (.A(_02900_),
    .Y(_04196_));
 sky130_fd_sc_hd__nor2_1 _08742_ (.A(_04196_),
    .B(_02920_),
    .Y(_04197_));
 sky130_fd_sc_hd__inv_2 _08743_ (.A(_02919_),
    .Y(_04198_));
 sky130_fd_sc_hd__o31a_1 _08744_ (.A1(_02895_),
    .A2(_02961_),
    .A3(_02939_),
    .B1(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__or2_1 _08745_ (.A(_04197_),
    .B(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _08746_ (.A(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08747_ (.A(_04201_),
    .X(_04202_));
 sky130_fd_sc_hd__mux2_1 _08748_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[5] ),
    .A1(_02973_),
    .S(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_1 _08749_ (.A(_04203_),
    .X(_00904_));
 sky130_fd_sc_hd__a211o_1 _08750_ (.A1(_02877_),
    .A2(\u_uart2wb.u_msg.TxMsgBuf[5] ),
    .B1(_02935_),
    .C1(_02954_),
    .X(_04204_));
 sky130_fd_sc_hd__mux2_1 _08751_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[13] ),
    .A1(_04204_),
    .S(_04202_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_1 _08752_ (.A(_04205_),
    .X(_00905_));
 sky130_fd_sc_hd__nor2_1 _08753_ (.A(_04197_),
    .B(_04199_),
    .Y(_04206_));
 sky130_fd_sc_hd__clkbuf_1 _08754_ (.A(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _08755_ (.A(_04207_),
    .X(_04208_));
 sky130_fd_sc_hd__o21a_1 _08756_ (.A1(_02930_),
    .A2(_02940_),
    .B1(_04201_),
    .X(_04209_));
 sky130_fd_sc_hd__or2_1 _08757_ (.A(_04197_),
    .B(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__a21o_1 _08758_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[18] ),
    .A2(_04208_),
    .B1(_04210_),
    .X(_00906_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08759_ (.A(_04207_),
    .X(_04211_));
 sky130_fd_sc_hd__nor2_1 _08760_ (.A(_02936_),
    .B(_02920_),
    .Y(_04212_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08761_ (.A(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__a221o_1 _08762_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[17] ),
    .A2(_04211_),
    .B1(_04213_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[11] ),
    .C1(_04209_),
    .X(_00907_));
 sky130_fd_sc_hd__a221o_1 _08763_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[20] ),
    .A2(_04211_),
    .B1(_04213_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[12] ),
    .C1(_04210_),
    .X(_00908_));
 sky130_fd_sc_hd__clkbuf_1 _08764_ (.A(_04202_),
    .X(_04214_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08765_ (.A(_02936_),
    .X(_04215_));
 sky130_fd_sc_hd__or2_1 _08766_ (.A(_04215_),
    .B(_02920_),
    .X(_04216_));
 sky130_fd_sc_hd__o22a_1 _08767_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[21] ),
    .A2(_04214_),
    .B1(_04216_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[13] ),
    .X(_00909_));
 sky130_fd_sc_hd__nor2_1 _08768_ (.A(_03132_),
    .B(_02972_),
    .Y(_04217_));
 sky130_fd_sc_hd__and2_1 _08769_ (.A(_04217_),
    .B(_04200_),
    .X(_04218_));
 sky130_fd_sc_hd__a21o_1 _08770_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[12] ),
    .A2(_04208_),
    .B1(_04218_),
    .X(_00910_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08771_ (.A(_04197_),
    .X(_04219_));
 sky130_fd_sc_hd__a21o_1 _08772_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[24] ),
    .A2(_04208_),
    .B1(_04219_),
    .X(_00911_));
 sky130_fd_sc_hd__clkbuf_1 _08773_ (.A(_04212_),
    .X(_04220_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08774_ (.A(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08775_ (.A(_02939_),
    .X(_04222_));
 sky130_fd_sc_hd__and3_1 _08776_ (.A(_02954_),
    .B(_04222_),
    .C(_04198_),
    .X(_04223_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08777_ (.A(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__a221o_1 _08778_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[26] ),
    .A2(_04211_),
    .B1(_04221_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[18] ),
    .C1(_04224_),
    .X(_00912_));
 sky130_fd_sc_hd__clkbuf_1 _08779_ (.A(_04206_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _08780_ (.A(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__a221o_1 _08781_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[25] ),
    .A2(_04226_),
    .B1(_04221_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[17] ),
    .C1(_04224_),
    .X(_00913_));
 sky130_fd_sc_hd__a221o_1 _08782_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[28] ),
    .A2(_04226_),
    .B1(_04221_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[20] ),
    .C1(_04224_),
    .X(_00914_));
 sky130_fd_sc_hd__o22a_1 _08783_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[29] ),
    .A2(_04214_),
    .B1(_04216_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[21] ),
    .X(_00915_));
 sky130_fd_sc_hd__a221o_1 _08784_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[11] ),
    .A2(_04226_),
    .B1(_04221_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[12] ),
    .C1(_04219_),
    .X(_00916_));
 sky130_fd_sc_hd__clkbuf_1 _08785_ (.A(_04220_),
    .X(_04227_));
 sky130_fd_sc_hd__a221o_1 _08786_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[32] ),
    .A2(_04226_),
    .B1(_04227_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[24] ),
    .C1(_04218_),
    .X(_00917_));
 sky130_fd_sc_hd__clkbuf_1 _08787_ (.A(_04225_),
    .X(_04228_));
 sky130_fd_sc_hd__a221o_1 _08788_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[33] ),
    .A2(_04228_),
    .B1(_04227_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[25] ),
    .C1(_04224_),
    .X(_00918_));
 sky130_fd_sc_hd__a221o_1 _08789_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[34] ),
    .A2(_04228_),
    .B1(_04227_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[26] ),
    .C1(_04219_),
    .X(_00919_));
 sky130_fd_sc_hd__or2_1 _08790_ (.A(_04218_),
    .B(_04223_),
    .X(_04229_));
 sky130_fd_sc_hd__a221o_1 _08791_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[35] ),
    .A2(_04228_),
    .B1(_04227_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[25] ),
    .C1(_04229_),
    .X(_00920_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08792_ (.A(_04201_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _08793_ (.A(_04220_),
    .X(_04231_));
 sky130_fd_sc_hd__and2_1 _08794_ (.A(\u_uart2wb.u_msg.TxMsgBuf[36] ),
    .B(_04207_),
    .X(_04232_));
 sky130_fd_sc_hd__a221o_1 _08795_ (.A1(_02980_),
    .A2(_04230_),
    .B1(_04231_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[28] ),
    .C1(_04232_),
    .X(_00921_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08796_ (.A(_04206_),
    .X(_04233_));
 sky130_fd_sc_hd__a211o_1 _08797_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[29] ),
    .A2(_03139_),
    .B1(_02965_),
    .C1(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08798_ (.A(_04217_),
    .X(_04235_));
 sky130_fd_sc_hd__o22a_1 _08799_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[37] ),
    .A2(_04214_),
    .B1(_04234_),
    .B2(_04235_),
    .X(_00922_));
 sky130_fd_sc_hd__a221o_1 _08800_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[38] ),
    .A2(_04228_),
    .B1(_04231_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[11] ),
    .C1(_04219_),
    .X(_00923_));
 sky130_fd_sc_hd__clkbuf_1 _08801_ (.A(_04225_),
    .X(_04236_));
 sky130_fd_sc_hd__a221o_1 _08802_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[40] ),
    .A2(_04236_),
    .B1(_04231_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[32] ),
    .C1(_04209_),
    .X(_00924_));
 sky130_fd_sc_hd__a221o_1 _08803_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[41] ),
    .A2(_04236_),
    .B1(_04231_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[33] ),
    .C1(_04229_),
    .X(_00925_));
 sky130_fd_sc_hd__a22o_1 _08804_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[42] ),
    .A2(_04208_),
    .B1(_04213_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[34] ),
    .X(_00926_));
 sky130_fd_sc_hd__a22o_1 _08805_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[43] ),
    .A2(_04211_),
    .B1(_04213_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[35] ),
    .X(_00927_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08806_ (.A(_04212_),
    .X(_04237_));
 sky130_fd_sc_hd__a221o_1 _08807_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[44] ),
    .A2(_04236_),
    .B1(_04237_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[36] ),
    .C1(_04229_),
    .X(_00928_));
 sky130_fd_sc_hd__o22a_1 _08808_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[45] ),
    .A2(_04214_),
    .B1(_04216_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[37] ),
    .X(_00929_));
 sky130_fd_sc_hd__a221o_1 _08809_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[46] ),
    .A2(_04236_),
    .B1(_04237_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[38] ),
    .C1(_04210_),
    .X(_00930_));
 sky130_fd_sc_hd__a221o_1 _08810_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[48] ),
    .A2(_04233_),
    .B1(_04237_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[40] ),
    .C1(_04229_),
    .X(_00931_));
 sky130_fd_sc_hd__a211o_1 _08811_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[41] ),
    .A2(_03139_),
    .B1(_04222_),
    .C1(_04233_),
    .X(_04238_));
 sky130_fd_sc_hd__o22a_1 _08812_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[49] ),
    .A2(_04230_),
    .B1(_04238_),
    .B2(_04235_),
    .X(_00932_));
 sky130_fd_sc_hd__a211o_1 _08813_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[42] ),
    .A2(_03138_),
    .B1(_02963_),
    .C1(_04235_),
    .X(_04239_));
 sky130_fd_sc_hd__mux2_1 _08814_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[50] ),
    .A1(_04239_),
    .S(_04201_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _08815_ (.A(_04240_),
    .X(_00933_));
 sky130_fd_sc_hd__a211o_1 _08816_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[43] ),
    .A2(_02928_),
    .B1(_02950_),
    .C1(_04225_),
    .X(_04241_));
 sky130_fd_sc_hd__o22a_1 _08817_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[51] ),
    .A2(_04230_),
    .B1(_04241_),
    .B2(_04235_),
    .X(_00934_));
 sky130_fd_sc_hd__and2_1 _08818_ (.A(\u_uart2wb.u_msg.TxMsgBuf[52] ),
    .B(_04207_),
    .X(_04242_));
 sky130_fd_sc_hd__a221o_1 _08819_ (.A1(_04222_),
    .A2(_04202_),
    .B1(_04237_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[44] ),
    .C1(_04242_),
    .X(_00935_));
 sky130_fd_sc_hd__o22a_1 _08820_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[53] ),
    .A2(_04230_),
    .B1(_04216_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[45] ),
    .X(_00936_));
 sky130_fd_sc_hd__a221o_1 _08821_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[54] ),
    .A2(_04233_),
    .B1(_04220_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[46] ),
    .C1(_04210_),
    .X(_00937_));
 sky130_fd_sc_hd__a22o_1 _08822_ (.A1(net21),
    .A2(_02695_),
    .B1(_02697_),
    .B2(_02525_),
    .X(_00938_));
 sky130_fd_sc_hd__o22a_1 _08823_ (.A1(net22),
    .A2(_03596_),
    .B1(_03597_),
    .B2(_03227_),
    .X(_00939_));
 sky130_fd_sc_hd__o22a_1 _08824_ (.A1(net24),
    .A2(_02698_),
    .B1(_02700_),
    .B2(_02529_),
    .X(_00940_));
 sky130_fd_sc_hd__a22o_1 _08825_ (.A1(net25),
    .A2(_02695_),
    .B1(_02697_),
    .B2(_02531_),
    .X(_00941_));
 sky130_fd_sc_hd__and2_1 _08826_ (.A(_02171_),
    .B(_03178_),
    .X(_04243_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08827_ (.A(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__mux2_1 _08828_ (.A0(\u_reg.cfg_glb_ctrl[0] ),
    .A1(_02285_),
    .S(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _08829_ (.A(_04245_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _08830_ (.A0(\u_reg.cfg_glb_ctrl[1] ),
    .A1(_02265_),
    .S(_04244_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _08831_ (.A(_04246_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _08832_ (.A0(\u_reg.cfg_glb_ctrl[2] ),
    .A1(_02258_),
    .S(_04244_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _08833_ (.A(_04247_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _08834_ (.A0(\u_reg.cfg_glb_ctrl[3] ),
    .A1(_02253_),
    .S(_04244_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _08835_ (.A(_04248_),
    .X(_00945_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08836_ (.A(_04243_),
    .X(_04249_));
 sky130_fd_sc_hd__mux2_1 _08837_ (.A0(\u_reg.cfg_glb_ctrl[4] ),
    .A1(_02245_),
    .S(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _08838_ (.A(_04250_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _08839_ (.A0(\u_reg.cfg_glb_ctrl[5] ),
    .A1(_02238_),
    .S(_04249_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _08840_ (.A(_04251_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _08841_ (.A0(\u_reg.cfg_glb_ctrl[6] ),
    .A1(_02233_),
    .S(_04249_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _08842_ (.A(_04252_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _08843_ (.A0(\u_reg.cfg_glb_ctrl[7] ),
    .A1(_02227_),
    .S(_04249_),
    .X(_04253_));
 sky130_fd_sc_hd__clkbuf_1 _08844_ (.A(_04253_),
    .X(_00949_));
 sky130_fd_sc_hd__clkbuf_1 _08845_ (.A(_01137_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _08846_ (.A(_03933_),
    .X(_04255_));
 sky130_fd_sc_hd__o211a_1 _08847_ (.A1(_04254_),
    .A2(_01184_),
    .B1(_04255_),
    .C1(_01140_),
    .X(_04256_));
 sky130_fd_sc_hd__a21oi_1 _08848_ (.A1(_04254_),
    .A2(_04255_),
    .B1(_01140_),
    .Y(_04257_));
 sky130_fd_sc_hd__nor2_1 _08849_ (.A(_04256_),
    .B(_04257_),
    .Y(_00950_));
 sky130_fd_sc_hd__o21ai_1 _08850_ (.A1(_01137_),
    .A2(_01184_),
    .B1(_04255_),
    .Y(_04258_));
 sky130_fd_sc_hd__a21o_1 _08851_ (.A1(_04254_),
    .A2(_01141_),
    .B1(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__o21a_1 _08852_ (.A1(_01139_),
    .A2(_04256_),
    .B1(_04259_),
    .X(_00951_));
 sky130_fd_sc_hd__nor2_1 _08853_ (.A(_01136_),
    .B(_01141_),
    .Y(_04260_));
 sky130_fd_sc_hd__a32o_1 _08854_ (.A1(_04254_),
    .A2(_04255_),
    .A3(_04260_),
    .B1(_04259_),
    .B2(_01136_),
    .X(_00952_));
 sky130_fd_sc_hd__nor2_1 _08855_ (.A(_02935_),
    .B(_02914_),
    .Y(_04261_));
 sky130_fd_sc_hd__clkbuf_2 _08856_ (.A(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__or3_1 _08857_ (.A(\u_uart2wb.rx_data[4] ),
    .B(\u_uart2wb.rx_data[7] ),
    .C(\u_uart2wb.rx_data[6] ),
    .X(_04263_));
 sky130_fd_sc_hd__or3b_1 _08858_ (.A(\u_uart2wb.rx_data[1] ),
    .B(\u_uart2wb.rx_data[0] ),
    .C_N(\u_uart2wb.rx_data[5] ),
    .X(_04264_));
 sky130_fd_sc_hd__nor4_2 _08859_ (.A(_04010_),
    .B(\u_uart2wb.rx_data[3] ),
    .C(_04263_),
    .D(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__or2b_1 _08860_ (.A(\u_uart2wb.rx_data[2] ),
    .B_N(\u_uart2wb.rx_data[3] ),
    .X(_04266_));
 sky130_fd_sc_hd__or2b_1 _08861_ (.A(\u_uart2wb.rx_data[0] ),
    .B_N(_04006_),
    .X(_04267_));
 sky130_fd_sc_hd__or4_1 _08862_ (.A(_04023_),
    .B(_04263_),
    .C(_04266_),
    .D(_04267_),
    .X(_04268_));
 sky130_fd_sc_hd__and2b_1 _08863_ (.A_N(_04265_),
    .B(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__or3_1 _08864_ (.A(\u_uart2wb.u_msg.RxMsgCnt[4] ),
    .B(\u_uart2wb.u_msg.RxMsgCnt[3] ),
    .C(\u_uart2wb.u_msg.RxMsgCnt[1] ),
    .X(_04270_));
 sky130_fd_sc_hd__nor3_1 _08865_ (.A(\u_uart2wb.u_msg.RxMsgCnt[2] ),
    .B(\u_uart2wb.u_msg.RxMsgCnt[0] ),
    .C(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__nor2_1 _08866_ (.A(_04269_),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__inv_2 _08867_ (.A(\u_uart2wb.rx_wr ),
    .Y(_04273_));
 sky130_fd_sc_hd__and2_1 _08868_ (.A(_04265_),
    .B(_04271_),
    .X(_04274_));
 sky130_fd_sc_hd__or2_1 _08869_ (.A(_02897_),
    .B(_02913_),
    .X(_04275_));
 sky130_fd_sc_hd__or3_1 _08870_ (.A(_04273_),
    .B(_04274_),
    .C(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__nor2_1 _08871_ (.A(_04272_),
    .B(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _08872_ (.A(_04273_),
    .X(_04278_));
 sky130_fd_sc_hd__clkbuf_1 _08873_ (.A(_02914_),
    .X(_04279_));
 sky130_fd_sc_hd__nor2_1 _08874_ (.A(_02898_),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__a21o_1 _08875_ (.A1(_04278_),
    .A2(_04280_),
    .B1(_02917_),
    .X(_04281_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08876_ (.A(_04268_),
    .X(_04282_));
 sky130_fd_sc_hd__nand2_1 _08877_ (.A(\u_uart2wb.u_msg.cmd[6] ),
    .B(\u_uart2wb.u_msg.cmd[9] ),
    .Y(_04283_));
 sky130_fd_sc_hd__and4b_1 _08878_ (.A_N(\u_uart2wb.u_msg.cmd[4] ),
    .B(\u_uart2wb.u_msg.cmd[5] ),
    .C(\u_uart2wb.u_msg.cmd[2] ),
    .D(\u_uart2wb.u_msg.cmd[3] ),
    .X(_04284_));
 sky130_fd_sc_hd__nand3b_1 _08879_ (.A_N(\u_uart2wb.u_msg.cmd[1] ),
    .B(\u_uart2wb.u_msg.cmd[0] ),
    .C(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__nand4b_1 _08880_ (.A_N(\u_uart2wb.u_msg.cmd[15] ),
    .B(\u_uart2wb.u_msg.cmd[14] ),
    .C(\u_uart2wb.u_msg.cmd[12] ),
    .D(\u_uart2wb.u_msg.cmd[13] ),
    .Y(_04286_));
 sky130_fd_sc_hd__or4_1 _08881_ (.A(\u_uart2wb.u_msg.cmd[7] ),
    .B(\u_uart2wb.u_msg.cmd[11] ),
    .C(_04285_),
    .D(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__or4_1 _08882_ (.A(\u_uart2wb.u_msg.cmd[8] ),
    .B(\u_uart2wb.u_msg.cmd[10] ),
    .C(_04283_),
    .D(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__nor2_1 _08883_ (.A(_04282_),
    .B(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__nor2_1 _08884_ (.A(_04276_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _08885_ (.A(_04272_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _08886_ (.A(_04265_),
    .X(_04292_));
 sky130_fd_sc_hd__or4bb_1 _08887_ (.A(\u_uart2wb.u_msg.cmd[7] ),
    .B(\u_uart2wb.u_msg.cmd[11] ),
    .C_N(\u_uart2wb.u_msg.cmd[9] ),
    .D_N(\u_uart2wb.u_msg.cmd[6] ),
    .X(_04293_));
 sky130_fd_sc_hd__or3_1 _08888_ (.A(_04285_),
    .B(_04286_),
    .C(_04293_),
    .X(_04294_));
 sky130_fd_sc_hd__clkinv_2 _08889_ (.A(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__and3_1 _08890_ (.A(\u_uart2wb.u_msg.cmd[8] ),
    .B(\u_uart2wb.u_msg.cmd[10] ),
    .C(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__and3_1 _08891_ (.A(_03984_),
    .B(_04292_),
    .C(_04296_),
    .X(_04297_));
 sky130_fd_sc_hd__and3_1 _08892_ (.A(_03983_),
    .B(_04265_),
    .C(_04261_),
    .X(_04298_));
 sky130_fd_sc_hd__o21a_1 _08893_ (.A1(_04278_),
    .A2(_04269_),
    .B1(_04261_),
    .X(_04299_));
 sky130_fd_sc_hd__a31o_1 _08894_ (.A1(_03983_),
    .A2(_04274_),
    .A3(_04280_),
    .B1(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__or2_1 _08895_ (.A(_04298_),
    .B(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__a31o_1 _08896_ (.A1(_04291_),
    .A2(_04280_),
    .A3(_04297_),
    .B1(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__or4_1 _08897_ (.A(_04277_),
    .B(_04281_),
    .C(_04290_),
    .D(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__or2_1 _08898_ (.A(_02899_),
    .B(_04279_),
    .X(_04304_));
 sky130_fd_sc_hd__nor2_1 _08899_ (.A(_04303_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__mux2_1 _08900_ (.A0(\u_uart2wb.reg_wr ),
    .A1(_04262_),
    .S(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_1 _08901_ (.A(_04306_),
    .X(_00953_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08902_ (.A(_04280_),
    .X(_04307_));
 sky130_fd_sc_hd__nor2_1 _08903_ (.A(_02875_),
    .B(_02914_),
    .Y(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _08904_ (.A(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__and2b_1 _08905_ (.A_N(_04271_),
    .B(_04292_),
    .X(_04310_));
 sky130_fd_sc_hd__and2_1 _08906_ (.A(_04309_),
    .B(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__or2_1 _08907_ (.A(_04277_),
    .B(_04304_),
    .X(_04312_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08908_ (.A(_04282_),
    .X(_04313_));
 sky130_fd_sc_hd__o2111ai_4 _08909_ (.A1(_04307_),
    .A2(_04311_),
    .B1(_04312_),
    .C1(_03984_),
    .D1(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _08910_ (.A(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08911_ (.A(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__inv_2 _08912_ (.A(_04023_),
    .Y(_04317_));
 sky130_fd_sc_hd__or3b_1 _08913_ (.A(_04029_),
    .B(_04026_),
    .C_N(_04019_),
    .X(_04318_));
 sky130_fd_sc_hd__nor3_1 _08914_ (.A(_04014_),
    .B(_04317_),
    .C(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__or3b_1 _08915_ (.A(_04019_),
    .B(_04029_),
    .C_N(_04026_),
    .X(_04320_));
 sky130_fd_sc_hd__or3b_1 _08916_ (.A(_04014_),
    .B(_04320_),
    .C_N(_04010_),
    .X(_04321_));
 sky130_fd_sc_hd__or3_1 _08917_ (.A(_04006_),
    .B(_04001_),
    .C(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__or2b_1 _08918_ (.A(_04006_),
    .B_N(_04001_),
    .X(_04323_));
 sky130_fd_sc_hd__or4_1 _08919_ (.A(_04317_),
    .B(_04266_),
    .C(_04323_),
    .D(_04318_),
    .X(_04324_));
 sky130_fd_sc_hd__nand2_1 _08920_ (.A(_04322_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__or3_2 _08921_ (.A(_04010_),
    .B(_04014_),
    .C(_04320_),
    .X(_04326_));
 sky130_fd_sc_hd__nor2_1 _08922_ (.A(_04267_),
    .B(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__nor2_1 _08923_ (.A(_04321_),
    .B(_04323_),
    .Y(_04328_));
 sky130_fd_sc_hd__nor3_1 _08924_ (.A(_04011_),
    .B(_04015_),
    .C(_04320_),
    .Y(_04329_));
 sky130_fd_sc_hd__nor3_1 _08925_ (.A(_04264_),
    .B(_04266_),
    .C(_04318_),
    .Y(_04330_));
 sky130_fd_sc_hd__a2111o_1 _08926_ (.A1(_04001_),
    .A2(_04329_),
    .B1(_04330_),
    .C1(_04319_),
    .D1(_04325_),
    .X(_04331_));
 sky130_fd_sc_hd__nor3_1 _08927_ (.A(_04327_),
    .B(_04328_),
    .C(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__a2111o_2 _08928_ (.A1(_04002_),
    .A2(_04319_),
    .B1(_04325_),
    .C1(_04332_),
    .D1(_04327_),
    .X(_04333_));
 sky130_fd_sc_hd__nor2_1 _08929_ (.A(_04275_),
    .B(_04314_),
    .Y(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _08930_ (.A(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__a22o_1 _08931_ (.A1(\u_uart2wb.reg_addr[0] ),
    .A2(_04316_),
    .B1(_04333_),
    .B2(_04335_),
    .X(_00954_));
 sky130_fd_sc_hd__clkbuf_1 _08932_ (.A(_04334_),
    .X(_04336_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08933_ (.A(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__nand2_1 _08934_ (.A(_04007_),
    .B(_04319_),
    .Y(_04338_));
 sky130_fd_sc_hd__o211ai_4 _08935_ (.A1(_04326_),
    .A2(_04323_),
    .B1(_04331_),
    .C1(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__a22o_1 _08936_ (.A1(\u_uart2wb.reg_addr[1] ),
    .A2(_04316_),
    .B1(_04337_),
    .B2(_04339_),
    .X(_00955_));
 sky130_fd_sc_hd__a311o_2 _08937_ (.A1(_04007_),
    .A2(_04002_),
    .A3(_04329_),
    .B1(_04332_),
    .C1(_04011_),
    .X(_04340_));
 sky130_fd_sc_hd__a22o_1 _08938_ (.A1(\u_uart2wb.reg_addr[2] ),
    .A2(_04316_),
    .B1(_04337_),
    .B2(_04340_),
    .X(_00956_));
 sky130_fd_sc_hd__or3_2 _08939_ (.A(_04015_),
    .B(_04317_),
    .C(_04318_),
    .X(_04341_));
 sky130_fd_sc_hd__a22o_1 _08940_ (.A1(\u_uart2wb.reg_addr[3] ),
    .A2(_04316_),
    .B1(_04341_),
    .B2(_04335_),
    .X(_00957_));
 sky130_fd_sc_hd__clkbuf_1 _08941_ (.A(_04315_),
    .X(_04342_));
 sky130_fd_sc_hd__a22o_1 _08942_ (.A1(\u_uart2wb.reg_addr[4] ),
    .A2(_04342_),
    .B1(_04337_),
    .B2(\u_uart2wb.reg_addr[0] ),
    .X(_00958_));
 sky130_fd_sc_hd__a22o_1 _08943_ (.A1(\u_uart2wb.reg_addr[5] ),
    .A2(_04342_),
    .B1(_04337_),
    .B2(\u_uart2wb.reg_addr[1] ),
    .X(_00959_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08944_ (.A(_04336_),
    .X(_04343_));
 sky130_fd_sc_hd__a22o_1 _08945_ (.A1(\u_uart2wb.reg_addr[6] ),
    .A2(_04342_),
    .B1(_04343_),
    .B2(\u_uart2wb.reg_addr[2] ),
    .X(_00960_));
 sky130_fd_sc_hd__a22o_1 _08946_ (.A1(\u_uart2wb.reg_addr[7] ),
    .A2(_04342_),
    .B1(_04343_),
    .B2(\u_uart2wb.reg_addr[3] ),
    .X(_00961_));
 sky130_fd_sc_hd__clkbuf_1 _08947_ (.A(_04315_),
    .X(_04344_));
 sky130_fd_sc_hd__a22o_1 _08948_ (.A1(\u_uart2wb.reg_addr[8] ),
    .A2(_04344_),
    .B1(_04343_),
    .B2(\u_uart2wb.reg_addr[4] ),
    .X(_00962_));
 sky130_fd_sc_hd__a22o_1 _08949_ (.A1(\u_uart2wb.reg_addr[9] ),
    .A2(_04344_),
    .B1(_04343_),
    .B2(\u_uart2wb.reg_addr[5] ),
    .X(_00963_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08950_ (.A(_04336_),
    .X(_04345_));
 sky130_fd_sc_hd__a22o_1 _08951_ (.A1(\u_uart2wb.reg_addr[10] ),
    .A2(_04344_),
    .B1(_04345_),
    .B2(\u_uart2wb.reg_addr[6] ),
    .X(_00964_));
 sky130_fd_sc_hd__a22o_1 _08952_ (.A1(\u_uart2wb.reg_addr[11] ),
    .A2(_04344_),
    .B1(_04345_),
    .B2(\u_uart2wb.reg_addr[7] ),
    .X(_00965_));
 sky130_fd_sc_hd__clkbuf_1 _08953_ (.A(_04315_),
    .X(_04346_));
 sky130_fd_sc_hd__a22o_1 _08954_ (.A1(\u_uart2wb.reg_addr[12] ),
    .A2(_04346_),
    .B1(_04345_),
    .B2(\u_uart2wb.reg_addr[8] ),
    .X(_00966_));
 sky130_fd_sc_hd__a22o_1 _08955_ (.A1(\u_uart2wb.reg_addr[13] ),
    .A2(_04346_),
    .B1(_04345_),
    .B2(\u_uart2wb.reg_addr[9] ),
    .X(_00967_));
 sky130_fd_sc_hd__clkbuf_1 _08956_ (.A(_04336_),
    .X(_04347_));
 sky130_fd_sc_hd__a22o_1 _08957_ (.A1(\u_uart2wb.reg_addr[14] ),
    .A2(_04346_),
    .B1(_04347_),
    .B2(\u_uart2wb.reg_addr[10] ),
    .X(_00968_));
 sky130_fd_sc_hd__a22o_1 _08958_ (.A1(\u_uart2wb.reg_addr[15] ),
    .A2(_04346_),
    .B1(_04347_),
    .B2(\u_uart2wb.reg_addr[11] ),
    .X(_00969_));
 sky130_fd_sc_hd__clkbuf_1 _08959_ (.A(_04314_),
    .X(_04348_));
 sky130_fd_sc_hd__a22o_1 _08960_ (.A1(\u_uart2wb.reg_addr[16] ),
    .A2(_04348_),
    .B1(_04347_),
    .B2(\u_uart2wb.reg_addr[12] ),
    .X(_00970_));
 sky130_fd_sc_hd__a22o_1 _08961_ (.A1(\u_uart2wb.reg_addr[17] ),
    .A2(_04348_),
    .B1(_04347_),
    .B2(\u_uart2wb.reg_addr[13] ),
    .X(_00971_));
 sky130_fd_sc_hd__a22o_1 _08962_ (.A1(\u_uart2wb.reg_addr[18] ),
    .A2(_04348_),
    .B1(_04335_),
    .B2(\u_uart2wb.reg_addr[14] ),
    .X(_00972_));
 sky130_fd_sc_hd__a22o_1 _08963_ (.A1(\u_uart2wb.reg_addr[19] ),
    .A2(_04348_),
    .B1(_04335_),
    .B2(\u_uart2wb.reg_addr[15] ),
    .X(_00973_));
 sky130_fd_sc_hd__a21bo_1 _08964_ (.A1(_04292_),
    .A2(_04296_),
    .B1_N(_04272_),
    .X(_04349_));
 sky130_fd_sc_hd__a21o_1 _08965_ (.A1(_02901_),
    .A2(_04282_),
    .B1(_04291_),
    .X(_04350_));
 sky130_fd_sc_hd__nand2_1 _08966_ (.A(_04349_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__or4_4 _08967_ (.A(_04278_),
    .B(_04298_),
    .C(_04312_),
    .D(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08968_ (.A(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _08969_ (.A(_04353_),
    .X(_04354_));
 sky130_fd_sc_hd__inv_2 _08970_ (.A(_04262_),
    .Y(_04355_));
 sky130_fd_sc_hd__nor2_1 _08971_ (.A(_04355_),
    .B(_04352_),
    .Y(_04356_));
 sky130_fd_sc_hd__clkbuf_1 _08972_ (.A(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _08973_ (.A(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__a22o_1 _08974_ (.A1(\u_uart2wb.reg_wdata[0] ),
    .A2(_04354_),
    .B1(_04358_),
    .B2(_04333_),
    .X(_00974_));
 sky130_fd_sc_hd__a22o_1 _08975_ (.A1(\u_uart2wb.reg_wdata[1] ),
    .A2(_04354_),
    .B1(_04358_),
    .B2(_04339_),
    .X(_00975_));
 sky130_fd_sc_hd__a22o_1 _08976_ (.A1(\u_uart2wb.reg_wdata[2] ),
    .A2(_04354_),
    .B1(_04358_),
    .B2(_04340_),
    .X(_00976_));
 sky130_fd_sc_hd__a22o_1 _08977_ (.A1(\u_uart2wb.reg_wdata[3] ),
    .A2(_04354_),
    .B1(_04358_),
    .B2(_04341_),
    .X(_00977_));
 sky130_fd_sc_hd__clkbuf_1 _08978_ (.A(_04353_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _08979_ (.A(_04357_),
    .X(_04360_));
 sky130_fd_sc_hd__a22o_1 _08980_ (.A1(\u_uart2wb.reg_wdata[4] ),
    .A2(_04359_),
    .B1(_04360_),
    .B2(\u_uart2wb.reg_wdata[0] ),
    .X(_00978_));
 sky130_fd_sc_hd__a22o_1 _08981_ (.A1(\u_uart2wb.reg_wdata[5] ),
    .A2(_04359_),
    .B1(_04360_),
    .B2(\u_uart2wb.reg_wdata[1] ),
    .X(_00979_));
 sky130_fd_sc_hd__a22o_1 _08982_ (.A1(\u_uart2wb.reg_wdata[6] ),
    .A2(_04359_),
    .B1(_04360_),
    .B2(\u_uart2wb.reg_wdata[2] ),
    .X(_00980_));
 sky130_fd_sc_hd__a22o_1 _08983_ (.A1(\u_uart2wb.reg_wdata[7] ),
    .A2(_04359_),
    .B1(_04360_),
    .B2(\u_uart2wb.reg_wdata[3] ),
    .X(_00981_));
 sky130_fd_sc_hd__clkbuf_1 _08984_ (.A(_04353_),
    .X(_04361_));
 sky130_fd_sc_hd__clkbuf_1 _08985_ (.A(_04357_),
    .X(_04362_));
 sky130_fd_sc_hd__a22o_1 _08986_ (.A1(\u_uart2wb.reg_wdata[8] ),
    .A2(_04361_),
    .B1(_04362_),
    .B2(\u_uart2wb.reg_wdata[4] ),
    .X(_00982_));
 sky130_fd_sc_hd__a22o_1 _08987_ (.A1(\u_uart2wb.reg_wdata[9] ),
    .A2(_04361_),
    .B1(_04362_),
    .B2(\u_uart2wb.reg_wdata[5] ),
    .X(_00983_));
 sky130_fd_sc_hd__a22o_1 _08988_ (.A1(\u_uart2wb.reg_wdata[10] ),
    .A2(_04361_),
    .B1(_04362_),
    .B2(\u_uart2wb.reg_wdata[6] ),
    .X(_00984_));
 sky130_fd_sc_hd__a22o_1 _08989_ (.A1(\u_uart2wb.reg_wdata[11] ),
    .A2(_04361_),
    .B1(_04362_),
    .B2(\u_uart2wb.reg_wdata[7] ),
    .X(_00985_));
 sky130_fd_sc_hd__clkbuf_1 _08990_ (.A(_04353_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _08991_ (.A(_04357_),
    .X(_04364_));
 sky130_fd_sc_hd__a22o_1 _08992_ (.A1(\u_uart2wb.reg_wdata[12] ),
    .A2(_04363_),
    .B1(_04364_),
    .B2(\u_uart2wb.reg_wdata[8] ),
    .X(_00986_));
 sky130_fd_sc_hd__a22o_1 _08993_ (.A1(\u_uart2wb.reg_wdata[13] ),
    .A2(_04363_),
    .B1(_04364_),
    .B2(\u_uart2wb.reg_wdata[9] ),
    .X(_00987_));
 sky130_fd_sc_hd__a22o_1 _08994_ (.A1(\u_uart2wb.reg_wdata[14] ),
    .A2(_04363_),
    .B1(_04364_),
    .B2(\u_uart2wb.reg_wdata[10] ),
    .X(_00988_));
 sky130_fd_sc_hd__a22o_1 _08995_ (.A1(\u_uart2wb.reg_wdata[15] ),
    .A2(_04363_),
    .B1(_04364_),
    .B2(\u_uart2wb.reg_wdata[11] ),
    .X(_00989_));
 sky130_fd_sc_hd__clkbuf_1 _08996_ (.A(_04352_),
    .X(_04365_));
 sky130_fd_sc_hd__clkbuf_1 _08997_ (.A(_04365_),
    .X(_04366_));
 sky130_fd_sc_hd__clkbuf_1 _08998_ (.A(_04356_),
    .X(_04367_));
 sky130_fd_sc_hd__clkbuf_1 _08999_ (.A(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__a22o_1 _09000_ (.A1(\u_uart2wb.reg_wdata[16] ),
    .A2(_04366_),
    .B1(_04368_),
    .B2(\u_uart2wb.reg_wdata[12] ),
    .X(_00990_));
 sky130_fd_sc_hd__a22o_1 _09001_ (.A1(\u_uart2wb.reg_wdata[17] ),
    .A2(_04366_),
    .B1(_04368_),
    .B2(\u_uart2wb.reg_wdata[13] ),
    .X(_00991_));
 sky130_fd_sc_hd__a22o_1 _09002_ (.A1(\u_uart2wb.reg_wdata[18] ),
    .A2(_04366_),
    .B1(_04368_),
    .B2(\u_uart2wb.reg_wdata[14] ),
    .X(_00992_));
 sky130_fd_sc_hd__a22o_1 _09003_ (.A1(\u_uart2wb.reg_wdata[19] ),
    .A2(_04366_),
    .B1(_04368_),
    .B2(\u_uart2wb.reg_wdata[15] ),
    .X(_00993_));
 sky130_fd_sc_hd__clkbuf_1 _09004_ (.A(_04365_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _09005_ (.A(_04367_),
    .X(_04370_));
 sky130_fd_sc_hd__a22o_1 _09006_ (.A1(\u_uart2wb.reg_wdata[20] ),
    .A2(_04369_),
    .B1(_04370_),
    .B2(\u_uart2wb.reg_wdata[16] ),
    .X(_00994_));
 sky130_fd_sc_hd__a22o_1 _09007_ (.A1(\u_uart2wb.reg_wdata[21] ),
    .A2(_04369_),
    .B1(_04370_),
    .B2(\u_uart2wb.reg_wdata[17] ),
    .X(_00995_));
 sky130_fd_sc_hd__a22o_1 _09008_ (.A1(\u_uart2wb.reg_wdata[22] ),
    .A2(_04369_),
    .B1(_04370_),
    .B2(\u_uart2wb.reg_wdata[18] ),
    .X(_00996_));
 sky130_fd_sc_hd__a22o_1 _09009_ (.A1(\u_uart2wb.reg_wdata[23] ),
    .A2(_04369_),
    .B1(_04370_),
    .B2(\u_uart2wb.reg_wdata[19] ),
    .X(_00997_));
 sky130_fd_sc_hd__clkbuf_1 _09010_ (.A(_04365_),
    .X(_04371_));
 sky130_fd_sc_hd__clkbuf_1 _09011_ (.A(_04367_),
    .X(_04372_));
 sky130_fd_sc_hd__a22o_1 _09012_ (.A1(\u_uart2wb.reg_wdata[24] ),
    .A2(_04371_),
    .B1(_04372_),
    .B2(\u_uart2wb.reg_wdata[20] ),
    .X(_00998_));
 sky130_fd_sc_hd__a22o_1 _09013_ (.A1(\u_uart2wb.reg_wdata[25] ),
    .A2(_04371_),
    .B1(_04372_),
    .B2(\u_uart2wb.reg_wdata[21] ),
    .X(_00999_));
 sky130_fd_sc_hd__a22o_1 _09014_ (.A1(\u_uart2wb.reg_wdata[26] ),
    .A2(_04371_),
    .B1(_04372_),
    .B2(\u_uart2wb.reg_wdata[22] ),
    .X(_01000_));
 sky130_fd_sc_hd__a22o_1 _09015_ (.A1(\u_uart2wb.reg_wdata[27] ),
    .A2(_04371_),
    .B1(_04372_),
    .B2(\u_uart2wb.reg_wdata[23] ),
    .X(_01001_));
 sky130_fd_sc_hd__clkbuf_1 _09016_ (.A(_04365_),
    .X(_04373_));
 sky130_fd_sc_hd__clkbuf_1 _09017_ (.A(_04367_),
    .X(_04374_));
 sky130_fd_sc_hd__a22o_1 _09018_ (.A1(\u_uart2wb.reg_wdata[28] ),
    .A2(_04373_),
    .B1(_04374_),
    .B2(\u_uart2wb.reg_wdata[24] ),
    .X(_01002_));
 sky130_fd_sc_hd__a22o_1 _09019_ (.A1(\u_uart2wb.reg_wdata[29] ),
    .A2(_04373_),
    .B1(_04374_),
    .B2(\u_uart2wb.reg_wdata[25] ),
    .X(_01003_));
 sky130_fd_sc_hd__a22o_1 _09020_ (.A1(\u_uart2wb.reg_wdata[30] ),
    .A2(_04373_),
    .B1(_04374_),
    .B2(\u_uart2wb.reg_wdata[26] ),
    .X(_01004_));
 sky130_fd_sc_hd__a22o_1 _09021_ (.A1(\u_uart2wb.reg_wdata[31] ),
    .A2(_04373_),
    .B1(_04374_),
    .B2(\u_uart2wb.reg_wdata[27] ),
    .X(_01005_));
 sky130_fd_sc_hd__o22a_1 _09022_ (.A1(_02916_),
    .A2(_04303_),
    .B1(_04305_),
    .B2(\u_uart2wb.reg_req ),
    .X(_01006_));
 sky130_fd_sc_hd__o21a_1 _09023_ (.A1(\u_uart2wb.u_msg.TxMsgSize[4] ),
    .A2(_02911_),
    .B1(_02895_),
    .X(_04375_));
 sky130_fd_sc_hd__o21a_1 _09024_ (.A1(_02909_),
    .A2(_02917_),
    .B1(\u_uart2wb.tx_data_avail ),
    .X(_04376_));
 sky130_fd_sc_hd__or2_1 _09025_ (.A(_04375_),
    .B(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_1 _09026_ (.A(_04377_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _09027_ (.A0(\u_uart2wb.tx_data[0] ),
    .A1(\u_uart2wb.u_core.u_txfsm.txdata[0] ),
    .S(_01161_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _09028_ (.A(_04378_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _09029_ (.A0(\u_uart2wb.tx_data[1] ),
    .A1(\u_uart2wb.u_core.u_txfsm.txdata[1] ),
    .S(_01161_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _09030_ (.A(_04379_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _09031_ (.A0(\u_uart2wb.tx_data[2] ),
    .A1(\u_uart2wb.u_core.u_txfsm.txdata[2] ),
    .S(_01161_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_1 _09032_ (.A(_04380_),
    .X(_01010_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09033_ (.A(_01160_),
    .X(_04381_));
 sky130_fd_sc_hd__mux2_1 _09034_ (.A0(\u_uart2wb.tx_data[3] ),
    .A1(\u_uart2wb.u_core.u_txfsm.txdata[3] ),
    .S(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _09035_ (.A(_04382_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _09036_ (.A0(\u_uart2wb.tx_data[4] ),
    .A1(\u_uart2wb.u_core.u_txfsm.txdata[4] ),
    .S(_04381_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _09037_ (.A(_04383_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _09038_ (.A0(\u_uart2wb.tx_data[5] ),
    .A1(\u_uart2wb.u_core.u_txfsm.txdata[5] ),
    .S(_04381_),
    .X(_04384_));
 sky130_fd_sc_hd__clkbuf_1 _09039_ (.A(_04384_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _09040_ (.A0(\u_uart2wb.tx_data[6] ),
    .A1(\u_uart2wb.u_core.u_txfsm.txdata[6] ),
    .S(_04381_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _09041_ (.A(_04385_),
    .X(_01014_));
 sky130_fd_sc_hd__o21a_1 _09042_ (.A1(\u_uart2wb.reg_rdata[1] ),
    .A2(\u_uart2wb.reg_rdata[2] ),
    .B1(\u_uart2wb.reg_rdata[3] ),
    .X(_04386_));
 sky130_fd_sc_hd__and2_1 _09043_ (.A(_02993_),
    .B(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__nor2_1 _09044_ (.A(_03091_),
    .B(_04386_),
    .Y(_04388_));
 sky130_fd_sc_hd__mux2_1 _09045_ (.A0(_04387_),
    .A1(_04388_),
    .S(\u_uart2wb.reg_rdata[0] ),
    .X(_04389_));
 sky130_fd_sc_hd__a211o_1 _09046_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[56] ),
    .A2(_03167_),
    .B1(_03021_),
    .C1(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__mux2_1 _09047_ (.A0(_04390_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[64] ),
    .S(_03174_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _09048_ (.A(_04391_),
    .X(_01015_));
 sky130_fd_sc_hd__or2b_1 _09049_ (.A(\u_uart2wb.reg_rdata[0] ),
    .B_N(\u_uart2wb.reg_rdata[3] ),
    .X(_04392_));
 sky130_fd_sc_hd__nor2_1 _09050_ (.A(_03629_),
    .B(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__a21o_1 _09051_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[57] ),
    .A2(_03132_),
    .B1(_02939_),
    .X(_04394_));
 sky130_fd_sc_hd__a31o_1 _09052_ (.A1(_03630_),
    .A2(_02959_),
    .A3(_04393_),
    .B1(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__a31o_1 _09053_ (.A1(_03629_),
    .A2(_02960_),
    .A3(_04392_),
    .B1(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__mux2_1 _09054_ (.A0(_04396_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[65] ),
    .S(_03174_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _09055_ (.A(_04397_),
    .X(_01016_));
 sky130_fd_sc_hd__and3b_1 _09056_ (.A_N(_04393_),
    .B(_03038_),
    .C(_03630_),
    .X(_04398_));
 sky130_fd_sc_hd__a211o_1 _09057_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[58] ),
    .A2(_03167_),
    .B1(_03145_),
    .C1(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_2 _09058_ (.A(_02948_),
    .X(_04400_));
 sky130_fd_sc_hd__mux2_1 _09059_ (.A0(_04399_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[66] ),
    .S(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_1 _09060_ (.A(_04401_),
    .X(_01017_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09061_ (.A(_02957_),
    .X(_04402_));
 sky130_fd_sc_hd__and4bb_1 _09062_ (.A_N(_03629_),
    .B_N(_03630_),
    .C(_03071_),
    .D(\u_uart2wb.reg_rdata[3] ),
    .X(_04403_));
 sky130_fd_sc_hd__a211o_1 _09063_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[59] ),
    .A2(_04402_),
    .B1(_02950_),
    .C1(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__mux2_1 _09064_ (.A0(_04404_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[67] ),
    .S(_04400_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _09065_ (.A(_04405_),
    .X(_01018_));
 sky130_fd_sc_hd__a211o_1 _09066_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[60] ),
    .A2(_02971_),
    .B1(_02967_),
    .C1(_04388_),
    .X(_04406_));
 sky130_fd_sc_hd__o21a_1 _09067_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[68] ),
    .A2(_03065_),
    .B1(_04406_),
    .X(_01019_));
 sky130_fd_sc_hd__o2bb2a_1 _09068_ (.A1_N(\u_uart2wb.u_msg.TxMsgBuf[61] ),
    .A2_N(_02982_),
    .B1(_04222_),
    .B2(_02938_),
    .X(_04407_));
 sky130_fd_sc_hd__or3b_1 _09069_ (.A(_03021_),
    .B(_04388_),
    .C_N(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__mux2_1 _09070_ (.A0(_04408_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[69] ),
    .S(_04400_),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_1 _09071_ (.A(_04409_),
    .X(_01020_));
 sky130_fd_sc_hd__a211o_1 _09072_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[62] ),
    .A2(_04402_),
    .B1(_03021_),
    .C1(_04387_),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_1 _09073_ (.A0(_04410_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[70] ),
    .S(_04400_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _09074_ (.A(_04411_),
    .X(_01021_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09075_ (.A(\u_uart2wb.u_msg.TxMsgSize[0] ),
    .X(_04412_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09076_ (.A(_02923_),
    .X(_04413_));
 sky130_fd_sc_hd__nor2_1 _09077_ (.A(_04412_),
    .B(_04215_),
    .Y(_04414_));
 sky130_fd_sc_hd__or4_1 _09078_ (.A(_02947_),
    .B(_02949_),
    .C(_02980_),
    .D(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__o21a_1 _09079_ (.A1(_04412_),
    .A2(_04413_),
    .B1(_04415_),
    .X(_01022_));
 sky130_fd_sc_hd__xnor2_1 _09080_ (.A(\u_uart2wb.u_msg.TxMsgSize[1] ),
    .B(_04412_),
    .Y(_04416_));
 sky130_fd_sc_hd__a211o_1 _09081_ (.A1(_02929_),
    .A2(_04416_),
    .B1(_02973_),
    .C1(_02933_),
    .X(_04417_));
 sky130_fd_sc_hd__o21a_1 _09082_ (.A1(\u_uart2wb.u_msg.TxMsgSize[1] ),
    .A2(_04413_),
    .B1(_04417_),
    .X(_01023_));
 sky130_fd_sc_hd__o21ai_1 _09083_ (.A1(\u_uart2wb.u_msg.TxMsgSize[1] ),
    .A2(_04412_),
    .B1(\u_uart2wb.u_msg.TxMsgSize[2] ),
    .Y(_04418_));
 sky130_fd_sc_hd__a21oi_1 _09084_ (.A1(_02910_),
    .A2(_04418_),
    .B1(_04215_),
    .Y(_04419_));
 sky130_fd_sc_hd__or4_1 _09085_ (.A(_02931_),
    .B(_02979_),
    .C(_02980_),
    .D(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__o21a_1 _09086_ (.A1(\u_uart2wb.u_msg.TxMsgSize[2] ),
    .A2(_04413_),
    .B1(_04420_),
    .X(_01024_));
 sky130_fd_sc_hd__nand2_1 _09087_ (.A(\u_uart2wb.u_msg.TxMsgSize[3] ),
    .B(_02910_),
    .Y(_04421_));
 sky130_fd_sc_hd__a21oi_1 _09088_ (.A1(_02911_),
    .A2(_04421_),
    .B1(_04215_),
    .Y(_04422_));
 sky130_fd_sc_hd__or4_1 _09089_ (.A(_02947_),
    .B(_02979_),
    .C(_02973_),
    .D(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__o21a_1 _09090_ (.A1(\u_uart2wb.u_msg.TxMsgSize[3] ),
    .A2(_04413_),
    .B1(_04423_),
    .X(_01025_));
 sky130_fd_sc_hd__a21o_1 _09091_ (.A1(_02929_),
    .A2(_02911_),
    .B1(_02933_),
    .X(_04424_));
 sky130_fd_sc_hd__a21o_1 _09092_ (.A1(\u_uart2wb.u_msg.TxMsgSize[4] ),
    .A2(_04424_),
    .B1(_04218_),
    .X(_01026_));
 sky130_fd_sc_hd__nor2_1 _09093_ (.A(_02901_),
    .B(_04279_),
    .Y(_04425_));
 sky130_fd_sc_hd__or2_1 _09094_ (.A(_02875_),
    .B(_04279_),
    .X(_04426_));
 sky130_fd_sc_hd__o221a_1 _09095_ (.A1(_02950_),
    .A2(_04425_),
    .B1(_04426_),
    .B2(_03983_),
    .C1(net239),
    .X(_04427_));
 sky130_fd_sc_hd__and3_1 _09096_ (.A(\u_uart2wb.rx_wr ),
    .B(_04274_),
    .C(_04308_),
    .X(_04428_));
 sky130_fd_sc_hd__clkinv_2 _09097_ (.A(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__and3_1 _09098_ (.A(_04312_),
    .B(_04427_),
    .C(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__and3_1 _09099_ (.A(\u_uart2wb.u_msg.RxMsgCnt[0] ),
    .B(_04313_),
    .C(_04430_),
    .X(_04431_));
 sky130_fd_sc_hd__clkbuf_1 _09100_ (.A(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__o211a_1 _09101_ (.A1(_04426_),
    .A2(_04310_),
    .B1(_04430_),
    .C1(_04275_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _09102_ (.A(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__a21oi_1 _09103_ (.A1(_04313_),
    .A2(_04430_),
    .B1(\u_uart2wb.u_msg.RxMsgCnt[0] ),
    .Y(_04435_));
 sky130_fd_sc_hd__nor3_1 _09104_ (.A(_04432_),
    .B(_04434_),
    .C(_04435_),
    .Y(_01027_));
 sky130_fd_sc_hd__clkbuf_1 _09105_ (.A(\u_uart2wb.u_msg.RxMsgCnt[1] ),
    .X(_04436_));
 sky130_fd_sc_hd__a21oi_1 _09106_ (.A1(_04436_),
    .A2(_04432_),
    .B1(_04434_),
    .Y(_04437_));
 sky130_fd_sc_hd__o21a_1 _09107_ (.A1(_04436_),
    .A2(_04432_),
    .B1(_04437_),
    .X(_01028_));
 sky130_fd_sc_hd__and3_1 _09108_ (.A(\u_uart2wb.u_msg.RxMsgCnt[2] ),
    .B(_04436_),
    .C(_04431_),
    .X(_04438_));
 sky130_fd_sc_hd__nor2_1 _09109_ (.A(_04426_),
    .B(_04310_),
    .Y(_04439_));
 sky130_fd_sc_hd__or2_1 _09110_ (.A(_04307_),
    .B(_04439_),
    .X(_04440_));
 sky130_fd_sc_hd__a31o_1 _09111_ (.A1(_04436_),
    .A2(_04432_),
    .A3(_04440_),
    .B1(\u_uart2wb.u_msg.RxMsgCnt[2] ),
    .X(_04441_));
 sky130_fd_sc_hd__nor3b_1 _09112_ (.A(_04434_),
    .B(_04438_),
    .C_N(_04441_),
    .Y(_01029_));
 sky130_fd_sc_hd__and2_1 _09113_ (.A(\u_uart2wb.u_msg.RxMsgCnt[3] ),
    .B(_04438_),
    .X(_04442_));
 sky130_fd_sc_hd__nor2_1 _09114_ (.A(_04433_),
    .B(_04442_),
    .Y(_04443_));
 sky130_fd_sc_hd__o21a_1 _09115_ (.A1(\u_uart2wb.u_msg.RxMsgCnt[3] ),
    .A2(_04438_),
    .B1(_04443_),
    .X(_01030_));
 sky130_fd_sc_hd__a21oi_1 _09116_ (.A1(\u_uart2wb.u_msg.RxMsgCnt[4] ),
    .A2(_04442_),
    .B1(_04434_),
    .Y(_04444_));
 sky130_fd_sc_hd__o21a_1 _09117_ (.A1(\u_uart2wb.u_msg.RxMsgCnt[4] ),
    .A2(_04442_),
    .B1(_04444_),
    .X(_01031_));
 sky130_fd_sc_hd__inv_2 _09118_ (.A(_04282_),
    .Y(_04445_));
 sky130_fd_sc_hd__nor3_1 _09119_ (.A(\u_uart2wb.u_msg.cmd[8] ),
    .B(\u_uart2wb.u_msg.cmd[10] ),
    .C(_04294_),
    .Y(_04446_));
 sky130_fd_sc_hd__a22o_1 _09120_ (.A1(_04445_),
    .A2(_04446_),
    .B1(_04296_),
    .B2(_04292_),
    .X(_04447_));
 sky130_fd_sc_hd__a21oi_1 _09121_ (.A1(_04291_),
    .A2(_04447_),
    .B1(_04275_),
    .Y(_04448_));
 sky130_fd_sc_hd__a31o_1 _09122_ (.A1(_02876_),
    .A2(_02891_),
    .A3(_02904_),
    .B1(_02926_),
    .X(_04449_));
 sky130_fd_sc_hd__nor2_1 _09123_ (.A(_02908_),
    .B(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__a221o_1 _09124_ (.A1(\u_uart2wb.u_msg.NextState[0] ),
    .A2(_03132_),
    .B1(_04445_),
    .B2(_04309_),
    .C1(_04261_),
    .X(_04451_));
 sky130_fd_sc_hd__or4_1 _09125_ (.A(_04311_),
    .B(_04448_),
    .C(_04450_),
    .D(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__a21boi_2 _09126_ (.A1(_01158_),
    .A2(_02874_),
    .B1_N(_02880_),
    .Y(_04453_));
 sky130_fd_sc_hd__a211o_1 _09127_ (.A1(_04278_),
    .A2(_04309_),
    .B1(_04375_),
    .C1(_04298_),
    .X(_04454_));
 sky130_fd_sc_hd__or4_1 _09128_ (.A(_04281_),
    .B(_04428_),
    .C(_04453_),
    .D(_04454_),
    .X(_04455_));
 sky130_fd_sc_hd__nor2_2 _09129_ (.A(_04300_),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__mux2_1 _09130_ (.A0(_02902_),
    .A1(_04452_),
    .S(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__clkbuf_1 _09131_ (.A(_04457_),
    .X(_01032_));
 sky130_fd_sc_hd__a211o_1 _09132_ (.A1(\u_uart2wb.u_msg.NextState[1] ),
    .A2(_03072_),
    .B1(_02908_),
    .C1(_04262_),
    .X(_04458_));
 sky130_fd_sc_hd__a31o_1 _09133_ (.A1(_04307_),
    .A2(_04349_),
    .A3(_04350_),
    .B1(_04458_),
    .X(_04459_));
 sky130_fd_sc_hd__mux2_1 _09134_ (.A0(_02901_),
    .A1(_04459_),
    .S(_04456_),
    .X(_04460_));
 sky130_fd_sc_hd__clkbuf_1 _09135_ (.A(_04460_),
    .X(_01033_));
 sky130_fd_sc_hd__or2_1 _09136_ (.A(_04349_),
    .B(_04439_),
    .X(_04461_));
 sky130_fd_sc_hd__a311o_1 _09137_ (.A1(_04313_),
    .A2(_04440_),
    .A3(_04461_),
    .B1(_04455_),
    .C1(_04300_),
    .X(_04462_));
 sky130_fd_sc_hd__o21a_1 _09138_ (.A1(_04446_),
    .A2(_04296_),
    .B1(_04311_),
    .X(_04463_));
 sky130_fd_sc_hd__a211o_1 _09139_ (.A1(\u_uart2wb.u_msg.NextState[2] ),
    .A2(_03139_),
    .B1(_04262_),
    .C1(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__a22o_1 _09140_ (.A1(_02954_),
    .A2(_04462_),
    .B1(_04464_),
    .B2(_04456_),
    .X(_01034_));
 sky130_fd_sc_hd__a21o_1 _09141_ (.A1(\u_uart2wb.u_msg.NextState[3] ),
    .A2(_02927_),
    .B1(_02908_),
    .X(_04465_));
 sky130_fd_sc_hd__a31o_1 _09142_ (.A1(_04291_),
    .A2(_04307_),
    .A3(_04289_),
    .B1(_04465_),
    .X(_04466_));
 sky130_fd_sc_hd__mux2_1 _09143_ (.A0(_02877_),
    .A1(_04466_),
    .S(_04456_),
    .X(_04467_));
 sky130_fd_sc_hd__clkbuf_1 _09144_ (.A(_04467_),
    .X(_01035_));
 sky130_fd_sc_hd__o21ai_1 _09145_ (.A1(_02900_),
    .A2(_02907_),
    .B1(_02902_),
    .Y(_04468_));
 sky130_fd_sc_hd__nor3_2 _09146_ (.A(_02880_),
    .B(_02917_),
    .C(_04449_),
    .Y(_04469_));
 sky130_fd_sc_hd__mux2_1 _09147_ (.A0(\u_uart2wb.u_msg.NextState[0] ),
    .A1(_04468_),
    .S(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__clkbuf_1 _09148_ (.A(_04470_),
    .X(_01036_));
 sky130_fd_sc_hd__inv_2 _09149_ (.A(\u_uart2wb.u_msg.NextState[1] ),
    .Y(_04471_));
 sky130_fd_sc_hd__o21ai_1 _09150_ (.A1(_04471_),
    .A2(_04469_),
    .B1(_04196_),
    .Y(_01037_));
 sky130_fd_sc_hd__mux2_1 _09151_ (.A0(\u_uart2wb.u_msg.NextState[2] ),
    .A1(_02907_),
    .S(_04469_),
    .X(_04472_));
 sky130_fd_sc_hd__clkbuf_1 _09152_ (.A(_04472_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _09153_ (.A0(\u_uart2wb.u_msg.NextState[3] ),
    .A1(_03145_),
    .S(_04469_),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_1 _09154_ (.A(_04473_),
    .X(_01039_));
 sky130_fd_sc_hd__and4_1 _09155_ (.A(net237),
    .B(_03984_),
    .C(_04269_),
    .D(_04309_),
    .X(_04474_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09156_ (.A(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__mux2_1 _09157_ (.A0(\u_uart2wb.u_msg.cmd[0] ),
    .A1(_04002_),
    .S(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__clkbuf_1 _09158_ (.A(_04476_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _09159_ (.A0(\u_uart2wb.u_msg.cmd[1] ),
    .A1(_04007_),
    .S(_04475_),
    .X(_04477_));
 sky130_fd_sc_hd__clkbuf_1 _09160_ (.A(_04477_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _09161_ (.A0(\u_uart2wb.u_msg.cmd[2] ),
    .A1(_04011_),
    .S(_04475_),
    .X(_04478_));
 sky130_fd_sc_hd__clkbuf_1 _09162_ (.A(_04478_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _09163_ (.A0(\u_uart2wb.u_msg.cmd[3] ),
    .A1(_04015_),
    .S(_04475_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _09164_ (.A(_04479_),
    .X(_01043_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09165_ (.A(_04474_),
    .X(_04480_));
 sky130_fd_sc_hd__mux2_1 _09166_ (.A0(\u_uart2wb.u_msg.cmd[4] ),
    .A1(_04019_),
    .S(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__clkbuf_1 _09167_ (.A(_04481_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _09168_ (.A0(\u_uart2wb.u_msg.cmd[5] ),
    .A1(_04023_),
    .S(_04480_),
    .X(_04482_));
 sky130_fd_sc_hd__clkbuf_1 _09169_ (.A(_04482_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(\u_uart2wb.u_msg.cmd[6] ),
    .A1(_04026_),
    .S(_04480_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_1 _09171_ (.A(_04483_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _09172_ (.A0(\u_uart2wb.u_msg.cmd[7] ),
    .A1(_04029_),
    .S(_04480_),
    .X(_04484_));
 sky130_fd_sc_hd__clkbuf_1 _09173_ (.A(_04484_),
    .X(_01047_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09174_ (.A(_04474_),
    .X(_04485_));
 sky130_fd_sc_hd__mux2_1 _09175_ (.A0(\u_uart2wb.u_msg.cmd[8] ),
    .A1(\u_uart2wb.u_msg.cmd[0] ),
    .S(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__clkbuf_1 _09176_ (.A(_04486_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _09177_ (.A0(\u_uart2wb.u_msg.cmd[9] ),
    .A1(\u_uart2wb.u_msg.cmd[1] ),
    .S(_04485_),
    .X(_04487_));
 sky130_fd_sc_hd__clkbuf_1 _09178_ (.A(_04487_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _09179_ (.A0(\u_uart2wb.u_msg.cmd[10] ),
    .A1(\u_uart2wb.u_msg.cmd[2] ),
    .S(_04485_),
    .X(_04488_));
 sky130_fd_sc_hd__clkbuf_1 _09180_ (.A(_04488_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _09181_ (.A0(\u_uart2wb.u_msg.cmd[11] ),
    .A1(\u_uart2wb.u_msg.cmd[3] ),
    .S(_04485_),
    .X(_04489_));
 sky130_fd_sc_hd__clkbuf_1 _09182_ (.A(_04489_),
    .X(_01051_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09183_ (.A(_04474_),
    .X(_04490_));
 sky130_fd_sc_hd__mux2_1 _09184_ (.A0(\u_uart2wb.u_msg.cmd[12] ),
    .A1(\u_uart2wb.u_msg.cmd[4] ),
    .S(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _09185_ (.A(_04491_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _09186_ (.A0(\u_uart2wb.u_msg.cmd[13] ),
    .A1(\u_uart2wb.u_msg.cmd[5] ),
    .S(_04490_),
    .X(_04492_));
 sky130_fd_sc_hd__clkbuf_1 _09187_ (.A(_04492_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _09188_ (.A0(\u_uart2wb.u_msg.cmd[14] ),
    .A1(\u_uart2wb.u_msg.cmd[6] ),
    .S(_04490_),
    .X(_04493_));
 sky130_fd_sc_hd__clkbuf_1 _09189_ (.A(_04493_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(\u_uart2wb.u_msg.cmd[15] ),
    .A1(\u_uart2wb.u_msg.cmd[7] ),
    .S(_04490_),
    .X(_04494_));
 sky130_fd_sc_hd__clkbuf_1 _09191_ (.A(_04494_),
    .X(_01055_));
 sky130_fd_sc_hd__nand2_1 _09192_ (.A(net249),
    .B(_02927_),
    .Y(_04495_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09193_ (.A(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[120] ),
    .A1(\u_uart2wb.tx_data[0] ),
    .S(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__clkbuf_1 _09195_ (.A(_04497_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[121] ),
    .A1(\u_uart2wb.tx_data[1] ),
    .S(_04496_),
    .X(_04498_));
 sky130_fd_sc_hd__clkbuf_1 _09197_ (.A(_04498_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[122] ),
    .A1(\u_uart2wb.tx_data[2] ),
    .S(_04496_),
    .X(_04499_));
 sky130_fd_sc_hd__clkbuf_1 _09199_ (.A(_04499_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[123] ),
    .A1(\u_uart2wb.tx_data[3] ),
    .S(_04496_),
    .X(_04500_));
 sky130_fd_sc_hd__clkbuf_1 _09201_ (.A(_04500_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _09202_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[124] ),
    .A1(\u_uart2wb.tx_data[4] ),
    .S(_04495_),
    .X(_04501_));
 sky130_fd_sc_hd__clkbuf_1 _09203_ (.A(_04501_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _09204_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[125] ),
    .A1(\u_uart2wb.tx_data[5] ),
    .S(_04495_),
    .X(_04502_));
 sky130_fd_sc_hd__clkbuf_1 _09205_ (.A(_04502_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _09206_ (.A0(\u_uart2wb.u_msg.TxMsgBuf[126] ),
    .A1(\u_uart2wb.tx_data[6] ),
    .S(_04495_),
    .X(_04503_));
 sky130_fd_sc_hd__clkbuf_1 _09207_ (.A(_04503_),
    .X(_01062_));
 sky130_fd_sc_hd__o21a_1 _09208_ (.A1(\u_uart2wb.reg_rdata[13] ),
    .A2(\u_uart2wb.reg_rdata[14] ),
    .B1(\u_uart2wb.reg_rdata[15] ),
    .X(_04504_));
 sky130_fd_sc_hd__nor2_1 _09209_ (.A(_03091_),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__inv_2 _09210_ (.A(\u_uart2wb.reg_rdata[12] ),
    .Y(_04506_));
 sky130_fd_sc_hd__a32o_1 _09211_ (.A1(_04506_),
    .A2(_03045_),
    .A3(_04504_),
    .B1(_02952_),
    .B2(\u_uart2wb.u_msg.TxMsgBuf[80] ),
    .X(_04507_));
 sky130_fd_sc_hd__a211o_1 _09212_ (.A1(\u_uart2wb.reg_rdata[12] ),
    .A2(_04505_),
    .B1(_04507_),
    .C1(_02996_),
    .X(_04508_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09213_ (.A(_02948_),
    .X(_04509_));
 sky130_fd_sc_hd__mux2_1 _09214_ (.A0(_04508_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[88] ),
    .S(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_1 _09215_ (.A(_04510_),
    .X(_01063_));
 sky130_fd_sc_hd__nand2_1 _09216_ (.A(_04506_),
    .B(\u_uart2wb.reg_rdata[15] ),
    .Y(_04511_));
 sky130_fd_sc_hd__a32o_1 _09217_ (.A1(_03638_),
    .A2(_03071_),
    .A3(_04511_),
    .B1(\u_uart2wb.u_msg.TxMsgBuf[81] ),
    .B2(_02982_),
    .X(_04512_));
 sky130_fd_sc_hd__inv_2 _09218_ (.A(\u_uart2wb.reg_rdata[14] ),
    .Y(_04513_));
 sky130_fd_sc_hd__or4_1 _09219_ (.A(\u_uart2wb.reg_rdata[13] ),
    .B(_04513_),
    .C(_03024_),
    .D(_04511_),
    .X(_04514_));
 sky130_fd_sc_hd__or3b_1 _09220_ (.A(_03020_),
    .B(_04512_),
    .C_N(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__mux2_1 _09221_ (.A0(_04515_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[89] ),
    .S(_04509_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_1 _09222_ (.A(_04516_),
    .X(_01064_));
 sky130_fd_sc_hd__o211a_1 _09223_ (.A1(_03638_),
    .A2(_04511_),
    .B1(_02959_),
    .C1(\u_uart2wb.reg_rdata[14] ),
    .X(_04517_));
 sky130_fd_sc_hd__a211o_1 _09224_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[82] ),
    .A2(_04402_),
    .B1(_03145_),
    .C1(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__mux2_1 _09225_ (.A0(_04518_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[90] ),
    .S(_04509_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _09226_ (.A(_04519_),
    .X(_01065_));
 sky130_fd_sc_hd__and4b_1 _09227_ (.A_N(_03638_),
    .B(_04513_),
    .C(_03045_),
    .D(\u_uart2wb.reg_rdata[15] ),
    .X(_04520_));
 sky130_fd_sc_hd__a211o_1 _09228_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[83] ),
    .A2(_04402_),
    .B1(_02962_),
    .C1(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__mux2_1 _09229_ (.A0(_04521_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[91] ),
    .S(_04509_),
    .X(_04522_));
 sky130_fd_sc_hd__clkbuf_1 _09230_ (.A(_04522_),
    .X(_01066_));
 sky130_fd_sc_hd__a211o_1 _09231_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[84] ),
    .A2(_03138_),
    .B1(_02930_),
    .C1(_04505_),
    .X(_04523_));
 sky130_fd_sc_hd__mux2_1 _09232_ (.A0(_04523_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[92] ),
    .S(_02992_),
    .X(_04524_));
 sky130_fd_sc_hd__clkbuf_1 _09233_ (.A(_04524_),
    .X(_01067_));
 sky130_fd_sc_hd__a211o_1 _09234_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[85] ),
    .A2(_03138_),
    .B1(_02995_),
    .C1(_04505_),
    .X(_04525_));
 sky130_fd_sc_hd__mux2_1 _09235_ (.A0(_04525_),
    .A1(\u_uart2wb.u_msg.TxMsgBuf[93] ),
    .S(_02992_),
    .X(_04526_));
 sky130_fd_sc_hd__clkbuf_1 _09236_ (.A(_04526_),
    .X(_01068_));
 sky130_fd_sc_hd__a22o_1 _09237_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[86] ),
    .A2(_02983_),
    .B1(_03067_),
    .B2(_04504_),
    .X(_04527_));
 sky130_fd_sc_hd__or3_1 _09238_ (.A(_02949_),
    .B(_02996_),
    .C(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__o21a_1 _09239_ (.A1(\u_uart2wb.u_msg.TxMsgBuf[94] ),
    .A2(_02924_),
    .B1(_04528_),
    .X(_01069_));
 sky130_fd_sc_hd__and3b_1 _09240_ (.A_N(\u_spi2wb.u_if.sck_l1 ),
    .B(\u_spi2wb.u_if.sck_l2 ),
    .C(\u_spi2wb.u_if.rd_phase ),
    .X(_04529_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09241_ (.A(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__mux2_1 _09242_ (.A0(net71),
    .A1(\u_spi2wb.u_if.RegSdOut[31] ),
    .S(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__clkbuf_1 _09243_ (.A(_04531_),
    .X(_01070_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09244_ (.A(_01836_),
    .X(_04532_));
 sky130_fd_sc_hd__nor2_1 _09245_ (.A(_04532_),
    .B(_04530_),
    .Y(_04533_));
 sky130_fd_sc_hd__a22o_1 _09246_ (.A1(\wb_dat_o[0] ),
    .A2(_04532_),
    .B1(_04533_),
    .B2(\u_spi2wb.u_if.RegSdOut[0] ),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _09247_ (.A0(\u_spi2wb.u_if.RegSdOut[1] ),
    .A1(\u_spi2wb.u_if.RegSdOut[0] ),
    .S(_04530_),
    .X(_04534_));
 sky130_fd_sc_hd__mux2_1 _09248_ (.A0(_04534_),
    .A1(\wb_dat_o[1] ),
    .S(_04532_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_1 _09249_ (.A(_04535_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _09250_ (.A0(\u_spi2wb.u_if.RegSdOut[2] ),
    .A1(\u_spi2wb.u_if.RegSdOut[1] ),
    .S(_04530_),
    .X(_04536_));
 sky130_fd_sc_hd__mux2_1 _09251_ (.A0(_04536_),
    .A1(\wb_dat_o[2] ),
    .S(_04532_),
    .X(_04537_));
 sky130_fd_sc_hd__clkbuf_1 _09252_ (.A(_04537_),
    .X(_01073_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09253_ (.A(_04529_),
    .X(_04538_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09254_ (.A(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__mux2_1 _09255_ (.A0(\u_spi2wb.u_if.RegSdOut[3] ),
    .A1(\u_spi2wb.u_if.RegSdOut[2] ),
    .S(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09256_ (.A(_01837_),
    .X(_04541_));
 sky130_fd_sc_hd__mux2_1 _09257_ (.A0(_04540_),
    .A1(\wb_dat_o[3] ),
    .S(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__clkbuf_1 _09258_ (.A(_04542_),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _09259_ (.A0(\u_spi2wb.u_if.RegSdOut[4] ),
    .A1(\u_spi2wb.u_if.RegSdOut[3] ),
    .S(_04539_),
    .X(_04543_));
 sky130_fd_sc_hd__mux2_1 _09260_ (.A0(_04543_),
    .A1(\wb_dat_o[4] ),
    .S(_04541_),
    .X(_04544_));
 sky130_fd_sc_hd__clkbuf_1 _09261_ (.A(_04544_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _09262_ (.A0(\u_spi2wb.u_if.RegSdOut[5] ),
    .A1(\u_spi2wb.u_if.RegSdOut[4] ),
    .S(_04539_),
    .X(_04545_));
 sky130_fd_sc_hd__mux2_1 _09263_ (.A0(_04545_),
    .A1(\wb_dat_o[5] ),
    .S(_04541_),
    .X(_04546_));
 sky130_fd_sc_hd__clkbuf_1 _09264_ (.A(_04546_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _09265_ (.A0(\u_spi2wb.u_if.RegSdOut[6] ),
    .A1(\u_spi2wb.u_if.RegSdOut[5] ),
    .S(_04539_),
    .X(_04547_));
 sky130_fd_sc_hd__mux2_1 _09266_ (.A0(_04547_),
    .A1(\wb_dat_o[6] ),
    .S(_04541_),
    .X(_04548_));
 sky130_fd_sc_hd__clkbuf_1 _09267_ (.A(_04548_),
    .X(_01077_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09268_ (.A(_04538_),
    .X(_04549_));
 sky130_fd_sc_hd__mux2_1 _09269_ (.A0(\u_spi2wb.u_if.RegSdOut[7] ),
    .A1(\u_spi2wb.u_if.RegSdOut[6] ),
    .S(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09270_ (.A(_01837_),
    .X(_04551_));
 sky130_fd_sc_hd__mux2_1 _09271_ (.A0(_04550_),
    .A1(\wb_dat_o[7] ),
    .S(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__clkbuf_1 _09272_ (.A(_04552_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _09273_ (.A0(\u_spi2wb.u_if.RegSdOut[8] ),
    .A1(\u_spi2wb.u_if.RegSdOut[7] ),
    .S(_04549_),
    .X(_04553_));
 sky130_fd_sc_hd__mux2_1 _09274_ (.A0(_04553_),
    .A1(\wb_dat_o[8] ),
    .S(_04551_),
    .X(_04554_));
 sky130_fd_sc_hd__clkbuf_1 _09275_ (.A(_04554_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _09276_ (.A0(\u_spi2wb.u_if.RegSdOut[9] ),
    .A1(\u_spi2wb.u_if.RegSdOut[8] ),
    .S(_04549_),
    .X(_04555_));
 sky130_fd_sc_hd__mux2_1 _09277_ (.A0(_04555_),
    .A1(\wb_dat_o[9] ),
    .S(_04551_),
    .X(_04556_));
 sky130_fd_sc_hd__clkbuf_1 _09278_ (.A(_04556_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _09279_ (.A0(\u_spi2wb.u_if.RegSdOut[10] ),
    .A1(\u_spi2wb.u_if.RegSdOut[9] ),
    .S(_04549_),
    .X(_04557_));
 sky130_fd_sc_hd__mux2_1 _09280_ (.A0(_04557_),
    .A1(\wb_dat_o[10] ),
    .S(_04551_),
    .X(_04558_));
 sky130_fd_sc_hd__clkbuf_1 _09281_ (.A(_04558_),
    .X(_01081_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09282_ (.A(_04538_),
    .X(_04559_));
 sky130_fd_sc_hd__mux2_1 _09283_ (.A0(\u_spi2wb.u_if.RegSdOut[11] ),
    .A1(\u_spi2wb.u_if.RegSdOut[10] ),
    .S(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_1 _09284_ (.A(_01836_),
    .X(_04561_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09285_ (.A(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__mux2_1 _09286_ (.A0(_04560_),
    .A1(\wb_dat_o[11] ),
    .S(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__clkbuf_1 _09287_ (.A(_04563_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _09288_ (.A0(\u_spi2wb.u_if.RegSdOut[12] ),
    .A1(\u_spi2wb.u_if.RegSdOut[11] ),
    .S(_04559_),
    .X(_04564_));
 sky130_fd_sc_hd__mux2_1 _09289_ (.A0(_04564_),
    .A1(\wb_dat_o[12] ),
    .S(_04562_),
    .X(_04565_));
 sky130_fd_sc_hd__clkbuf_1 _09290_ (.A(_04565_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _09291_ (.A0(\u_spi2wb.u_if.RegSdOut[13] ),
    .A1(\u_spi2wb.u_if.RegSdOut[12] ),
    .S(_04559_),
    .X(_04566_));
 sky130_fd_sc_hd__mux2_1 _09292_ (.A0(_04566_),
    .A1(\wb_dat_o[13] ),
    .S(_04562_),
    .X(_04567_));
 sky130_fd_sc_hd__clkbuf_1 _09293_ (.A(_04567_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _09294_ (.A0(\u_spi2wb.u_if.RegSdOut[14] ),
    .A1(\u_spi2wb.u_if.RegSdOut[13] ),
    .S(_04559_),
    .X(_04568_));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(_04568_),
    .A1(\wb_dat_o[14] ),
    .S(_04562_),
    .X(_04569_));
 sky130_fd_sc_hd__clkbuf_1 _09296_ (.A(_04569_),
    .X(_01085_));
 sky130_fd_sc_hd__clkbuf_1 _09297_ (.A(_04529_),
    .X(_04570_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09298_ (.A(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(\u_spi2wb.u_if.RegSdOut[15] ),
    .A1(\u_spi2wb.u_if.RegSdOut[14] ),
    .S(_04571_),
    .X(_04572_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09300_ (.A(_04561_),
    .X(_04573_));
 sky130_fd_sc_hd__mux2_1 _09301_ (.A0(_04572_),
    .A1(\wb_dat_o[15] ),
    .S(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__clkbuf_1 _09302_ (.A(_04574_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _09303_ (.A0(\u_spi2wb.u_if.RegSdOut[16] ),
    .A1(\u_spi2wb.u_if.RegSdOut[15] ),
    .S(_04571_),
    .X(_04575_));
 sky130_fd_sc_hd__mux2_1 _09304_ (.A0(_04575_),
    .A1(\wb_dat_o[16] ),
    .S(_04573_),
    .X(_04576_));
 sky130_fd_sc_hd__clkbuf_1 _09305_ (.A(_04576_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _09306_ (.A0(\u_spi2wb.u_if.RegSdOut[17] ),
    .A1(\u_spi2wb.u_if.RegSdOut[16] ),
    .S(_04571_),
    .X(_04577_));
 sky130_fd_sc_hd__mux2_1 _09307_ (.A0(_04577_),
    .A1(\wb_dat_o[17] ),
    .S(_04573_),
    .X(_04578_));
 sky130_fd_sc_hd__clkbuf_1 _09308_ (.A(_04578_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _09309_ (.A0(\u_spi2wb.u_if.RegSdOut[18] ),
    .A1(\u_spi2wb.u_if.RegSdOut[17] ),
    .S(_04571_),
    .X(_04579_));
 sky130_fd_sc_hd__mux2_1 _09310_ (.A0(_04579_),
    .A1(\wb_dat_o[18] ),
    .S(_04573_),
    .X(_04580_));
 sky130_fd_sc_hd__clkbuf_1 _09311_ (.A(_04580_),
    .X(_01089_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09312_ (.A(_04570_),
    .X(_04581_));
 sky130_fd_sc_hd__mux2_1 _09313_ (.A0(\u_spi2wb.u_if.RegSdOut[19] ),
    .A1(\u_spi2wb.u_if.RegSdOut[18] ),
    .S(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09314_ (.A(_04561_),
    .X(_04583_));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(_04582_),
    .A1(\wb_dat_o[19] ),
    .S(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__clkbuf_1 _09316_ (.A(_04584_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(\u_spi2wb.u_if.RegSdOut[20] ),
    .A1(\u_spi2wb.u_if.RegSdOut[19] ),
    .S(_04581_),
    .X(_04585_));
 sky130_fd_sc_hd__mux2_1 _09318_ (.A0(_04585_),
    .A1(\wb_dat_o[20] ),
    .S(_04583_),
    .X(_04586_));
 sky130_fd_sc_hd__clkbuf_1 _09319_ (.A(_04586_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _09320_ (.A0(\u_spi2wb.u_if.RegSdOut[21] ),
    .A1(\u_spi2wb.u_if.RegSdOut[20] ),
    .S(_04581_),
    .X(_04587_));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(_04587_),
    .A1(\wb_dat_o[21] ),
    .S(_04583_),
    .X(_04588_));
 sky130_fd_sc_hd__clkbuf_1 _09322_ (.A(_04588_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(\u_spi2wb.u_if.RegSdOut[22] ),
    .A1(\u_spi2wb.u_if.RegSdOut[21] ),
    .S(_04581_),
    .X(_04589_));
 sky130_fd_sc_hd__mux2_1 _09324_ (.A0(_04589_),
    .A1(\wb_dat_o[22] ),
    .S(_04583_),
    .X(_04590_));
 sky130_fd_sc_hd__clkbuf_1 _09325_ (.A(_04590_),
    .X(_01093_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09326_ (.A(_04570_),
    .X(_04591_));
 sky130_fd_sc_hd__mux2_1 _09327_ (.A0(\u_spi2wb.u_if.RegSdOut[23] ),
    .A1(\u_spi2wb.u_if.RegSdOut[22] ),
    .S(_04591_),
    .X(_04592_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09328_ (.A(_04561_),
    .X(_04593_));
 sky130_fd_sc_hd__mux2_1 _09329_ (.A0(_04592_),
    .A1(\wb_dat_o[23] ),
    .S(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__clkbuf_1 _09330_ (.A(_04594_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _09331_ (.A0(\u_spi2wb.u_if.RegSdOut[24] ),
    .A1(\u_spi2wb.u_if.RegSdOut[23] ),
    .S(_04591_),
    .X(_04595_));
 sky130_fd_sc_hd__mux2_1 _09332_ (.A0(_04595_),
    .A1(\wb_dat_o[24] ),
    .S(_04593_),
    .X(_04596_));
 sky130_fd_sc_hd__clkbuf_1 _09333_ (.A(_04596_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _09334_ (.A0(\u_spi2wb.u_if.RegSdOut[25] ),
    .A1(\u_spi2wb.u_if.RegSdOut[24] ),
    .S(_04591_),
    .X(_04597_));
 sky130_fd_sc_hd__mux2_1 _09335_ (.A0(_04597_),
    .A1(\wb_dat_o[25] ),
    .S(_04593_),
    .X(_04598_));
 sky130_fd_sc_hd__clkbuf_1 _09336_ (.A(_04598_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _09337_ (.A0(\u_spi2wb.u_if.RegSdOut[26] ),
    .A1(\u_spi2wb.u_if.RegSdOut[25] ),
    .S(_04591_),
    .X(_04599_));
 sky130_fd_sc_hd__mux2_1 _09338_ (.A0(_04599_),
    .A1(\wb_dat_o[26] ),
    .S(_04593_),
    .X(_04600_));
 sky130_fd_sc_hd__clkbuf_1 _09339_ (.A(_04600_),
    .X(_01097_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09340_ (.A(_04570_),
    .X(_04601_));
 sky130_fd_sc_hd__mux2_1 _09341_ (.A0(\u_spi2wb.u_if.RegSdOut[27] ),
    .A1(\u_spi2wb.u_if.RegSdOut[26] ),
    .S(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09342_ (.A(_01836_),
    .X(_04603_));
 sky130_fd_sc_hd__mux2_1 _09343_ (.A0(_04602_),
    .A1(\wb_dat_o[27] ),
    .S(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__clkbuf_1 _09344_ (.A(_04604_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _09345_ (.A0(\u_spi2wb.u_if.RegSdOut[28] ),
    .A1(\u_spi2wb.u_if.RegSdOut[27] ),
    .S(_04601_),
    .X(_04605_));
 sky130_fd_sc_hd__mux2_1 _09346_ (.A0(_04605_),
    .A1(\wb_dat_o[28] ),
    .S(_04603_),
    .X(_04606_));
 sky130_fd_sc_hd__clkbuf_1 _09347_ (.A(_04606_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _09348_ (.A0(\u_spi2wb.u_if.RegSdOut[29] ),
    .A1(\u_spi2wb.u_if.RegSdOut[28] ),
    .S(_04601_),
    .X(_04607_));
 sky130_fd_sc_hd__mux2_1 _09349_ (.A0(_04607_),
    .A1(\wb_dat_o[29] ),
    .S(_04603_),
    .X(_04608_));
 sky130_fd_sc_hd__clkbuf_1 _09350_ (.A(_04608_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _09351_ (.A0(\u_spi2wb.u_if.RegSdOut[30] ),
    .A1(\u_spi2wb.u_if.RegSdOut[29] ),
    .S(_04601_),
    .X(_04609_));
 sky130_fd_sc_hd__mux2_1 _09352_ (.A0(_04609_),
    .A1(\wb_dat_o[30] ),
    .S(_04603_),
    .X(_04610_));
 sky130_fd_sc_hd__clkbuf_1 _09353_ (.A(_04610_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _09354_ (.A0(\u_spi2wb.u_if.RegSdOut[31] ),
    .A1(\u_spi2wb.u_if.RegSdOut[30] ),
    .S(_04538_),
    .X(_04611_));
 sky130_fd_sc_hd__mux2_1 _09355_ (.A0(_04611_),
    .A1(\wb_dat_o[31] ),
    .S(_01837_),
    .X(_04612_));
 sky130_fd_sc_hd__clkbuf_1 _09356_ (.A(_04612_),
    .X(_01102_));
 sky130_fd_sc_hd__o41a_1 _09357_ (.A1(_01122_),
    .A2(\u_spi2wb.u_if.spi_if_st[0] ),
    .A3(_01120_),
    .A4(_01450_),
    .B1(_01460_),
    .X(_04613_));
 sky130_fd_sc_hd__o21ai_1 _09358_ (.A1(\u_spi2wb.u_if.ssn_l1 ),
    .A2(_04613_),
    .B1(_01454_),
    .Y(_04614_));
 sky130_fd_sc_hd__mux2_1 _09359_ (.A0(_01452_),
    .A1(net72),
    .S(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__clkbuf_1 _09360_ (.A(_04615_),
    .X(_01103_));
 sky130_fd_sc_hd__or2b_1 _09361_ (.A(_01835_),
    .B_N(_01112_),
    .X(_04616_));
 sky130_fd_sc_hd__o31a_1 _09362_ (.A1(_01111_),
    .A2(_01112_),
    .A3(_03598_),
    .B1(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__nor2_1 _09363_ (.A(_01459_),
    .B(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__o21a_1 _09364_ (.A1(_01457_),
    .A2(_04618_),
    .B1(\u_spi2wb.reg_wr ),
    .X(_04619_));
 sky130_fd_sc_hd__a21o_1 _09365_ (.A1(_01449_),
    .A2(_04617_),
    .B1(_04619_),
    .X(_01104_));
 sky130_fd_sc_hd__dfrtp_4 _09366_ (.CLK(clknet_leaf_74_wbm_clk_i),
    .D(_00038_),
    .RESET_B(net270),
    .Q(\u_spi2wb.reg_rd ));
 sky130_fd_sc_hd__dfrtp_4 _09367_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_00039_),
    .RESET_B(net294),
    .Q(\wb_dat_o[0] ));
 sky130_fd_sc_hd__dfrtp_4 _09368_ (.CLK(clknet_leaf_89_wbm_clk_i),
    .D(_00040_),
    .RESET_B(net294),
    .Q(\wb_dat_o[1] ));
 sky130_fd_sc_hd__dfrtp_4 _09369_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00041_),
    .RESET_B(net292),
    .Q(\wb_dat_o[2] ));
 sky130_fd_sc_hd__dfrtp_4 _09370_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00042_),
    .RESET_B(net292),
    .Q(\wb_dat_o[3] ));
 sky130_fd_sc_hd__dfrtp_4 _09371_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00043_),
    .RESET_B(net292),
    .Q(\wb_dat_o[4] ));
 sky130_fd_sc_hd__dfrtp_4 _09372_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00044_),
    .RESET_B(net292),
    .Q(\wb_dat_o[5] ));
 sky130_fd_sc_hd__dfrtp_4 _09373_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_00045_),
    .RESET_B(net292),
    .Q(\wb_dat_o[6] ));
 sky130_fd_sc_hd__dfrtp_4 _09374_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00046_),
    .RESET_B(net292),
    .Q(\wb_dat_o[7] ));
 sky130_fd_sc_hd__dfrtp_4 _09375_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00047_),
    .RESET_B(net292),
    .Q(\wb_dat_o[8] ));
 sky130_fd_sc_hd__dfrtp_4 _09376_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00048_),
    .RESET_B(net292),
    .Q(\wb_dat_o[9] ));
 sky130_fd_sc_hd__dfrtp_4 _09377_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00049_),
    .RESET_B(net294),
    .Q(\wb_dat_o[10] ));
 sky130_fd_sc_hd__dfrtp_4 _09378_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00050_),
    .RESET_B(net294),
    .Q(\wb_dat_o[11] ));
 sky130_fd_sc_hd__dfrtp_4 _09379_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00051_),
    .RESET_B(net294),
    .Q(\wb_dat_o[12] ));
 sky130_fd_sc_hd__dfrtp_4 _09380_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_00052_),
    .RESET_B(net294),
    .Q(\wb_dat_o[13] ));
 sky130_fd_sc_hd__dfrtp_4 _09381_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_00053_),
    .RESET_B(net294),
    .Q(\wb_dat_o[14] ));
 sky130_fd_sc_hd__dfrtp_4 _09382_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_00054_),
    .RESET_B(net294),
    .Q(\wb_dat_o[15] ));
 sky130_fd_sc_hd__dfrtp_4 _09383_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_00055_),
    .RESET_B(net293),
    .Q(\wb_dat_o[16] ));
 sky130_fd_sc_hd__dfrtp_4 _09384_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_00056_),
    .RESET_B(net292),
    .Q(\wb_dat_o[17] ));
 sky130_fd_sc_hd__dfrtp_4 _09385_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_00057_),
    .RESET_B(net293),
    .Q(\wb_dat_o[18] ));
 sky130_fd_sc_hd__dfrtp_4 _09386_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00058_),
    .RESET_B(net292),
    .Q(\wb_dat_o[19] ));
 sky130_fd_sc_hd__dfrtp_4 _09387_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_00059_),
    .RESET_B(net293),
    .Q(\wb_dat_o[20] ));
 sky130_fd_sc_hd__dfrtp_4 _09388_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(_00060_),
    .RESET_B(net300),
    .Q(\wb_dat_o[21] ));
 sky130_fd_sc_hd__dfrtp_4 _09389_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00061_),
    .RESET_B(net300),
    .Q(\wb_dat_o[22] ));
 sky130_fd_sc_hd__dfrtp_4 _09390_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00062_),
    .RESET_B(net293),
    .Q(\wb_dat_o[23] ));
 sky130_fd_sc_hd__dfrtp_4 _09391_ (.CLK(clknet_leaf_70_wbm_clk_i),
    .D(_00063_),
    .RESET_B(net300),
    .Q(\wb_dat_o[24] ));
 sky130_fd_sc_hd__dfrtp_4 _09392_ (.CLK(clknet_leaf_71_wbm_clk_i),
    .D(_00064_),
    .RESET_B(net300),
    .Q(\wb_dat_o[25] ));
 sky130_fd_sc_hd__dfrtp_4 _09393_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(_00065_),
    .RESET_B(net300),
    .Q(\wb_dat_o[26] ));
 sky130_fd_sc_hd__dfrtp_4 _09394_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(_00066_),
    .RESET_B(net300),
    .Q(\wb_dat_o[27] ));
 sky130_fd_sc_hd__dfrtp_4 _09395_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(_00067_),
    .RESET_B(net300),
    .Q(\wb_dat_o[28] ));
 sky130_fd_sc_hd__dfrtp_4 _09396_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(_00068_),
    .RESET_B(net300),
    .Q(\wb_dat_o[29] ));
 sky130_fd_sc_hd__dfrtp_4 _09397_ (.CLK(clknet_leaf_70_wbm_clk_i),
    .D(_00069_),
    .RESET_B(net302),
    .Q(\wb_dat_o[30] ));
 sky130_fd_sc_hd__dfrtp_4 _09398_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(_00070_),
    .RESET_B(net300),
    .Q(\wb_dat_o[31] ));
 sky130_fd_sc_hd__dfstp_1 _09399_ (.CLK(clknet_leaf_61_wbm_clk_i),
    .D(sclk),
    .SET_B(net272),
    .Q(\u_spi2wb.u_if.sck_l0 ));
 sky130_fd_sc_hd__dfstp_2 _09400_ (.CLK(clknet_leaf_62_wbm_clk_i),
    .D(net344),
    .SET_B(net272),
    .Q(\u_spi2wb.u_if.sck_l1 ));
 sky130_fd_sc_hd__dfstp_1 _09401_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(net364),
    .SET_B(net270),
    .Q(\u_spi2wb.u_if.sck_l2 ));
 sky130_fd_sc_hd__dfstp_1 _09402_ (.CLK(clknet_leaf_62_wbm_clk_i),
    .D(ssn),
    .SET_B(net272),
    .Q(\u_spi2wb.u_if.ssn_l0 ));
 sky130_fd_sc_hd__dfstp_2 _09403_ (.CLK(clknet_leaf_62_wbm_clk_i),
    .D(net363),
    .SET_B(net272),
    .Q(\u_spi2wb.u_if.ssn_l1 ));
 sky130_fd_sc_hd__dfrtp_1 _09404_ (.CLK(clknet_leaf_61_wbm_clk_i),
    .D(_00071_),
    .RESET_B(net274),
    .Q(\u_reset_fsm.clk_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09405_ (.CLK(clknet_leaf_61_wbm_clk_i),
    .D(_00072_),
    .RESET_B(net274),
    .Q(\u_reset_fsm.clk_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09406_ (.CLK(clknet_leaf_61_wbm_clk_i),
    .D(_00073_),
    .RESET_B(net274),
    .Q(\u_reset_fsm.clk_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09407_ (.CLK(clknet_leaf_60_wbm_clk_i),
    .D(_00074_),
    .RESET_B(net273),
    .Q(\u_reset_fsm.clk_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09408_ (.CLK(clknet_leaf_60_wbm_clk_i),
    .D(_00075_),
    .RESET_B(net273),
    .Q(\u_reset_fsm.clk_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09409_ (.CLK(clknet_leaf_60_wbm_clk_i),
    .D(_00076_),
    .RESET_B(net273),
    .Q(\u_reset_fsm.clk_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09410_ (.CLK(clknet_leaf_60_wbm_clk_i),
    .D(_00077_),
    .RESET_B(net273),
    .Q(\u_reset_fsm.clk_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09411_ (.CLK(clknet_leaf_60_wbm_clk_i),
    .D(_00078_),
    .RESET_B(net273),
    .Q(\u_reset_fsm.clk_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09412_ (.CLK(clknet_leaf_63_wbm_clk_i),
    .D(_00079_),
    .RESET_B(net272),
    .Q(\u_reset_fsm.clk_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09413_ (.CLK(clknet_leaf_62_wbm_clk_i),
    .D(_00080_),
    .RESET_B(net272),
    .Q(\u_reset_fsm.clk_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09414_ (.CLK(clknet_leaf_62_wbm_clk_i),
    .D(_00081_),
    .RESET_B(net272),
    .Q(\u_reset_fsm.clk_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09415_ (.CLK(clknet_leaf_62_wbm_clk_i),
    .D(_00082_),
    .RESET_B(net272),
    .Q(\u_reset_fsm.clk_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09416_ (.CLK(clknet_leaf_63_wbm_clk_i),
    .D(_00083_),
    .RESET_B(net275),
    .Q(\u_reset_fsm.clk_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09417_ (.CLK(clknet_leaf_61_wbm_clk_i),
    .D(_00084_),
    .RESET_B(net272),
    .Q(\u_reset_fsm.clk_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09418_ (.CLK(clknet_leaf_62_wbm_clk_i),
    .D(_00085_),
    .RESET_B(net272),
    .Q(\u_reset_fsm.clk_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09419_ (.CLK(clknet_leaf_62_wbm_clk_i),
    .D(_00086_),
    .RESET_B(net275),
    .Q(\u_reset_fsm.clk_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09420_ (.CLK(clknet_leaf_90_wbm_clk_i),
    .D(_00087_),
    .RESET_B(net260),
    .Q(\u_spi2wb.reg_be[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09421_ (.CLK(clknet_leaf_9_wbm_clk_i),
    .D(_00088_),
    .RESET_B(net260),
    .Q(\u_spi2wb.reg_be[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09422_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_00089_),
    .RESET_B(net260),
    .Q(\u_spi2wb.reg_be[2] ));
 sky130_fd_sc_hd__dfrtp_2 _09423_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_00090_),
    .RESET_B(net260),
    .Q(\u_spi2wb.reg_be[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09424_ (.CLK(clknet_leaf_75_wbm_clk_i),
    .D(_00091_),
    .RESET_B(net270),
    .Q(\u_spi2wb.u_if.cmd_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09425_ (.CLK(clknet_leaf_75_wbm_clk_i),
    .D(_00092_),
    .RESET_B(net271),
    .Q(\u_spi2wb.u_if.cmd_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09426_ (.CLK(clknet_leaf_74_wbm_clk_i),
    .D(_00093_),
    .RESET_B(net271),
    .Q(\u_spi2wb.u_if.cmd_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09427_ (.CLK(clknet_leaf_74_wbm_clk_i),
    .D(_00094_),
    .RESET_B(net270),
    .Q(\u_spi2wb.u_if.cmd_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09428_ (.CLK(clknet_leaf_1_wbm_clk_i),
    .D(_00095_),
    .RESET_B(net255),
    .Q(\u_spi2wb.reg_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09429_ (.CLK(clknet_leaf_0_wbm_clk_i),
    .D(_00096_),
    .RESET_B(net255),
    .Q(\u_spi2wb.reg_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09430_ (.CLK(clknet_leaf_1_wbm_clk_i),
    .D(_00097_),
    .RESET_B(net255),
    .Q(\u_spi2wb.reg_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09431_ (.CLK(clknet_leaf_1_wbm_clk_i),
    .D(_00098_),
    .RESET_B(net255),
    .Q(\u_spi2wb.reg_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09432_ (.CLK(clknet_leaf_1_wbm_clk_i),
    .D(_00099_),
    .RESET_B(net255),
    .Q(\u_spi2wb.reg_addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09433_ (.CLK(clknet_leaf_0_wbm_clk_i),
    .D(_00100_),
    .RESET_B(net255),
    .Q(\u_spi2wb.reg_addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09434_ (.CLK(clknet_leaf_0_wbm_clk_i),
    .D(_00101_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09435_ (.CLK(clknet_leaf_0_wbm_clk_i),
    .D(_00102_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09436_ (.CLK(clknet_leaf_0_wbm_clk_i),
    .D(_00103_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09437_ (.CLK(clknet_leaf_0_wbm_clk_i),
    .D(_00104_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09438_ (.CLK(clknet_leaf_94_wbm_clk_i),
    .D(_00105_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09439_ (.CLK(clknet_leaf_94_wbm_clk_i),
    .D(_00106_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09440_ (.CLK(clknet_leaf_0_wbm_clk_i),
    .D(_00107_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09441_ (.CLK(clknet_leaf_94_wbm_clk_i),
    .D(_00108_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09442_ (.CLK(clknet_leaf_94_wbm_clk_i),
    .D(_00109_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09443_ (.CLK(clknet_leaf_94_wbm_clk_i),
    .D(_00110_),
    .RESET_B(net254),
    .Q(\u_spi2wb.reg_addr[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09444_ (.CLK(clknet_leaf_93_wbm_clk_i),
    .D(_00111_),
    .RESET_B(net255),
    .Q(\u_spi2wb.reg_addr[16] ));
 sky130_fd_sc_hd__dfrtp_1 _09445_ (.CLK(clknet_leaf_93_wbm_clk_i),
    .D(_00112_),
    .RESET_B(net256),
    .Q(\u_spi2wb.reg_addr[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09446_ (.CLK(clknet_leaf_93_wbm_clk_i),
    .D(_00113_),
    .RESET_B(net256),
    .Q(\u_spi2wb.reg_addr[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09447_ (.CLK(clknet_leaf_93_wbm_clk_i),
    .D(_00114_),
    .RESET_B(net256),
    .Q(\u_spi2wb.reg_addr[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09448_ (.CLK(clknet_leaf_1_wbm_clk_i),
    .D(_00115_),
    .RESET_B(net255),
    .Q(\u_spi2wb.reg_wdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09449_ (.CLK(clknet_leaf_1_wbm_clk_i),
    .D(_00116_),
    .RESET_B(net255),
    .Q(\u_spi2wb.reg_wdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09450_ (.CLK(clknet_leaf_3_wbm_clk_i),
    .D(_00117_),
    .RESET_B(net256),
    .Q(\u_spi2wb.reg_wdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09451_ (.CLK(clknet_leaf_3_wbm_clk_i),
    .D(_00118_),
    .RESET_B(net256),
    .Q(\u_spi2wb.reg_wdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09452_ (.CLK(clknet_leaf_3_wbm_clk_i),
    .D(_00119_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09453_ (.CLK(clknet_leaf_3_wbm_clk_i),
    .D(_00120_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09454_ (.CLK(clknet_leaf_3_wbm_clk_i),
    .D(_00121_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09455_ (.CLK(clknet_leaf_3_wbm_clk_i),
    .D(_00122_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09456_ (.CLK(clknet_leaf_3_wbm_clk_i),
    .D(_00123_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09457_ (.CLK(clknet_leaf_3_wbm_clk_i),
    .D(_00124_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09458_ (.CLK(clknet_leaf_4_wbm_clk_i),
    .D(_00125_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09459_ (.CLK(clknet_leaf_4_wbm_clk_i),
    .D(_00126_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09460_ (.CLK(clknet_leaf_4_wbm_clk_i),
    .D(_00127_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09461_ (.CLK(clknet_leaf_4_wbm_clk_i),
    .D(_00128_),
    .RESET_B(net258),
    .Q(\u_spi2wb.reg_wdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09462_ (.CLK(clknet_leaf_4_wbm_clk_i),
    .D(_00129_),
    .RESET_B(net258),
    .Q(\u_spi2wb.reg_wdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09463_ (.CLK(clknet_leaf_6_wbm_clk_i),
    .D(_00130_),
    .RESET_B(net258),
    .Q(\u_spi2wb.reg_wdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09464_ (.CLK(clknet_leaf_6_wbm_clk_i),
    .D(_00131_),
    .RESET_B(net257),
    .Q(\u_spi2wb.reg_wdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 _09465_ (.CLK(clknet_leaf_6_wbm_clk_i),
    .D(_00132_),
    .RESET_B(net258),
    .Q(\u_spi2wb.reg_wdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09466_ (.CLK(clknet_leaf_6_wbm_clk_i),
    .D(_00133_),
    .RESET_B(net258),
    .Q(\u_spi2wb.reg_wdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09467_ (.CLK(clknet_leaf_8_wbm_clk_i),
    .D(_00134_),
    .RESET_B(net258),
    .Q(\u_spi2wb.reg_wdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09468_ (.CLK(clknet_leaf_2_wbm_clk_i),
    .D(_00135_),
    .RESET_B(net256),
    .Q(\u_spi2wb.reg_wdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 _09469_ (.CLK(clknet_leaf_2_wbm_clk_i),
    .D(_00136_),
    .RESET_B(net256),
    .Q(\u_spi2wb.reg_wdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 _09470_ (.CLK(clknet_leaf_2_wbm_clk_i),
    .D(_00137_),
    .RESET_B(net256),
    .Q(\u_spi2wb.reg_wdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 _09471_ (.CLK(clknet_leaf_2_wbm_clk_i),
    .D(_00138_),
    .RESET_B(net256),
    .Q(\u_spi2wb.reg_wdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 _09472_ (.CLK(clknet_leaf_2_wbm_clk_i),
    .D(_00139_),
    .RESET_B(net259),
    .Q(\u_spi2wb.reg_wdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 _09473_ (.CLK(clknet_leaf_92_wbm_clk_i),
    .D(_00140_),
    .RESET_B(net259),
    .Q(\u_spi2wb.reg_wdata[25] ));
 sky130_fd_sc_hd__dfrtp_1 _09474_ (.CLK(clknet_leaf_91_wbm_clk_i),
    .D(_00141_),
    .RESET_B(net264),
    .Q(\u_spi2wb.reg_wdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 _09475_ (.CLK(clknet_leaf_90_wbm_clk_i),
    .D(_00142_),
    .RESET_B(net264),
    .Q(\u_spi2wb.reg_wdata[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09476_ (.CLK(clknet_leaf_9_wbm_clk_i),
    .D(_00143_),
    .RESET_B(net264),
    .Q(\u_spi2wb.reg_wdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 _09477_ (.CLK(clknet_leaf_9_wbm_clk_i),
    .D(_00144_),
    .RESET_B(net260),
    .Q(\u_spi2wb.reg_wdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 _09478_ (.CLK(clknet_leaf_90_wbm_clk_i),
    .D(_00145_),
    .RESET_B(net264),
    .Q(\u_spi2wb.reg_wdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 _09479_ (.CLK(clknet_leaf_2_wbm_clk_i),
    .D(_00146_),
    .RESET_B(net258),
    .Q(\u_spi2wb.reg_wdata[31] ));
 sky130_fd_sc_hd__dfrtp_1 _09480_ (.CLK(clknet_leaf_61_wbm_clk_i),
    .D(net348),
    .RESET_B(net274),
    .Q(\u_reset_fsm.boot_req_ss ));
 sky130_fd_sc_hd__dfrtp_1 _09481_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(strap_sticky[31]),
    .RESET_B(net274),
    .Q(\u_reset_fsm.boot_req_s ));
 sky130_fd_sc_hd__dfrtp_1 _09482_ (.CLK(clknet_leaf_59_wbm_clk_i),
    .D(_00147_),
    .RESET_B(net273),
    .Q(\u_reset_fsm.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09483_ (.CLK(clknet_leaf_59_wbm_clk_i),
    .D(_00148_),
    .RESET_B(net273),
    .Q(\u_reset_fsm.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09484_ (.CLK(clknet_leaf_60_wbm_clk_i),
    .D(_00149_),
    .RESET_B(net273),
    .Q(\u_reset_fsm.state[2] ));
 sky130_fd_sc_hd__dfstp_1 _09485_ (.CLK(clknet_leaf_59_wbm_clk_i),
    .D(_00150_),
    .SET_B(net273),
    .Q(\u_reg.force_refclk ));
 sky130_fd_sc_hd__dfrtp_1 _09486_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(_00151_),
    .RESET_B(net273),
    .Q(\u_reg.clk_enb ));
 sky130_fd_sc_hd__dfrtp_1 _09487_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(_00152_),
    .RESET_B(net274),
    .Q(\u_reg.soft_reboot ));
 sky130_fd_sc_hd__dfrtp_4 _09488_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(_00153_),
    .RESET_B(net274),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _09489_ (.CLK(clknet_leaf_59_wbm_clk_i),
    .D(_00154_),
    .RESET_B(net274),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_4 _09490_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00155_),
    .RESET_B(net265),
    .Q(\u_reg.cfg_glb_ctrl[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09491_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00156_),
    .RESET_B(net265),
    .Q(\u_reg.cfg_glb_ctrl[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09492_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00157_),
    .RESET_B(net265),
    .Q(\u_reg.cfg_glb_ctrl[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09493_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00158_),
    .RESET_B(net265),
    .Q(\u_reg.cfg_glb_ctrl[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09494_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00159_),
    .RESET_B(net265),
    .Q(\u_reg.cfg_glb_ctrl[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09495_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00160_),
    .RESET_B(net266),
    .Q(\u_reg.cfg_glb_ctrl[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09496_ (.CLK(clknet_leaf_31_wbm_clk_i),
    .D(_00161_),
    .RESET_B(net266),
    .Q(\u_reg.cfg_glb_ctrl[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09497_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00162_),
    .RESET_B(net266),
    .Q(\u_reg.cfg_glb_ctrl[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09498_ (.CLK(clknet_leaf_28_wbm_clk_i),
    .D(_00163_),
    .RESET_B(net265),
    .Q(\u_async_wb.m_cmd_wr_data[61] ));
 sky130_fd_sc_hd__dfrtp_1 _09499_ (.CLK(clknet_leaf_28_wbm_clk_i),
    .D(_00164_),
    .RESET_B(net265),
    .Q(\u_async_wb.m_cmd_wr_data[60] ));
 sky130_fd_sc_hd__dfrtp_2 _09500_ (.CLK(clknet_leaf_23_wbm_clk_i),
    .D(_00165_),
    .RESET_B(net267),
    .Q(\u_async_wb.m_cmd_wr_data[59] ));
 sky130_fd_sc_hd__dfrtp_2 _09501_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00166_),
    .RESET_B(net267),
    .Q(\u_async_wb.m_cmd_wr_data[58] ));
 sky130_fd_sc_hd__dfrtp_1 _09502_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00167_),
    .RESET_B(net267),
    .Q(\u_async_wb.m_cmd_wr_data[57] ));
 sky130_fd_sc_hd__dfrtp_2 _09503_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00168_),
    .RESET_B(net267),
    .Q(\u_async_wb.m_cmd_wr_data[56] ));
 sky130_fd_sc_hd__dfrtp_1 _09504_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00169_),
    .RESET_B(net268),
    .Q(\u_reg.u_bank_sel.gen_bit_reg[2].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09505_ (.CLK(clknet_leaf_42_wbm_clk_i),
    .D(_00170_),
    .RESET_B(net268),
    .Q(\u_reg.u_bank_sel.gen_bit_reg[1].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09506_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00171_),
    .RESET_B(net266),
    .Q(\u_async_wb.m_cmd_wr_data[68] ));
 sky130_fd_sc_hd__dfrtp_1 _09507_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00172_),
    .RESET_B(net266),
    .Q(\u_async_wb.m_cmd_wr_data[67] ));
 sky130_fd_sc_hd__dfrtp_1 _09508_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00173_),
    .RESET_B(net266),
    .Q(\u_async_wb.m_cmd_wr_data[66] ));
 sky130_fd_sc_hd__dfstp_1 _09509_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00174_),
    .SET_B(net266),
    .Q(\u_async_wb.m_cmd_wr_data[65] ));
 sky130_fd_sc_hd__dfrtp_1 _09510_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00175_),
    .RESET_B(net265),
    .Q(\u_async_wb.m_cmd_wr_data[64] ));
 sky130_fd_sc_hd__dfrtp_1 _09511_ (.CLK(clknet_leaf_28_wbm_clk_i),
    .D(_00176_),
    .RESET_B(net265),
    .Q(\u_async_wb.m_cmd_wr_data[63] ));
 sky130_fd_sc_hd__dfrtp_1 _09512_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00177_),
    .RESET_B(net268),
    .Q(\u_reg.u_bank_sel.gen_bit_reg[0].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfxtp_1 _09513_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(_00178_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _09514_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(_00179_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _09515_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(_00180_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _09516_ (.CLK(clknet_leaf_59_wbm_clk_i),
    .D(_00181_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _09517_ (.CLK(clknet_leaf_57_wbm_clk_i),
    .D(_00182_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _09518_ (.CLK(clknet_leaf_57_wbm_clk_i),
    .D(_00183_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _09519_ (.CLK(clknet_leaf_57_wbm_clk_i),
    .D(_00184_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _09520_ (.CLK(clknet_leaf_57_wbm_clk_i),
    .D(_00185_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _09521_ (.CLK(clknet_leaf_58_wbm_clk_i),
    .D(_00186_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_1 _09522_ (.CLK(clknet_leaf_58_wbm_clk_i),
    .D(_00187_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _09523_ (.CLK(clknet_leaf_58_wbm_clk_i),
    .D(_00188_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _09524_ (.CLK(clknet_leaf_58_wbm_clk_i),
    .D(_00189_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _09525_ (.CLK(clknet_leaf_58_wbm_clk_i),
    .D(_00190_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _09526_ (.CLK(clknet_leaf_58_wbm_clk_i),
    .D(_00191_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _09527_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00192_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _09528_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00193_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _09529_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00194_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _09530_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00195_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _09531_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00196_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _09532_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00197_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _09533_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00198_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _09534_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00199_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _09535_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00200_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _09536_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00201_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _09537_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00202_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _09538_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00203_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _09539_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00204_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _09540_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00205_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_1 _09541_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00206_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _09542_ (.CLK(clknet_leaf_54_wbm_clk_i),
    .D(_00207_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _09543_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(_00208_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _09544_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(_00209_),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _09545_ (.CLK(\u_reg.cpu_ref_clk ),
    .D(_00022_),
    .RESET_B(net289),
    .Q(\u_reg.cpu_ref_clk_div_2 ));
 sky130_fd_sc_hd__dfrtp_1 _09546_ (.CLK(\u_reg.cpu_ref_clk ),
    .D(_00023_),
    .RESET_B(net290),
    .Q(\u_reg.cpu_ref_clk_div_4 ));
 sky130_fd_sc_hd__dfrtp_1 _09547_ (.CLK(\u_reg.cpu_ref_clk ),
    .D(_00024_),
    .RESET_B(net290),
    .Q(\u_reg.cpu_ref_clk_div_8 ));
 sky130_fd_sc_hd__dfrtp_1 _09548_ (.CLK(clknet_leaf_28_wbm_clk_i),
    .D(_00210_),
    .RESET_B(net265),
    .Q(\u_async_wb.m_cmd_wr_data[62] ));
 sky130_fd_sc_hd__dfrtp_1 _09549_ (.CLK(\u_reg.u_wbclk.mclk ),
    .D(_00025_),
    .RESET_B(net290),
    .Q(\u_reg.u_wbclk.clk_div_2 ));
 sky130_fd_sc_hd__dfrtp_1 _09550_ (.CLK(\u_reg.u_wbclk.mclk ),
    .D(_00026_),
    .RESET_B(net290),
    .Q(\u_reg.u_wbclk.clk_div_4 ));
 sky130_fd_sc_hd__dfrtp_1 _09551_ (.CLK(\u_reg.u_wbclk.mclk ),
    .D(_00027_),
    .RESET_B(net290),
    .Q(\u_reg.u_wbclk.clk_div_8 ));
 sky130_fd_sc_hd__dfxtp_1 _09552_ (.CLK(clknet_leaf_57_wbm_clk_i),
    .D(_00211_),
    .Q(\u_reg.cfg_clk_ctrl[0] ));
 sky130_fd_sc_hd__dfxtp_1 _09553_ (.CLK(clknet_leaf_58_wbm_clk_i),
    .D(_00212_),
    .Q(\u_reg.cfg_clk_ctrl[1] ));
 sky130_fd_sc_hd__dfxtp_1 _09554_ (.CLK(clknet_leaf_58_wbm_clk_i),
    .D(_00213_),
    .Q(\u_reg.cfg_clk_ctrl[2] ));
 sky130_fd_sc_hd__dfxtp_1 _09555_ (.CLK(clknet_leaf_57_wbm_clk_i),
    .D(_00214_),
    .Q(\u_reg.cfg_clk_ctrl[3] ));
 sky130_fd_sc_hd__dfxtp_1 _09556_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00215_),
    .Q(\u_reg.cfg_clk_ctrl[4] ));
 sky130_fd_sc_hd__dfxtp_1 _09557_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00216_),
    .Q(\u_reg.cfg_clk_ctrl[5] ));
 sky130_fd_sc_hd__dfxtp_1 _09558_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00217_),
    .Q(\u_reg.cfg_clk_ctrl[6] ));
 sky130_fd_sc_hd__dfxtp_1 _09559_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00218_),
    .Q(\u_reg.cfg_clk_ctrl[7] ));
 sky130_fd_sc_hd__dfxtp_1 _09560_ (.CLK(clknet_leaf_34_wbm_clk_i),
    .D(_00219_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _09561_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00220_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _09562_ (.CLK(clknet_leaf_34_wbm_clk_i),
    .D(_00221_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _09563_ (.CLK(clknet_leaf_34_wbm_clk_i),
    .D(_00222_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _09564_ (.CLK(clknet_leaf_31_wbm_clk_i),
    .D(_00223_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _09565_ (.CLK(clknet_leaf_31_wbm_clk_i),
    .D(_00224_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _09566_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00225_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _09567_ (.CLK(clknet_leaf_31_wbm_clk_i),
    .D(_00226_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _09568_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00227_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _09569_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00228_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _09570_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00229_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _09571_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00230_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _09572_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00231_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _09573_ (.CLK(clknet_leaf_31_wbm_clk_i),
    .D(_00232_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _09574_ (.CLK(clknet_leaf_31_wbm_clk_i),
    .D(_00233_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _09575_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00234_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _09576_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00235_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _09577_ (.CLK(clknet_leaf_36_wbm_clk_i),
    .D(_00236_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _09578_ (.CLK(clknet_leaf_36_wbm_clk_i),
    .D(_00237_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_2 _09579_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00238_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _09580_ (.CLK(clknet_leaf_52_wbm_clk_i),
    .D(_00239_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _09581_ (.CLK(clknet_leaf_52_wbm_clk_i),
    .D(_00240_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _09582_ (.CLK(clknet_leaf_52_wbm_clk_i),
    .D(_00241_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _09583_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00242_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _09584_ (.CLK(clknet_leaf_52_wbm_clk_i),
    .D(_00243_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _09585_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00244_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _09586_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00245_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _09587_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00246_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _09588_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00247_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _09589_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00248_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _09590_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00249_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _09591_ (.CLK(clknet_leaf_52_wbm_clk_i),
    .D(_00250_),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _09592_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00251_),
    .RESET_B(net289),
    .Q(\u_reg.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09593_ (.CLK(clknet_leaf_49_wbm_clk_i),
    .D(_00252_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09594_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00253_),
    .RESET_B(net289),
    .Q(\u_reg.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09595_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00254_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09596_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00255_),
    .RESET_B(net289),
    .Q(\u_reg.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09597_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00256_),
    .RESET_B(net289),
    .Q(\u_reg.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09598_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00257_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09599_ (.CLK(clknet_leaf_56_wbm_clk_i),
    .D(_00258_),
    .RESET_B(net289),
    .Q(\u_reg.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09600_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00259_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09601_ (.CLK(clknet_leaf_57_wbm_clk_i),
    .D(_00260_),
    .RESET_B(net289),
    .Q(\u_reg.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09602_ (.CLK(clknet_leaf_57_wbm_clk_i),
    .D(_00261_),
    .RESET_B(net289),
    .Q(\u_reg.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09603_ (.CLK(clknet_leaf_39_wbm_clk_i),
    .D(_00262_),
    .RESET_B(net286),
    .Q(\u_reg.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09604_ (.CLK(clknet_leaf_39_wbm_clk_i),
    .D(_00263_),
    .RESET_B(net286),
    .Q(\u_reg.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09605_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00264_),
    .RESET_B(net286),
    .Q(\u_reg.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09606_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00265_),
    .RESET_B(net289),
    .Q(\u_reg.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09607_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00266_),
    .RESET_B(net286),
    .Q(\u_reg.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09608_ (.CLK(clknet_leaf_50_wbm_clk_i),
    .D(_00267_),
    .RESET_B(net286),
    .Q(\u_reg.reg_rdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 _09609_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00268_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09610_ (.CLK(clknet_leaf_50_wbm_clk_i),
    .D(_00269_),
    .RESET_B(net286),
    .Q(\u_reg.reg_rdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09611_ (.CLK(clknet_leaf_48_wbm_clk_i),
    .D(_00270_),
    .RESET_B(net286),
    .Q(\u_reg.reg_rdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09612_ (.CLK(clknet_leaf_50_wbm_clk_i),
    .D(_00271_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 _09613_ (.CLK(clknet_leaf_50_wbm_clk_i),
    .D(_00272_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 _09614_ (.CLK(clknet_leaf_50_wbm_clk_i),
    .D(_00273_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 _09615_ (.CLK(clknet_leaf_50_wbm_clk_i),
    .D(_00274_),
    .RESET_B(net286),
    .Q(\u_reg.reg_rdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 _09616_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00275_),
    .RESET_B(net288),
    .Q(\u_reg.reg_rdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 _09617_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00276_),
    .RESET_B(net288),
    .Q(\u_reg.reg_rdata[25] ));
 sky130_fd_sc_hd__dfrtp_1 _09618_ (.CLK(clknet_leaf_53_wbm_clk_i),
    .D(_00277_),
    .RESET_B(net288),
    .Q(\u_reg.reg_rdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 _09619_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00278_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09620_ (.CLK(clknet_leaf_49_wbm_clk_i),
    .D(_00279_),
    .RESET_B(net287),
    .Q(\u_reg.reg_rdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 _09621_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00280_),
    .RESET_B(net288),
    .Q(\u_reg.reg_rdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 _09622_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00281_),
    .RESET_B(net288),
    .Q(\u_reg.reg_rdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 _09623_ (.CLK(clknet_leaf_55_wbm_clk_i),
    .D(_00282_),
    .RESET_B(net289),
    .Q(\u_reg.reg_rdata[31] ));
 sky130_fd_sc_hd__dfrtp_1 _09624_ (.CLK(clknet_leaf_48_wbm_clk_i),
    .D(_00020_),
    .RESET_B(net286),
    .Q(\u_reg.reg_ack ));
 sky130_fd_sc_hd__dfrtp_1 _09625_ (.CLK(clknet_leaf_68_wbm_clk_i),
    .D(_00283_),
    .RESET_B(net303),
    .Q(\u_async_wb.u_resp_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09626_ (.CLK(clknet_leaf_68_wbm_clk_i),
    .D(_00284_),
    .RESET_B(net302),
    .Q(\u_async_wb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _09627_ (.CLK(clknet_leaf_36_wbm_clk_i),
    .D(_00285_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _09628_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00286_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _09629_ (.CLK(clknet_leaf_34_wbm_clk_i),
    .D(_00287_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_2 _09630_ (.CLK(clknet_leaf_36_wbm_clk_i),
    .D(_00288_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_2 _09631_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00289_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_2 _09632_ (.CLK(clknet_leaf_34_wbm_clk_i),
    .D(_00290_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _09633_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00291_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _09634_ (.CLK(clknet_leaf_34_wbm_clk_i),
    .D(_00292_),
    .Q(net2));
 sky130_fd_sc_hd__dfxtp_1 _09635_ (.CLK(clknet_leaf_37_wbm_clk_i),
    .D(_00293_),
    .Q(net3));
 sky130_fd_sc_hd__dfxtp_1 _09636_ (.CLK(clknet_leaf_36_wbm_clk_i),
    .D(_00294_),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_1 _09637_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00295_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_1 _09638_ (.CLK(clknet_leaf_35_wbm_clk_i),
    .D(_00296_),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_1 _09639_ (.CLK(clknet_leaf_37_wbm_clk_i),
    .D(_00297_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _09640_ (.CLK(clknet_leaf_37_wbm_clk_i),
    .D(_00298_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _09641_ (.CLK(clknet_leaf_37_wbm_clk_i),
    .D(_00299_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _09642_ (.CLK(clknet_leaf_37_wbm_clk_i),
    .D(_00300_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _09643_ (.CLK(clknet_leaf_37_wbm_clk_i),
    .D(_00301_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _09644_ (.CLK(clknet_leaf_37_wbm_clk_i),
    .D(_00302_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _09645_ (.CLK(clknet_leaf_52_wbm_clk_i),
    .D(_00303_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _09646_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00304_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_2 _09647_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00305_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _09648_ (.CLK(\clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00306_),
    .Q(\u_async_wb.u_resp_if.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _09649_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00307_),
    .Q(\u_async_wb.u_resp_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _09650_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00308_),
    .Q(\u_async_wb.u_resp_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _09651_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00309_),
    .Q(\u_async_wb.u_resp_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _09652_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00310_),
    .Q(\u_async_wb.u_resp_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _09653_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00311_),
    .Q(\u_async_wb.u_resp_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _09654_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00312_),
    .Q(\u_async_wb.u_resp_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _09655_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00313_),
    .Q(\u_async_wb.u_resp_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _09656_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00314_),
    .Q(\u_async_wb.u_resp_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _09657_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00315_),
    .Q(\u_async_wb.u_resp_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _09658_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00316_),
    .Q(\u_async_wb.u_resp_if.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _09659_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00317_),
    .Q(\u_async_wb.u_resp_if.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _09660_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00318_),
    .Q(\u_async_wb.u_resp_if.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _09661_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00319_),
    .Q(\u_async_wb.u_resp_if.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _09662_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00320_),
    .Q(\u_async_wb.u_resp_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _09663_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00321_),
    .Q(\u_async_wb.u_resp_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _09664_ (.CLK(\clknet_3_3__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00322_),
    .Q(\u_async_wb.u_resp_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _09665_ (.CLK(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00323_),
    .Q(\u_async_wb.u_resp_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _09666_ (.CLK(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00324_),
    .Q(\u_async_wb.u_resp_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _09667_ (.CLK(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00325_),
    .Q(\u_async_wb.u_resp_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _09668_ (.CLK(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00326_),
    .Q(\u_async_wb.u_resp_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _09669_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00327_),
    .Q(\u_async_wb.u_resp_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _09670_ (.CLK(\clknet_3_3__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00328_),
    .Q(\u_async_wb.u_resp_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _09671_ (.CLK(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00329_),
    .Q(\u_async_wb.u_resp_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _09672_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00330_),
    .Q(\u_async_wb.u_resp_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _09673_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00331_),
    .Q(\u_async_wb.u_resp_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _09674_ (.CLK(\clknet_3_3__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00332_),
    .Q(\u_async_wb.u_resp_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _09675_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00333_),
    .Q(\u_async_wb.u_resp_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _09676_ (.CLK(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00334_),
    .Q(\u_async_wb.u_resp_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _09677_ (.CLK(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00335_),
    .Q(\u_async_wb.u_resp_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _09678_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00336_),
    .Q(\u_async_wb.u_resp_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _09679_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00337_),
    .Q(\u_async_wb.u_resp_if.mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _09680_ (.CLK(\clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00338_),
    .Q(\u_async_wb.u_resp_if.mem[1][32] ));
 sky130_fd_sc_hd__dfstp_1 _09681_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00015_),
    .SET_B(net246),
    .Q(\u_uart2wb.u_core.u_txfsm.txstate[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09682_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00016_),
    .RESET_B(net247),
    .Q(\u_uart2wb.u_core.u_txfsm.txstate[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09683_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00017_),
    .RESET_B(net246),
    .Q(\u_uart2wb.u_core.u_txfsm.txstate[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09684_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_00018_),
    .RESET_B(net247),
    .Q(\u_uart2wb.u_core.u_txfsm.txstate[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09685_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00019_),
    .RESET_B(net247),
    .Q(\u_uart2wb.u_core.u_txfsm.txstate[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09686_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(net362),
    .RESET_B(net252),
    .Q(\u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09687_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(net361),
    .RESET_B(net253),
    .Q(\u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09688_ (.CLK(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(net353),
    .RESET_B(\u_async_wb.u_cmd_if.rd_reset_n ),
    .Q(\u_async_wb.u_cmd_if.sync_wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09689_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(\u_async_wb.u_cmd_if.grey_wr_ptr[0] ),
    .RESET_B(net252),
    .Q(\u_async_wb.u_cmd_if.sync_wr_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09690_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(\u_async_wb.u_cmd_if.grey_wr_ptr[1] ),
    .RESET_B(net252),
    .Q(\u_async_wb.u_cmd_if.sync_wr_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09691_ (.CLK(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(\u_async_wb.u_cmd_if.grey_wr_ptr[2] ),
    .RESET_B(net252),
    .Q(\u_async_wb.u_cmd_if.sync_wr_ptr_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09692_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00339_),
    .RESET_B(net252),
    .Q(\u_async_wb.u_cmd_if.grey_rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09693_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00340_),
    .RESET_B(net252),
    .Q(\u_async_wb.u_cmd_if.grey_rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09694_ (.CLK(clknet_leaf_46_wbm_clk_i),
    .D(_00341_),
    .RESET_B(net305),
    .Q(\u_async_wb.PendingRd ));
 sky130_fd_sc_hd__dfrtp_1 _09695_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00342_),
    .RESET_B(net305),
    .Q(\u_async_wb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09696_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00343_),
    .RESET_B(net305),
    .Q(\u_async_wb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09697_ (.CLK(clknet_leaf_46_wbm_clk_i),
    .D(\u_async_wb.u_cmd_if.grey_rd_ptr[0] ),
    .RESET_B(net305),
    .Q(\u_async_wb.u_cmd_if.sync_rd_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09698_ (.CLK(clknet_leaf_70_wbm_clk_i),
    .D(\u_async_wb.u_cmd_if.grey_rd_ptr[1] ),
    .RESET_B(net305),
    .Q(\u_async_wb.u_cmd_if.sync_rd_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09699_ (.CLK(clknet_leaf_70_wbm_clk_i),
    .D(\u_async_wb.u_cmd_if.grey_rd_ptr[2] ),
    .RESET_B(net302),
    .Q(\u_async_wb.u_cmd_if.sync_rd_ptr_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09700_ (.CLK(clknet_leaf_70_wbm_clk_i),
    .D(net343),
    .RESET_B(net305),
    .Q(\u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09701_ (.CLK(clknet_leaf_70_wbm_clk_i),
    .D(net356),
    .RESET_B(net305),
    .Q(\u_async_wb.u_cmd_if.sync_rd_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09702_ (.CLK(clknet_leaf_70_wbm_clk_i),
    .D(net357),
    .RESET_B(net302),
    .Q(\u_async_wb.u_cmd_if.sync_rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09703_ (.CLK(clknet_leaf_46_wbm_clk_i),
    .D(_00344_),
    .RESET_B(net305),
    .Q(\u_async_wb.u_cmd_if.grey_wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09704_ (.CLK(clknet_leaf_46_wbm_clk_i),
    .D(_00345_),
    .RESET_B(net305),
    .Q(\u_async_wb.u_cmd_if.grey_wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _09705_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00346_),
    .RESET_B(net305),
    .Q(\u_async_wb.u_cmd_if.grey_wr_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _09706_ (.CLK(\clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00347_),
    .Q(\u_async_wb.u_resp_if.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _09707_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00348_),
    .Q(\u_async_wb.u_resp_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _09708_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00349_),
    .Q(\u_async_wb.u_resp_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _09709_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00350_),
    .Q(\u_async_wb.u_resp_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _09710_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00351_),
    .Q(\u_async_wb.u_resp_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _09711_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00352_),
    .Q(\u_async_wb.u_resp_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _09712_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00353_),
    .Q(\u_async_wb.u_resp_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _09713_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00354_),
    .Q(\u_async_wb.u_resp_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _09714_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00355_),
    .Q(\u_async_wb.u_resp_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _09715_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00356_),
    .Q(\u_async_wb.u_resp_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _09716_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00357_),
    .Q(\u_async_wb.u_resp_if.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _09717_ (.CLK(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00358_),
    .Q(\u_async_wb.u_resp_if.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _09718_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00359_),
    .Q(\u_async_wb.u_resp_if.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _09719_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00360_),
    .Q(\u_async_wb.u_resp_if.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _09720_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00361_),
    .Q(\u_async_wb.u_resp_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _09721_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00362_),
    .Q(\u_async_wb.u_resp_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _09722_ (.CLK(\clknet_3_3__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00363_),
    .Q(\u_async_wb.u_resp_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _09723_ (.CLK(\clknet_3_3__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00364_),
    .Q(\u_async_wb.u_resp_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _09724_ (.CLK(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00365_),
    .Q(\u_async_wb.u_resp_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _09725_ (.CLK(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00366_),
    .Q(\u_async_wb.u_resp_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _09726_ (.CLK(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00367_),
    .Q(\u_async_wb.u_resp_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _09727_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00368_),
    .Q(\u_async_wb.u_resp_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _09728_ (.CLK(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00369_),
    .Q(\u_async_wb.u_resp_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _09729_ (.CLK(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00370_),
    .Q(\u_async_wb.u_resp_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _09730_ (.CLK(\clknet_3_3__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00371_),
    .Q(\u_async_wb.u_resp_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _09731_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00372_),
    .Q(\u_async_wb.u_resp_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _09732_ (.CLK(\clknet_3_3__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00373_),
    .Q(\u_async_wb.u_resp_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _09733_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00374_),
    .Q(\u_async_wb.u_resp_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _09734_ (.CLK(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00375_),
    .Q(\u_async_wb.u_resp_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _09735_ (.CLK(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00376_),
    .Q(\u_async_wb.u_resp_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _09736_ (.CLK(\clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00377_),
    .Q(\u_async_wb.u_resp_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _09737_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00378_),
    .Q(\u_async_wb.u_resp_if.mem[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _09738_ (.CLK(\clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00379_),
    .Q(\u_async_wb.u_resp_if.mem[0][32] ));
 sky130_fd_sc_hd__dfrtp_1 _09739_ (.CLK(clknet_leaf_68_wbm_clk_i),
    .D(_00380_),
    .RESET_B(net302),
    .Q(\u_async_wb.u_resp_if.grey_rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09740_ (.CLK(clknet_leaf_67_wbm_clk_i),
    .D(_00381_),
    .RESET_B(net302),
    .Q(\u_async_wb.u_resp_if.grey_rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09741_ (.CLK(clknet_leaf_67_wbm_clk_i),
    .D(net346),
    .RESET_B(net302),
    .Q(\u_async_wb.u_resp_if.sync_wr_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09742_ (.CLK(clknet_leaf_69_wbm_clk_i),
    .D(net358),
    .RESET_B(net302),
    .Q(\u_async_wb.u_resp_if.sync_wr_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09743_ (.CLK(clknet_leaf_69_wbm_clk_i),
    .D(\u_async_wb.u_resp_if.grey_wr_ptr[0] ),
    .RESET_B(net302),
    .Q(\u_async_wb.u_resp_if.sync_wr_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09744_ (.CLK(clknet_leaf_69_wbm_clk_i),
    .D(\u_async_wb.u_resp_if.grey_wr_ptr[1] ),
    .RESET_B(net302),
    .Q(\u_async_wb.u_resp_if.sync_wr_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09745_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00382_),
    .RESET_B(net252),
    .Q(\u_async_wb.u_cmd_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09746_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00383_),
    .RESET_B(net252),
    .Q(\u_async_wb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _09747_ (.CLK(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00384_),
    .RESET_B(net252),
    .Q(\u_async_wb.u_cmd_if.grey_rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09748_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00385_),
    .RESET_B(net253),
    .Q(\u_async_wb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09749_ (.CLK(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00386_),
    .RESET_B(net253),
    .Q(\u_async_wb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09750_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(\u_async_wb.u_resp_if.grey_rd_ptr[0] ),
    .RESET_B(net253),
    .Q(\u_async_wb.u_resp_if.sync_rd_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09751_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(\u_async_wb.u_resp_if.grey_rd_ptr[1] ),
    .RESET_B(net253),
    .Q(\u_async_wb.u_resp_if.sync_rd_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09752_ (.CLK(\clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(net351),
    .RESET_B(net253),
    .Q(\u_async_wb.u_resp_if.sync_rd_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09753_ (.CLK(\clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(net350),
    .RESET_B(net253),
    .Q(\u_async_wb.u_resp_if.sync_rd_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09754_ (.CLK(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00387_),
    .RESET_B(net253),
    .Q(\u_async_wb.u_resp_if.grey_wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09755_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(_00388_),
    .RESET_B(net253),
    .Q(\u_async_wb.u_resp_if.grey_wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09756_ (.CLK(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(wbs_ack_i),
    .RESET_B(net252),
    .Q(\u_async_wb.wbs_ack_f ));
 sky130_fd_sc_hd__dfrtp_1 _09757_ (.CLK(clknet_leaf_92_wbm_clk_i),
    .D(_00389_),
    .RESET_B(net295),
    .Q(\u_arb.gnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09758_ (.CLK(clknet_leaf_92_wbm_clk_i),
    .D(_00390_),
    .RESET_B(net295),
    .Q(\u_arb.gnt[1] ));
 sky130_fd_sc_hd__dfstp_1 _09759_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(net368),
    .SET_B(net270),
    .Q(\u_spi2wb.u_if.spi_if_st[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09760_ (.CLK(clknet_leaf_73_wbm_clk_i),
    .D(_00002_),
    .RESET_B(net271),
    .Q(\u_spi2wb.u_if.spi_if_st[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09761_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(_00003_),
    .RESET_B(net271),
    .Q(\u_spi2wb.u_if.adr_phase ));
 sky130_fd_sc_hd__dfrtp_1 _09762_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(_00004_),
    .RESET_B(net270),
    .Q(\u_spi2wb.u_if.rd_phase ));
 sky130_fd_sc_hd__dfrtp_1 _09763_ (.CLK(clknet_leaf_73_wbm_clk_i),
    .D(_00005_),
    .RESET_B(net271),
    .Q(\u_spi2wb.u_if.cmd_phase ));
 sky130_fd_sc_hd__dfrtp_1 _09764_ (.CLK(clknet_leaf_73_wbm_clk_i),
    .D(_00006_),
    .RESET_B(net270),
    .Q(\u_spi2wb.u_if.spi_if_st[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09765_ (.CLK(clknet_leaf_74_wbm_clk_i),
    .D(_00007_),
    .RESET_B(net270),
    .Q(\u_spi2wb.u_if.wr_phase ));
 sky130_fd_sc_hd__dfrtp_1 _09766_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00391_),
    .RESET_B(net246),
    .Q(\u_uart2wb.u_msg.wait_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09767_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00392_),
    .RESET_B(net246),
    .Q(\u_uart2wb.u_msg.wait_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09768_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00393_),
    .RESET_B(net246),
    .Q(\u_uart2wb.u_msg.wait_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09769_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00394_),
    .RESET_B(net247),
    .Q(\u_uart2wb.u_msg.wait_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09770_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00395_),
    .RESET_B(net246),
    .Q(\u_uart2wb.u_msg.wait_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09771_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00396_),
    .RESET_B(net246),
    .Q(\u_uart2wb.u_msg.wait_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09772_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00397_),
    .RESET_B(net248),
    .Q(\u_uart2wb.u_msg.wait_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09773_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00398_),
    .RESET_B(net248),
    .Q(\u_uart2wb.u_msg.wait_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09774_ (.CLK(clknet_leaf_90_wbm_clk_i),
    .D(wb_ack_o1),
    .RESET_B(net295),
    .Q(wb_ack_o));
 sky130_fd_sc_hd__dfrtp_1 _09775_ (.CLK(clknet_leaf_93_wbm_clk_i),
    .D(wb_err_o1),
    .RESET_B(net295),
    .Q(wb_err_o));
 sky130_fd_sc_hd__dfrtp_4 _09776_ (.CLK(clknet_leaf_90_wbm_clk_i),
    .D(_00000_),
    .RESET_B(net295),
    .Q(wb_req));
 sky130_fd_sc_hd__dfrtp_1 _09777_ (.CLK(\clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(net347),
    .RESET_B(net303),
    .Q(\u_wbs_rst.in_data_2s ));
 sky130_fd_sc_hd__dfrtp_1 _09778_ (.CLK(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ),
    .D(net318),
    .RESET_B(net303),
    .Q(\u_wbs_rst.in_data_s ));
 sky130_fd_sc_hd__conb_1 _09778__318 (.HI(net318));
 sky130_fd_sc_hd__dfrtp_1 _09779_ (.CLK(clknet_leaf_94_wbm_clk_i),
    .D(net352),
    .RESET_B(_00036_),
    .Q(\u_wbm_rst.in_data_2s ));
 sky130_fd_sc_hd__dfrtp_1 _09780_ (.CLK(clknet_leaf_94_wbm_clk_i),
    .D(net317),
    .RESET_B(_00037_),
    .Q(\u_wbm_rst.in_data_s ));
 sky130_fd_sc_hd__conb_1 _09780__317 (.HI(net317));
 sky130_fd_sc_hd__dfxtp_1 _09781_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_00399_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[56] ));
 sky130_fd_sc_hd__dfxtp_1 _09782_ (.CLK(\clknet_leaf_14_u_uart2wb.baud_clk_16x ),
    .D(_00400_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[57] ));
 sky130_fd_sc_hd__dfxtp_1 _09783_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_00401_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[58] ));
 sky130_fd_sc_hd__dfxtp_1 _09784_ (.CLK(\clknet_leaf_14_u_uart2wb.baud_clk_16x ),
    .D(_00402_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[59] ));
 sky130_fd_sc_hd__dfxtp_1 _09785_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_00403_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[60] ));
 sky130_fd_sc_hd__dfxtp_1 _09786_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_00404_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[61] ));
 sky130_fd_sc_hd__dfxtp_1 _09787_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_00405_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[62] ));
 sky130_fd_sc_hd__dfxtp_1 _09788_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_00406_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[120] ));
 sky130_fd_sc_hd__dfxtp_1 _09789_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_00407_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[121] ));
 sky130_fd_sc_hd__dfxtp_1 _09790_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00408_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[122] ));
 sky130_fd_sc_hd__dfxtp_1 _09791_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00409_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[123] ));
 sky130_fd_sc_hd__dfxtp_1 _09792_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00410_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[124] ));
 sky130_fd_sc_hd__dfxtp_1 _09793_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00411_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[125] ));
 sky130_fd_sc_hd__dfxtp_1 _09794_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00412_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[126] ));
 sky130_fd_sc_hd__dfxtp_1 _09795_ (.CLK(\clknet_leaf_8_u_uart2wb.baud_clk_16x ),
    .D(_00413_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[72] ));
 sky130_fd_sc_hd__dfxtp_1 _09796_ (.CLK(\clknet_leaf_14_u_uart2wb.baud_clk_16x ),
    .D(_00414_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[73] ));
 sky130_fd_sc_hd__dfxtp_1 _09797_ (.CLK(\clknet_leaf_8_u_uart2wb.baud_clk_16x ),
    .D(_00415_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[74] ));
 sky130_fd_sc_hd__dfxtp_1 _09798_ (.CLK(\clknet_leaf_7_u_uart2wb.baud_clk_16x ),
    .D(_00416_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[75] ));
 sky130_fd_sc_hd__dfxtp_1 _09799_ (.CLK(\clknet_leaf_7_u_uart2wb.baud_clk_16x ),
    .D(_00417_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[76] ));
 sky130_fd_sc_hd__dfxtp_1 _09800_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00418_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[77] ));
 sky130_fd_sc_hd__dfxtp_1 _09801_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00419_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[78] ));
 sky130_fd_sc_hd__dfxtp_1 _09802_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00420_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[80] ));
 sky130_fd_sc_hd__dfxtp_1 _09803_ (.CLK(\clknet_leaf_9_u_uart2wb.baud_clk_16x ),
    .D(_00421_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[81] ));
 sky130_fd_sc_hd__dfxtp_1 _09804_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_00422_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[82] ));
 sky130_fd_sc_hd__dfxtp_1 _09805_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00423_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[83] ));
 sky130_fd_sc_hd__dfxtp_1 _09806_ (.CLK(\clknet_leaf_7_u_uart2wb.baud_clk_16x ),
    .D(_00424_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[84] ));
 sky130_fd_sc_hd__dfxtp_1 _09807_ (.CLK(\clknet_leaf_7_u_uart2wb.baud_clk_16x ),
    .D(_00425_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[85] ));
 sky130_fd_sc_hd__dfxtp_1 _09808_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00426_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[86] ));
 sky130_fd_sc_hd__dfxtp_1 _09809_ (.CLK(\clknet_leaf_9_u_uart2wb.baud_clk_16x ),
    .D(_00427_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[96] ));
 sky130_fd_sc_hd__dfxtp_1 _09810_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00428_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[97] ));
 sky130_fd_sc_hd__dfxtp_1 _09811_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_00429_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[98] ));
 sky130_fd_sc_hd__dfxtp_1 _09812_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_00430_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[99] ));
 sky130_fd_sc_hd__dfxtp_1 _09813_ (.CLK(\clknet_leaf_9_u_uart2wb.baud_clk_16x ),
    .D(_00431_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[100] ));
 sky130_fd_sc_hd__dfxtp_1 _09814_ (.CLK(\clknet_leaf_9_u_uart2wb.baud_clk_16x ),
    .D(_00432_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[101] ));
 sky130_fd_sc_hd__dfxtp_1 _09815_ (.CLK(\clknet_leaf_14_u_uart2wb.baud_clk_16x ),
    .D(_00433_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[102] ));
 sky130_fd_sc_hd__dfxtp_1 _09816_ (.CLK(\clknet_leaf_9_u_uart2wb.baud_clk_16x ),
    .D(_00434_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[104] ));
 sky130_fd_sc_hd__dfxtp_1 _09817_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00435_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[105] ));
 sky130_fd_sc_hd__dfxtp_1 _09818_ (.CLK(\clknet_leaf_14_u_uart2wb.baud_clk_16x ),
    .D(_00436_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[106] ));
 sky130_fd_sc_hd__dfxtp_1 _09819_ (.CLK(\clknet_leaf_9_u_uart2wb.baud_clk_16x ),
    .D(_00437_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[107] ));
 sky130_fd_sc_hd__dfxtp_1 _09820_ (.CLK(\clknet_leaf_14_u_uart2wb.baud_clk_16x ),
    .D(_00438_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[108] ));
 sky130_fd_sc_hd__dfxtp_1 _09821_ (.CLK(\clknet_leaf_9_u_uart2wb.baud_clk_16x ),
    .D(_00439_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[109] ));
 sky130_fd_sc_hd__dfxtp_1 _09822_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00440_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[110] ));
 sky130_fd_sc_hd__dfxtp_1 _09823_ (.CLK(\clknet_leaf_14_u_uart2wb.baud_clk_16x ),
    .D(_00441_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[112] ));
 sky130_fd_sc_hd__dfxtp_1 _09824_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00442_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[113] ));
 sky130_fd_sc_hd__dfxtp_1 _09825_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00443_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[114] ));
 sky130_fd_sc_hd__dfxtp_1 _09826_ (.CLK(\clknet_leaf_12_u_uart2wb.baud_clk_16x ),
    .D(_00444_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[115] ));
 sky130_fd_sc_hd__dfxtp_1 _09827_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00445_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[116] ));
 sky130_fd_sc_hd__dfxtp_1 _09828_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00446_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[117] ));
 sky130_fd_sc_hd__dfxtp_1 _09829_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00447_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[118] ));
 sky130_fd_sc_hd__dfxtp_1 _09830_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00448_),
    .Q(\u_async_wb.u_cmd_if.mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _09831_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00449_),
    .Q(\u_async_wb.u_cmd_if.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _09832_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00450_),
    .Q(\u_async_wb.u_cmd_if.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _09833_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00451_),
    .Q(\u_async_wb.u_cmd_if.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _09834_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00452_),
    .Q(\u_async_wb.u_cmd_if.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _09835_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00453_),
    .Q(\u_async_wb.u_cmd_if.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _09836_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00454_),
    .Q(\u_async_wb.u_cmd_if.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _09837_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00455_),
    .Q(\u_async_wb.u_cmd_if.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _09838_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00456_),
    .Q(\u_async_wb.u_cmd_if.mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _09839_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00457_),
    .Q(\u_async_wb.u_cmd_if.mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _09840_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00458_),
    .Q(\u_async_wb.u_cmd_if.mem[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _09841_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00459_),
    .Q(\u_async_wb.u_cmd_if.mem[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _09842_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00460_),
    .Q(\u_async_wb.u_cmd_if.mem[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _09843_ (.CLK(clknet_leaf_29_wbm_clk_i),
    .D(_00461_),
    .Q(\u_async_wb.u_cmd_if.mem[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _09844_ (.CLK(clknet_leaf_29_wbm_clk_i),
    .D(_00462_),
    .Q(\u_async_wb.u_cmd_if.mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _09845_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00463_),
    .Q(\u_async_wb.u_cmd_if.mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _09846_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00464_),
    .Q(\u_async_wb.u_cmd_if.mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _09847_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00465_),
    .Q(\u_async_wb.u_cmd_if.mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _09848_ (.CLK(clknet_leaf_31_wbm_clk_i),
    .D(_00466_),
    .Q(\u_async_wb.u_cmd_if.mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _09849_ (.CLK(clknet_leaf_41_wbm_clk_i),
    .D(_00467_),
    .Q(\u_async_wb.u_cmd_if.mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _09850_ (.CLK(clknet_leaf_41_wbm_clk_i),
    .D(_00468_),
    .Q(\u_async_wb.u_cmd_if.mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _09851_ (.CLK(clknet_leaf_41_wbm_clk_i),
    .D(_00469_),
    .Q(\u_async_wb.u_cmd_if.mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _09852_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00470_),
    .Q(\u_async_wb.u_cmd_if.mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _09853_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00471_),
    .Q(\u_async_wb.u_cmd_if.mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _09854_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00472_),
    .Q(\u_async_wb.u_cmd_if.mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _09855_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00473_),
    .Q(\u_async_wb.u_cmd_if.mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _09856_ (.CLK(clknet_leaf_43_wbm_clk_i),
    .D(_00474_),
    .Q(\u_async_wb.u_cmd_if.mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _09857_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00475_),
    .Q(\u_async_wb.u_cmd_if.mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _09858_ (.CLK(clknet_leaf_43_wbm_clk_i),
    .D(_00476_),
    .Q(\u_async_wb.u_cmd_if.mem[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _09859_ (.CLK(clknet_leaf_47_wbm_clk_i),
    .D(_00477_),
    .Q(\u_async_wb.u_cmd_if.mem[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _09860_ (.CLK(clknet_leaf_47_wbm_clk_i),
    .D(_00478_),
    .Q(\u_async_wb.u_cmd_if.mem[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _09861_ (.CLK(clknet_leaf_47_wbm_clk_i),
    .D(_00479_),
    .Q(\u_async_wb.u_cmd_if.mem[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _09862_ (.CLK(clknet_leaf_45_wbm_clk_i),
    .D(_00480_),
    .Q(\u_async_wb.u_cmd_if.mem[3][32] ));
 sky130_fd_sc_hd__dfxtp_1 _09863_ (.CLK(clknet_leaf_45_wbm_clk_i),
    .D(_00481_),
    .Q(\u_async_wb.u_cmd_if.mem[3][33] ));
 sky130_fd_sc_hd__dfxtp_1 _09864_ (.CLK(clknet_leaf_45_wbm_clk_i),
    .D(_00482_),
    .Q(\u_async_wb.u_cmd_if.mem[3][34] ));
 sky130_fd_sc_hd__dfxtp_1 _09865_ (.CLK(clknet_leaf_45_wbm_clk_i),
    .D(_00483_),
    .Q(\u_async_wb.u_cmd_if.mem[3][35] ));
 sky130_fd_sc_hd__dfxtp_1 _09866_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00484_),
    .Q(\u_async_wb.u_cmd_if.mem[3][36] ));
 sky130_fd_sc_hd__dfxtp_1 _09867_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_00485_),
    .Q(\u_async_wb.u_cmd_if.mem[3][37] ));
 sky130_fd_sc_hd__dfxtp_1 _09868_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00486_),
    .Q(\u_async_wb.u_cmd_if.mem[3][38] ));
 sky130_fd_sc_hd__dfxtp_1 _09869_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00487_),
    .Q(\u_async_wb.u_cmd_if.mem[3][39] ));
 sky130_fd_sc_hd__dfxtp_1 _09870_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_00488_),
    .Q(\u_async_wb.u_cmd_if.mem[3][40] ));
 sky130_fd_sc_hd__dfxtp_1 _09871_ (.CLK(clknet_leaf_15_wbm_clk_i),
    .D(_00489_),
    .Q(\u_async_wb.u_cmd_if.mem[3][41] ));
 sky130_fd_sc_hd__dfxtp_1 _09872_ (.CLK(clknet_leaf_7_wbm_clk_i),
    .D(_00490_),
    .Q(\u_async_wb.u_cmd_if.mem[3][42] ));
 sky130_fd_sc_hd__dfxtp_1 _09873_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00491_),
    .Q(\u_async_wb.u_cmd_if.mem[3][43] ));
 sky130_fd_sc_hd__dfxtp_1 _09874_ (.CLK(clknet_leaf_7_wbm_clk_i),
    .D(_00492_),
    .Q(\u_async_wb.u_cmd_if.mem[3][44] ));
 sky130_fd_sc_hd__dfxtp_1 _09875_ (.CLK(clknet_leaf_6_wbm_clk_i),
    .D(_00493_),
    .Q(\u_async_wb.u_cmd_if.mem[3][45] ));
 sky130_fd_sc_hd__dfxtp_1 _09876_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00494_),
    .Q(\u_async_wb.u_cmd_if.mem[3][46] ));
 sky130_fd_sc_hd__dfxtp_1 _09877_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00495_),
    .Q(\u_async_wb.u_cmd_if.mem[3][47] ));
 sky130_fd_sc_hd__dfxtp_1 _09878_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00496_),
    .Q(\u_async_wb.u_cmd_if.mem[3][48] ));
 sky130_fd_sc_hd__dfxtp_1 _09879_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00497_),
    .Q(\u_async_wb.u_cmd_if.mem[3][49] ));
 sky130_fd_sc_hd__dfxtp_1 _09880_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00498_),
    .Q(\u_async_wb.u_cmd_if.mem[3][50] ));
 sky130_fd_sc_hd__dfxtp_1 _09881_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00499_),
    .Q(\u_async_wb.u_cmd_if.mem[3][51] ));
 sky130_fd_sc_hd__dfxtp_1 _09882_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00500_),
    .Q(\u_async_wb.u_cmd_if.mem[3][52] ));
 sky130_fd_sc_hd__dfxtp_1 _09883_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00501_),
    .Q(\u_async_wb.u_cmd_if.mem[3][53] ));
 sky130_fd_sc_hd__dfxtp_1 _09884_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00502_),
    .Q(\u_async_wb.u_cmd_if.mem[3][54] ));
 sky130_fd_sc_hd__dfxtp_1 _09885_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00503_),
    .Q(\u_async_wb.u_cmd_if.mem[3][55] ));
 sky130_fd_sc_hd__dfxtp_1 _09886_ (.CLK(clknet_leaf_22_wbm_clk_i),
    .D(_00504_),
    .Q(\u_async_wb.u_cmd_if.mem[3][56] ));
 sky130_fd_sc_hd__dfxtp_1 _09887_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00505_),
    .Q(\u_async_wb.u_cmd_if.mem[3][57] ));
 sky130_fd_sc_hd__dfxtp_1 _09888_ (.CLK(clknet_leaf_22_wbm_clk_i),
    .D(_00506_),
    .Q(\u_async_wb.u_cmd_if.mem[3][58] ));
 sky130_fd_sc_hd__dfxtp_1 _09889_ (.CLK(clknet_leaf_23_wbm_clk_i),
    .D(_00507_),
    .Q(\u_async_wb.u_cmd_if.mem[3][59] ));
 sky130_fd_sc_hd__dfxtp_1 _09890_ (.CLK(clknet_leaf_23_wbm_clk_i),
    .D(_00508_),
    .Q(\u_async_wb.u_cmd_if.mem[3][60] ));
 sky130_fd_sc_hd__dfxtp_1 _09891_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00509_),
    .Q(\u_async_wb.u_cmd_if.mem[3][61] ));
 sky130_fd_sc_hd__dfxtp_1 _09892_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00510_),
    .Q(\u_async_wb.u_cmd_if.mem[3][62] ));
 sky130_fd_sc_hd__dfxtp_1 _09893_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00511_),
    .Q(\u_async_wb.u_cmd_if.mem[3][63] ));
 sky130_fd_sc_hd__dfxtp_1 _09894_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00512_),
    .Q(\u_async_wb.u_cmd_if.mem[3][64] ));
 sky130_fd_sc_hd__dfxtp_1 _09895_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00513_),
    .Q(\u_async_wb.u_cmd_if.mem[3][65] ));
 sky130_fd_sc_hd__dfxtp_1 _09896_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00514_),
    .Q(\u_async_wb.u_cmd_if.mem[3][66] ));
 sky130_fd_sc_hd__dfxtp_1 _09897_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00515_),
    .Q(\u_async_wb.u_cmd_if.mem[3][67] ));
 sky130_fd_sc_hd__dfxtp_1 _09898_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00516_),
    .Q(\u_async_wb.u_cmd_if.mem[3][68] ));
 sky130_fd_sc_hd__dfrtp_1 _09899_ (.CLK(clknet_leaf_68_wbm_clk_i),
    .D(net316),
    .RESET_B(net304),
    .Q(\u_uart2wb.u_arst_sync.in_data_s ));
 sky130_fd_sc_hd__conb_1 _09899__316 (.HI(net316));
 sky130_fd_sc_hd__dfrtp_1 _09900_ (.CLK(clknet_leaf_68_wbm_clk_i),
    .D(net354),
    .RESET_B(net304),
    .Q(\u_uart2wb.u_arst_sync.in_data_2s ));
 sky130_fd_sc_hd__dfrtp_1 _09901_ (.CLK(clknet_leaf_91_wbm_clk_i),
    .D(net365),
    .RESET_B(net285),
    .Q(\u_uart2wb.u_async_reg_bus.in_flag_ss ));
 sky130_fd_sc_hd__dfrtp_1 _09902_ (.CLK(clknet_leaf_91_wbm_clk_i),
    .D(\u_uart2wb.u_async_reg_bus.in_flag ),
    .RESET_B(net285),
    .Q(\u_uart2wb.u_async_reg_bus.in_flag_s ));
 sky130_fd_sc_hd__dfxtp_1 _09903_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00517_),
    .Q(\u_async_wb.u_cmd_if.mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _09904_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00518_),
    .Q(\u_async_wb.u_cmd_if.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _09905_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00519_),
    .Q(\u_async_wb.u_cmd_if.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _09906_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00520_),
    .Q(\u_async_wb.u_cmd_if.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _09907_ (.CLK(clknet_leaf_43_wbm_clk_i),
    .D(_00521_),
    .Q(\u_async_wb.u_cmd_if.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _09908_ (.CLK(clknet_leaf_42_wbm_clk_i),
    .D(_00522_),
    .Q(\u_async_wb.u_cmd_if.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _09909_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00523_),
    .Q(\u_async_wb.u_cmd_if.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _09910_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00524_),
    .Q(\u_async_wb.u_cmd_if.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _09911_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00525_),
    .Q(\u_async_wb.u_cmd_if.mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _09912_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00526_),
    .Q(\u_async_wb.u_cmd_if.mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _09913_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00527_),
    .Q(\u_async_wb.u_cmd_if.mem[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _09914_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00528_),
    .Q(\u_async_wb.u_cmd_if.mem[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _09915_ (.CLK(clknet_leaf_29_wbm_clk_i),
    .D(_00529_),
    .Q(\u_async_wb.u_cmd_if.mem[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _09916_ (.CLK(clknet_leaf_29_wbm_clk_i),
    .D(_00530_),
    .Q(\u_async_wb.u_cmd_if.mem[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _09917_ (.CLK(clknet_leaf_29_wbm_clk_i),
    .D(_00531_),
    .Q(\u_async_wb.u_cmd_if.mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _09918_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00532_),
    .Q(\u_async_wb.u_cmd_if.mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _09919_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00533_),
    .Q(\u_async_wb.u_cmd_if.mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _09920_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00534_),
    .Q(\u_async_wb.u_cmd_if.mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _09921_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00535_),
    .Q(\u_async_wb.u_cmd_if.mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _09922_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00536_),
    .Q(\u_async_wb.u_cmd_if.mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _09923_ (.CLK(clknet_leaf_41_wbm_clk_i),
    .D(_00537_),
    .Q(\u_async_wb.u_cmd_if.mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _09924_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00538_),
    .Q(\u_async_wb.u_cmd_if.mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _09925_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00539_),
    .Q(\u_async_wb.u_cmd_if.mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _09926_ (.CLK(clknet_leaf_39_wbm_clk_i),
    .D(_00540_),
    .Q(\u_async_wb.u_cmd_if.mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _09927_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00541_),
    .Q(\u_async_wb.u_cmd_if.mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _09928_ (.CLK(clknet_leaf_41_wbm_clk_i),
    .D(_00542_),
    .Q(\u_async_wb.u_cmd_if.mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _09929_ (.CLK(clknet_leaf_43_wbm_clk_i),
    .D(_00543_),
    .Q(\u_async_wb.u_cmd_if.mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _09930_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00544_),
    .Q(\u_async_wb.u_cmd_if.mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _09931_ (.CLK(clknet_leaf_43_wbm_clk_i),
    .D(_00545_),
    .Q(\u_async_wb.u_cmd_if.mem[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _09932_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00546_),
    .Q(\u_async_wb.u_cmd_if.mem[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _09933_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00547_),
    .Q(\u_async_wb.u_cmd_if.mem[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _09934_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00548_),
    .Q(\u_async_wb.u_cmd_if.mem[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _09935_ (.CLK(clknet_leaf_46_wbm_clk_i),
    .D(_00549_),
    .Q(\u_async_wb.u_cmd_if.mem[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _09936_ (.CLK(clknet_leaf_45_wbm_clk_i),
    .D(_00550_),
    .Q(\u_async_wb.u_cmd_if.mem[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _09937_ (.CLK(clknet_leaf_45_wbm_clk_i),
    .D(_00551_),
    .Q(\u_async_wb.u_cmd_if.mem[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _09938_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00552_),
    .Q(\u_async_wb.u_cmd_if.mem[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _09939_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00553_),
    .Q(\u_async_wb.u_cmd_if.mem[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _09940_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00554_),
    .Q(\u_async_wb.u_cmd_if.mem[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _09941_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_00555_),
    .Q(\u_async_wb.u_cmd_if.mem[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _09942_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00556_),
    .Q(\u_async_wb.u_cmd_if.mem[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _09943_ (.CLK(clknet_leaf_15_wbm_clk_i),
    .D(_00557_),
    .Q(\u_async_wb.u_cmd_if.mem[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _09944_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00558_),
    .Q(\u_async_wb.u_cmd_if.mem[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _09945_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00559_),
    .Q(\u_async_wb.u_cmd_if.mem[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _09946_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00560_),
    .Q(\u_async_wb.u_cmd_if.mem[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _09947_ (.CLK(clknet_leaf_7_wbm_clk_i),
    .D(_00561_),
    .Q(\u_async_wb.u_cmd_if.mem[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _09948_ (.CLK(clknet_leaf_7_wbm_clk_i),
    .D(_00562_),
    .Q(\u_async_wb.u_cmd_if.mem[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _09949_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00563_),
    .Q(\u_async_wb.u_cmd_if.mem[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _09950_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00564_),
    .Q(\u_async_wb.u_cmd_if.mem[2][47] ));
 sky130_fd_sc_hd__dfxtp_1 _09951_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00565_),
    .Q(\u_async_wb.u_cmd_if.mem[2][48] ));
 sky130_fd_sc_hd__dfxtp_1 _09952_ (.CLK(clknet_leaf_4_wbm_clk_i),
    .D(_00566_),
    .Q(\u_async_wb.u_cmd_if.mem[2][49] ));
 sky130_fd_sc_hd__dfxtp_1 _09953_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00567_),
    .Q(\u_async_wb.u_cmd_if.mem[2][50] ));
 sky130_fd_sc_hd__dfxtp_1 _09954_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00568_),
    .Q(\u_async_wb.u_cmd_if.mem[2][51] ));
 sky130_fd_sc_hd__dfxtp_1 _09955_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00569_),
    .Q(\u_async_wb.u_cmd_if.mem[2][52] ));
 sky130_fd_sc_hd__dfxtp_1 _09956_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00570_),
    .Q(\u_async_wb.u_cmd_if.mem[2][53] ));
 sky130_fd_sc_hd__dfxtp_1 _09957_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00571_),
    .Q(\u_async_wb.u_cmd_if.mem[2][54] ));
 sky130_fd_sc_hd__dfxtp_1 _09958_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00572_),
    .Q(\u_async_wb.u_cmd_if.mem[2][55] ));
 sky130_fd_sc_hd__dfxtp_1 _09959_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00573_),
    .Q(\u_async_wb.u_cmd_if.mem[2][56] ));
 sky130_fd_sc_hd__dfxtp_1 _09960_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00574_),
    .Q(\u_async_wb.u_cmd_if.mem[2][57] ));
 sky130_fd_sc_hd__dfxtp_1 _09961_ (.CLK(clknet_leaf_22_wbm_clk_i),
    .D(_00575_),
    .Q(\u_async_wb.u_cmd_if.mem[2][58] ));
 sky130_fd_sc_hd__dfxtp_1 _09962_ (.CLK(clknet_leaf_22_wbm_clk_i),
    .D(_00576_),
    .Q(\u_async_wb.u_cmd_if.mem[2][59] ));
 sky130_fd_sc_hd__dfxtp_1 _09963_ (.CLK(clknet_leaf_23_wbm_clk_i),
    .D(_00577_),
    .Q(\u_async_wb.u_cmd_if.mem[2][60] ));
 sky130_fd_sc_hd__dfxtp_1 _09964_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00578_),
    .Q(\u_async_wb.u_cmd_if.mem[2][61] ));
 sky130_fd_sc_hd__dfxtp_1 _09965_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00579_),
    .Q(\u_async_wb.u_cmd_if.mem[2][62] ));
 sky130_fd_sc_hd__dfxtp_1 _09966_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00580_),
    .Q(\u_async_wb.u_cmd_if.mem[2][63] ));
 sky130_fd_sc_hd__dfxtp_1 _09967_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00581_),
    .Q(\u_async_wb.u_cmd_if.mem[2][64] ));
 sky130_fd_sc_hd__dfxtp_1 _09968_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00582_),
    .Q(\u_async_wb.u_cmd_if.mem[2][65] ));
 sky130_fd_sc_hd__dfxtp_1 _09969_ (.CLK(clknet_leaf_23_wbm_clk_i),
    .D(_00583_),
    .Q(\u_async_wb.u_cmd_if.mem[2][66] ));
 sky130_fd_sc_hd__dfxtp_1 _09970_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00584_),
    .Q(\u_async_wb.u_cmd_if.mem[2][67] ));
 sky130_fd_sc_hd__dfxtp_1 _09971_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00585_),
    .Q(\u_async_wb.u_cmd_if.mem[2][68] ));
 sky130_fd_sc_hd__dfxtp_1 _09972_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00586_),
    .Q(\u_async_wb.u_cmd_if.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _09973_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00587_),
    .Q(\u_async_wb.u_cmd_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _09974_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00588_),
    .Q(\u_async_wb.u_cmd_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _09975_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00589_),
    .Q(\u_async_wb.u_cmd_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _09976_ (.CLK(clknet_leaf_43_wbm_clk_i),
    .D(_00590_),
    .Q(\u_async_wb.u_cmd_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _09977_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00591_),
    .Q(\u_async_wb.u_cmd_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _09978_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00592_),
    .Q(\u_async_wb.u_cmd_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _09979_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00593_),
    .Q(\u_async_wb.u_cmd_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _09980_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00594_),
    .Q(\u_async_wb.u_cmd_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _09981_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00595_),
    .Q(\u_async_wb.u_cmd_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _09982_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00596_),
    .Q(\u_async_wb.u_cmd_if.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _09983_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00597_),
    .Q(\u_async_wb.u_cmd_if.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _09984_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00598_),
    .Q(\u_async_wb.u_cmd_if.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _09985_ (.CLK(clknet_leaf_29_wbm_clk_i),
    .D(_00599_),
    .Q(\u_async_wb.u_cmd_if.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _09986_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00600_),
    .Q(\u_async_wb.u_cmd_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _09987_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00601_),
    .Q(\u_async_wb.u_cmd_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _09988_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00602_),
    .Q(\u_async_wb.u_cmd_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _09989_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00603_),
    .Q(\u_async_wb.u_cmd_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _09990_ (.CLK(clknet_leaf_31_wbm_clk_i),
    .D(_00604_),
    .Q(\u_async_wb.u_cmd_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _09991_ (.CLK(clknet_leaf_41_wbm_clk_i),
    .D(_00605_),
    .Q(\u_async_wb.u_cmd_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _09992_ (.CLK(clknet_leaf_41_wbm_clk_i),
    .D(_00606_),
    .Q(\u_async_wb.u_cmd_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _09993_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00607_),
    .Q(\u_async_wb.u_cmd_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _09994_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00608_),
    .Q(\u_async_wb.u_cmd_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _09995_ (.CLK(clknet_leaf_39_wbm_clk_i),
    .D(_00609_),
    .Q(\u_async_wb.u_cmd_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _09996_ (.CLK(clknet_leaf_39_wbm_clk_i),
    .D(_00610_),
    .Q(\u_async_wb.u_cmd_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _09997_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00611_),
    .Q(\u_async_wb.u_cmd_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _09998_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00612_),
    .Q(\u_async_wb.u_cmd_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _09999_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00613_),
    .Q(\u_async_wb.u_cmd_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10000_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00614_),
    .Q(\u_async_wb.u_cmd_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10001_ (.CLK(clknet_leaf_48_wbm_clk_i),
    .D(_00615_),
    .Q(\u_async_wb.u_cmd_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10002_ (.CLK(clknet_leaf_47_wbm_clk_i),
    .D(_00616_),
    .Q(\u_async_wb.u_cmd_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _10003_ (.CLK(clknet_leaf_47_wbm_clk_i),
    .D(_00617_),
    .Q(\u_async_wb.u_cmd_if.mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _10004_ (.CLK(clknet_leaf_46_wbm_clk_i),
    .D(_00618_),
    .Q(\u_async_wb.u_cmd_if.mem[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _10005_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00619_),
    .Q(\u_async_wb.u_cmd_if.mem[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _10006_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00620_),
    .Q(\u_async_wb.u_cmd_if.mem[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _10007_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00621_),
    .Q(\u_async_wb.u_cmd_if.mem[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _10008_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00622_),
    .Q(\u_async_wb.u_cmd_if.mem[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _10009_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00623_),
    .Q(\u_async_wb.u_cmd_if.mem[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _10010_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00624_),
    .Q(\u_async_wb.u_cmd_if.mem[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _10011_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00625_),
    .Q(\u_async_wb.u_cmd_if.mem[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _10012_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_00626_),
    .Q(\u_async_wb.u_cmd_if.mem[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _10013_ (.CLK(clknet_leaf_15_wbm_clk_i),
    .D(_00627_),
    .Q(\u_async_wb.u_cmd_if.mem[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _10014_ (.CLK(clknet_leaf_15_wbm_clk_i),
    .D(_00628_),
    .Q(\u_async_wb.u_cmd_if.mem[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _10015_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00629_),
    .Q(\u_async_wb.u_cmd_if.mem[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _10016_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00630_),
    .Q(\u_async_wb.u_cmd_if.mem[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _10017_ (.CLK(clknet_leaf_7_wbm_clk_i),
    .D(_00631_),
    .Q(\u_async_wb.u_cmd_if.mem[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _10018_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00632_),
    .Q(\u_async_wb.u_cmd_if.mem[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _10019_ (.CLK(clknet_leaf_6_wbm_clk_i),
    .D(_00633_),
    .Q(\u_async_wb.u_cmd_if.mem[1][47] ));
 sky130_fd_sc_hd__dfxtp_1 _10020_ (.CLK(clknet_leaf_6_wbm_clk_i),
    .D(_00634_),
    .Q(\u_async_wb.u_cmd_if.mem[1][48] ));
 sky130_fd_sc_hd__dfxtp_1 _10021_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00635_),
    .Q(\u_async_wb.u_cmd_if.mem[1][49] ));
 sky130_fd_sc_hd__dfxtp_1 _10022_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00636_),
    .Q(\u_async_wb.u_cmd_if.mem[1][50] ));
 sky130_fd_sc_hd__dfxtp_1 _10023_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00637_),
    .Q(\u_async_wb.u_cmd_if.mem[1][51] ));
 sky130_fd_sc_hd__dfxtp_1 _10024_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00638_),
    .Q(\u_async_wb.u_cmd_if.mem[1][52] ));
 sky130_fd_sc_hd__dfxtp_1 _10025_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00639_),
    .Q(\u_async_wb.u_cmd_if.mem[1][53] ));
 sky130_fd_sc_hd__dfxtp_1 _10026_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00640_),
    .Q(\u_async_wb.u_cmd_if.mem[1][54] ));
 sky130_fd_sc_hd__dfxtp_1 _10027_ (.CLK(clknet_leaf_22_wbm_clk_i),
    .D(_00641_),
    .Q(\u_async_wb.u_cmd_if.mem[1][55] ));
 sky130_fd_sc_hd__dfxtp_1 _10028_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00642_),
    .Q(\u_async_wb.u_cmd_if.mem[1][56] ));
 sky130_fd_sc_hd__dfxtp_1 _10029_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00643_),
    .Q(\u_async_wb.u_cmd_if.mem[1][57] ));
 sky130_fd_sc_hd__dfxtp_1 _10030_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00644_),
    .Q(\u_async_wb.u_cmd_if.mem[1][58] ));
 sky130_fd_sc_hd__dfxtp_1 _10031_ (.CLK(clknet_leaf_23_wbm_clk_i),
    .D(_00645_),
    .Q(\u_async_wb.u_cmd_if.mem[1][59] ));
 sky130_fd_sc_hd__dfxtp_1 _10032_ (.CLK(clknet_leaf_23_wbm_clk_i),
    .D(_00646_),
    .Q(\u_async_wb.u_cmd_if.mem[1][60] ));
 sky130_fd_sc_hd__dfxtp_1 _10033_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00647_),
    .Q(\u_async_wb.u_cmd_if.mem[1][61] ));
 sky130_fd_sc_hd__dfxtp_1 _10034_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00648_),
    .Q(\u_async_wb.u_cmd_if.mem[1][62] ));
 sky130_fd_sc_hd__dfxtp_1 _10035_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00649_),
    .Q(\u_async_wb.u_cmd_if.mem[1][63] ));
 sky130_fd_sc_hd__dfxtp_1 _10036_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00650_),
    .Q(\u_async_wb.u_cmd_if.mem[1][64] ));
 sky130_fd_sc_hd__dfxtp_1 _10037_ (.CLK(clknet_leaf_23_wbm_clk_i),
    .D(_00651_),
    .Q(\u_async_wb.u_cmd_if.mem[1][65] ));
 sky130_fd_sc_hd__dfxtp_1 _10038_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00652_),
    .Q(\u_async_wb.u_cmd_if.mem[1][66] ));
 sky130_fd_sc_hd__dfxtp_1 _10039_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00653_),
    .Q(\u_async_wb.u_cmd_if.mem[1][67] ));
 sky130_fd_sc_hd__dfxtp_1 _10040_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00654_),
    .Q(\u_async_wb.u_cmd_if.mem[1][68] ));
 sky130_fd_sc_hd__dfxtp_1 _10041_ (.CLK(clknet_leaf_14_wbm_clk_i),
    .D(_00655_),
    .Q(\u_async_wb.u_cmd_if.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10042_ (.CLK(clknet_leaf_15_wbm_clk_i),
    .D(_00656_),
    .Q(\u_async_wb.u_cmd_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10043_ (.CLK(clknet_leaf_16_wbm_clk_i),
    .D(_00657_),
    .Q(\u_async_wb.u_cmd_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10044_ (.CLK(clknet_leaf_15_wbm_clk_i),
    .D(_00658_),
    .Q(\u_async_wb.u_cmd_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10045_ (.CLK(clknet_leaf_43_wbm_clk_i),
    .D(_00659_),
    .Q(\u_async_wb.u_cmd_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10046_ (.CLK(clknet_leaf_42_wbm_clk_i),
    .D(_00660_),
    .Q(\u_async_wb.u_cmd_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10047_ (.CLK(clknet_leaf_42_wbm_clk_i),
    .D(_00661_),
    .Q(\u_async_wb.u_cmd_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10048_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00662_),
    .Q(\u_async_wb.u_cmd_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10049_ (.CLK(clknet_leaf_42_wbm_clk_i),
    .D(_00663_),
    .Q(\u_async_wb.u_cmd_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10050_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00664_),
    .Q(\u_async_wb.u_cmd_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10051_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00665_),
    .Q(\u_async_wb.u_cmd_if.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10052_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00666_),
    .Q(\u_async_wb.u_cmd_if.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10053_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00667_),
    .Q(\u_async_wb.u_cmd_if.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10054_ (.CLK(clknet_leaf_28_wbm_clk_i),
    .D(_00668_),
    .Q(\u_async_wb.u_cmd_if.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10055_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00669_),
    .Q(\u_async_wb.u_cmd_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10056_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00670_),
    .Q(\u_async_wb.u_cmd_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10057_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00671_),
    .Q(\u_async_wb.u_cmd_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10058_ (.CLK(clknet_leaf_30_wbm_clk_i),
    .D(_00672_),
    .Q(\u_async_wb.u_cmd_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10059_ (.CLK(clknet_leaf_31_wbm_clk_i),
    .D(_00673_),
    .Q(\u_async_wb.u_cmd_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10060_ (.CLK(clknet_leaf_32_wbm_clk_i),
    .D(_00674_),
    .Q(\u_async_wb.u_cmd_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10061_ (.CLK(clknet_leaf_41_wbm_clk_i),
    .D(_00675_),
    .Q(\u_async_wb.u_cmd_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10062_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00676_),
    .Q(\u_async_wb.u_cmd_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10063_ (.CLK(clknet_leaf_40_wbm_clk_i),
    .D(_00677_),
    .Q(\u_async_wb.u_cmd_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10064_ (.CLK(clknet_leaf_39_wbm_clk_i),
    .D(_00678_),
    .Q(\u_async_wb.u_cmd_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10065_ (.CLK(clknet_leaf_50_wbm_clk_i),
    .D(_00679_),
    .Q(\u_async_wb.u_cmd_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10066_ (.CLK(clknet_leaf_41_wbm_clk_i),
    .D(_00680_),
    .Q(\u_async_wb.u_cmd_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10067_ (.CLK(clknet_leaf_43_wbm_clk_i),
    .D(_00681_),
    .Q(\u_async_wb.u_cmd_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10068_ (.CLK(clknet_leaf_48_wbm_clk_i),
    .D(_00682_),
    .Q(\u_async_wb.u_cmd_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10069_ (.CLK(clknet_leaf_44_wbm_clk_i),
    .D(_00683_),
    .Q(\u_async_wb.u_cmd_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10070_ (.CLK(clknet_leaf_48_wbm_clk_i),
    .D(_00684_),
    .Q(\u_async_wb.u_cmd_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10071_ (.CLK(clknet_leaf_47_wbm_clk_i),
    .D(_00685_),
    .Q(\u_async_wb.u_cmd_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _10072_ (.CLK(clknet_leaf_47_wbm_clk_i),
    .D(_00686_),
    .Q(\u_async_wb.u_cmd_if.mem[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _10073_ (.CLK(clknet_leaf_46_wbm_clk_i),
    .D(_00687_),
    .Q(\u_async_wb.u_cmd_if.mem[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _10074_ (.CLK(clknet_leaf_45_wbm_clk_i),
    .D(_00688_),
    .Q(\u_async_wb.u_cmd_if.mem[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _10075_ (.CLK(clknet_leaf_45_wbm_clk_i),
    .D(_00689_),
    .Q(\u_async_wb.u_cmd_if.mem[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _10076_ (.CLK(clknet_leaf_45_wbm_clk_i),
    .D(_00690_),
    .Q(\u_async_wb.u_cmd_if.mem[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _10077_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00691_),
    .Q(\u_async_wb.u_cmd_if.mem[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _10078_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00692_),
    .Q(\u_async_wb.u_cmd_if.mem[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _10079_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00693_),
    .Q(\u_async_wb.u_cmd_if.mem[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _10080_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_00694_),
    .Q(\u_async_wb.u_cmd_if.mem[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _10081_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_00695_),
    .Q(\u_async_wb.u_cmd_if.mem[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _10082_ (.CLK(clknet_leaf_15_wbm_clk_i),
    .D(_00696_),
    .Q(\u_async_wb.u_cmd_if.mem[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _10083_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_00697_),
    .Q(\u_async_wb.u_cmd_if.mem[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _10084_ (.CLK(clknet_leaf_15_wbm_clk_i),
    .D(_00698_),
    .Q(\u_async_wb.u_cmd_if.mem[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _10085_ (.CLK(clknet_leaf_7_wbm_clk_i),
    .D(_00699_),
    .Q(\u_async_wb.u_cmd_if.mem[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _10086_ (.CLK(clknet_leaf_8_wbm_clk_i),
    .D(_00700_),
    .Q(\u_async_wb.u_cmd_if.mem[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _10087_ (.CLK(clknet_leaf_19_wbm_clk_i),
    .D(_00701_),
    .Q(\u_async_wb.u_cmd_if.mem[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _10088_ (.CLK(clknet_leaf_6_wbm_clk_i),
    .D(_00702_),
    .Q(\u_async_wb.u_cmd_if.mem[0][47] ));
 sky130_fd_sc_hd__dfxtp_1 _10089_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00703_),
    .Q(\u_async_wb.u_cmd_if.mem[0][48] ));
 sky130_fd_sc_hd__dfxtp_1 _10090_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00704_),
    .Q(\u_async_wb.u_cmd_if.mem[0][49] ));
 sky130_fd_sc_hd__dfxtp_1 _10091_ (.CLK(clknet_leaf_5_wbm_clk_i),
    .D(_00705_),
    .Q(\u_async_wb.u_cmd_if.mem[0][50] ));
 sky130_fd_sc_hd__dfxtp_1 _10092_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00706_),
    .Q(\u_async_wb.u_cmd_if.mem[0][51] ));
 sky130_fd_sc_hd__dfxtp_1 _10093_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00707_),
    .Q(\u_async_wb.u_cmd_if.mem[0][52] ));
 sky130_fd_sc_hd__dfxtp_1 _10094_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00708_),
    .Q(\u_async_wb.u_cmd_if.mem[0][53] ));
 sky130_fd_sc_hd__dfxtp_1 _10095_ (.CLK(clknet_leaf_20_wbm_clk_i),
    .D(_00709_),
    .Q(\u_async_wb.u_cmd_if.mem[0][54] ));
 sky130_fd_sc_hd__dfxtp_1 _10096_ (.CLK(clknet_leaf_21_wbm_clk_i),
    .D(_00710_),
    .Q(\u_async_wb.u_cmd_if.mem[0][55] ));
 sky130_fd_sc_hd__dfxtp_1 _10097_ (.CLK(clknet_leaf_18_wbm_clk_i),
    .D(_00711_),
    .Q(\u_async_wb.u_cmd_if.mem[0][56] ));
 sky130_fd_sc_hd__dfxtp_1 _10098_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00712_),
    .Q(\u_async_wb.u_cmd_if.mem[0][57] ));
 sky130_fd_sc_hd__dfxtp_1 _10099_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00713_),
    .Q(\u_async_wb.u_cmd_if.mem[0][58] ));
 sky130_fd_sc_hd__dfxtp_1 _10100_ (.CLK(clknet_leaf_22_wbm_clk_i),
    .D(_00714_),
    .Q(\u_async_wb.u_cmd_if.mem[0][59] ));
 sky130_fd_sc_hd__dfxtp_1 _10101_ (.CLK(clknet_leaf_28_wbm_clk_i),
    .D(_00715_),
    .Q(\u_async_wb.u_cmd_if.mem[0][60] ));
 sky130_fd_sc_hd__dfxtp_1 _10102_ (.CLK(clknet_leaf_27_wbm_clk_i),
    .D(_00716_),
    .Q(\u_async_wb.u_cmd_if.mem[0][61] ));
 sky130_fd_sc_hd__dfxtp_1 _10103_ (.CLK(clknet_leaf_28_wbm_clk_i),
    .D(_00717_),
    .Q(\u_async_wb.u_cmd_if.mem[0][62] ));
 sky130_fd_sc_hd__dfxtp_1 _10104_ (.CLK(clknet_leaf_26_wbm_clk_i),
    .D(_00718_),
    .Q(\u_async_wb.u_cmd_if.mem[0][63] ));
 sky130_fd_sc_hd__dfxtp_1 _10105_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00719_),
    .Q(\u_async_wb.u_cmd_if.mem[0][64] ));
 sky130_fd_sc_hd__dfxtp_1 _10106_ (.CLK(clknet_leaf_24_wbm_clk_i),
    .D(_00720_),
    .Q(\u_async_wb.u_cmd_if.mem[0][65] ));
 sky130_fd_sc_hd__dfxtp_1 _10107_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00721_),
    .Q(\u_async_wb.u_cmd_if.mem[0][66] ));
 sky130_fd_sc_hd__dfxtp_1 _10108_ (.CLK(clknet_leaf_25_wbm_clk_i),
    .D(_00722_),
    .Q(\u_async_wb.u_cmd_if.mem[0][67] ));
 sky130_fd_sc_hd__dfxtp_1 _10109_ (.CLK(clknet_leaf_17_wbm_clk_i),
    .D(_00723_),
    .Q(\u_async_wb.u_cmd_if.mem[0][68] ));
 sky130_fd_sc_hd__dfxtp_1 _10110_ (.CLK(clknet_leaf_36_wbm_clk_i),
    .D(_00724_),
    .Q(net1));
 sky130_fd_sc_hd__dfxtp_1 _10111_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00725_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _10112_ (.CLK(clknet_leaf_36_wbm_clk_i),
    .D(_00726_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _10113_ (.CLK(clknet_leaf_34_wbm_clk_i),
    .D(_00727_),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_1 _10114_ (.CLK(clknet_leaf_36_wbm_clk_i),
    .D(_00728_),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _10115_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00729_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _10116_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00730_),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_1 _10117_ (.CLK(clknet_leaf_69_wbm_clk_i),
    .D(_00731_),
    .RESET_B(net270),
    .Q(\u_spi2wb.u_if.bitcnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10118_ (.CLK(clknet_leaf_67_wbm_clk_i),
    .D(_00732_),
    .RESET_B(net271),
    .Q(\u_spi2wb.u_if.bitcnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10119_ (.CLK(clknet_leaf_69_wbm_clk_i),
    .D(_00733_),
    .RESET_B(net270),
    .Q(\u_spi2wb.u_if.bitcnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10120_ (.CLK(clknet_leaf_73_wbm_clk_i),
    .D(_00734_),
    .RESET_B(net271),
    .Q(\u_spi2wb.u_if.bitcnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10121_ (.CLK(clknet_leaf_73_wbm_clk_i),
    .D(_00735_),
    .RESET_B(net275),
    .Q(\u_spi2wb.u_if.bitcnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10122_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(_00736_),
    .RESET_B(net275),
    .Q(\u_spi2wb.u_if.bitcnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10123_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00737_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10124_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00738_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10125_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00739_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10126_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00740_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10127_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00741_),
    .RESET_B(net241),
    .Q(\u_uart2wb.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10128_ (.CLK(\clknet_leaf_7_u_uart2wb.baud_clk_16x ),
    .D(_00742_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10129_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00743_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10130_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00744_),
    .RESET_B(net241),
    .Q(\u_uart2wb.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10131_ (.CLK(\clknet_leaf_7_u_uart2wb.baud_clk_16x ),
    .D(_00745_),
    .RESET_B(net241),
    .Q(\u_uart2wb.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10132_ (.CLK(\clknet_leaf_7_u_uart2wb.baud_clk_16x ),
    .D(_00746_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10133_ (.CLK(\clknet_leaf_7_u_uart2wb.baud_clk_16x ),
    .D(_00747_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10134_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00748_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10135_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00749_),
    .RESET_B(net242),
    .Q(\u_uart2wb.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10136_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00750_),
    .RESET_B(net242),
    .Q(\u_uart2wb.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10137_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00751_),
    .RESET_B(net240),
    .Q(\u_uart2wb.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10138_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_00752_),
    .RESET_B(net242),
    .Q(\u_uart2wb.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10139_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_00753_),
    .RESET_B(net245),
    .Q(\u_uart2wb.reg_rdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10140_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_00754_),
    .RESET_B(net245),
    .Q(\u_uart2wb.reg_rdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10141_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_00755_),
    .RESET_B(net245),
    .Q(\u_uart2wb.reg_rdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10142_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_00756_),
    .RESET_B(net245),
    .Q(\u_uart2wb.reg_rdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10143_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00757_),
    .RESET_B(net245),
    .Q(\u_uart2wb.reg_rdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10144_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00758_),
    .RESET_B(net245),
    .Q(\u_uart2wb.reg_rdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10145_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00759_),
    .RESET_B(net245),
    .Q(\u_uart2wb.reg_rdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10146_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00760_),
    .RESET_B(net245),
    .Q(\u_uart2wb.reg_rdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10147_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00761_),
    .RESET_B(net249),
    .Q(\u_uart2wb.reg_rdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10148_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00762_),
    .RESET_B(net249),
    .Q(\u_uart2wb.reg_rdata[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10149_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00763_),
    .RESET_B(net249),
    .Q(\u_uart2wb.reg_rdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10150_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00764_),
    .RESET_B(net249),
    .Q(\u_uart2wb.reg_rdata[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10151_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00765_),
    .RESET_B(net249),
    .Q(\u_uart2wb.reg_rdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10152_ (.CLK(\clknet_leaf_12_u_uart2wb.baud_clk_16x ),
    .D(_00766_),
    .RESET_B(net249),
    .Q(\u_uart2wb.reg_rdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10153_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(_00767_),
    .RESET_B(net249),
    .Q(\u_uart2wb.reg_rdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10154_ (.CLK(\clknet_leaf_12_u_uart2wb.baud_clk_16x ),
    .D(_00768_),
    .RESET_B(net249),
    .Q(\u_uart2wb.reg_rdata[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10155_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(_00769_),
    .RESET_B(net239),
    .Q(\u_uart2wb.reg_ack ));
 sky130_fd_sc_hd__dfrtp_1 _10156_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(_00770_),
    .RESET_B(net242),
    .Q(\u_uart2wb.u_async_reg_bus.in_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10157_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00771_),
    .RESET_B(net241),
    .Q(\u_uart2wb.u_async_reg_bus.in_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10158_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_00772_),
    .RESET_B(net237),
    .Q(\u_uart2wb.u_async_reg_bus.in_timer[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10159_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_00773_),
    .RESET_B(net237),
    .Q(\u_uart2wb.u_async_reg_bus.in_timer[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10160_ (.CLK(\clknet_leaf_24_u_uart2wb.baud_clk_16x ),
    .D(_00774_),
    .RESET_B(net237),
    .Q(\u_uart2wb.u_async_reg_bus.in_timer[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10161_ (.CLK(\clknet_leaf_24_u_uart2wb.baud_clk_16x ),
    .D(_00775_),
    .RESET_B(net237),
    .Q(\u_uart2wb.u_async_reg_bus.in_timer[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10162_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(_00776_),
    .RESET_B(net237),
    .Q(\u_uart2wb.u_async_reg_bus.in_timer[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10163_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(_00777_),
    .RESET_B(net237),
    .Q(\u_uart2wb.u_async_reg_bus.in_timer[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10164_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(_00778_),
    .RESET_B(net237),
    .Q(\u_uart2wb.u_async_reg_bus.in_timer[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10165_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00779_),
    .RESET_B(net241),
    .Q(\u_uart2wb.u_async_reg_bus.in_timer[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10166_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_00780_),
    .RESET_B(net241),
    .Q(\u_uart2wb.u_async_reg_bus.in_timer[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10167_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_00781_),
    .RESET_B(net239),
    .Q(\u_uart2wb.u_async_reg_bus.in_flag ));
 sky130_fd_sc_hd__dfrtp_1 _10168_ (.CLK(clknet_leaf_92_wbm_clk_i),
    .D(_00782_),
    .RESET_B(net285),
    .Q(\u_uart2wb.u_async_reg_bus.out_reg_cs ));
 sky130_fd_sc_hd__dfrtp_1 _10169_ (.CLK(clknet_leaf_92_wbm_clk_i),
    .D(_00783_),
    .RESET_B(net285),
    .Q(\u_uart2wb.u_async_reg_bus.out_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10170_ (.CLK(clknet_leaf_92_wbm_clk_i),
    .D(_00784_),
    .RESET_B(net285),
    .Q(\u_uart2wb.u_async_reg_bus.out_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10171_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(\u_uart2wb.u_async_reg_bus.out_flag ),
    .RESET_B(net232),
    .Q(\u_uart2wb.u_async_reg_bus.out_flag_s ));
 sky130_fd_sc_hd__dfrtp_1 _10172_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(net360),
    .RESET_B(net241),
    .Q(\u_uart2wb.u_async_reg_bus.out_flag_ss ));
 sky130_fd_sc_hd__dfrtp_2 _10173_ (.CLK(clknet_leaf_75_wbm_clk_i),
    .D(_00785_),
    .RESET_B(net278),
    .Q(\u_uart2wb.auto_rx_enb ));
 sky130_fd_sc_hd__dfrtp_1 _10174_ (.CLK(clknet_leaf_64_wbm_clk_i),
    .D(_00786_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10175_ (.CLK(clknet_leaf_64_wbm_clk_i),
    .D(_00787_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10176_ (.CLK(clknet_leaf_64_wbm_clk_i),
    .D(_00788_),
    .RESET_B(net282),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10177_ (.CLK(clknet_leaf_65_wbm_clk_i),
    .D(_00789_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10178_ (.CLK(clknet_leaf_79_wbm_clk_i),
    .D(_00790_),
    .RESET_B(net280),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10179_ (.CLK(clknet_leaf_65_wbm_clk_i),
    .D(_00791_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10180_ (.CLK(clknet_leaf_79_wbm_clk_i),
    .D(_00792_),
    .RESET_B(net283),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10181_ (.CLK(clknet_leaf_78_wbm_clk_i),
    .D(_00793_),
    .RESET_B(net280),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10182_ (.CLK(clknet_leaf_80_wbm_clk_i),
    .D(_00794_),
    .RESET_B(net277),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10183_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00795_),
    .RESET_B(net277),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10184_ (.CLK(clknet_leaf_81_wbm_clk_i),
    .D(_00796_),
    .RESET_B(net277),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10185_ (.CLK(clknet_leaf_81_wbm_clk_i),
    .D(_00797_),
    .RESET_B(net276),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10186_ (.CLK(clknet_leaf_81_wbm_clk_i),
    .D(_00798_),
    .RESET_B(net277),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10187_ (.CLK(clknet_leaf_75_wbm_clk_i),
    .D(_00799_),
    .RESET_B(net278),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10188_ (.CLK(clknet_leaf_75_wbm_clk_i),
    .D(_00800_),
    .RESET_B(net278),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10189_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(_00801_),
    .RESET_B(net280),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10190_ (.CLK(clknet_leaf_78_wbm_clk_i),
    .D(_00802_),
    .RESET_B(net280),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10191_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(_00803_),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10192_ (.CLK(clknet_leaf_78_wbm_clk_i),
    .D(_00804_),
    .RESET_B(net280),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10193_ (.CLK(clknet_leaf_78_wbm_clk_i),
    .D(_00805_),
    .RESET_B(net283),
    .Q(\u_uart2wb.u_aut_det.ref1_cnt[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10194_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(uartm_rxd),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.rxd_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10195_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(net355),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.rxd_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10196_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(\u_uart2wb.u_aut_det.rxd_sync[1] ),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.rxd_sync[2] ));
 sky130_fd_sc_hd__dfstp_1 _10197_ (.CLK(clknet_leaf_78_wbm_clk_i),
    .D(_00008_),
    .SET_B(net280),
    .Q(\u_uart2wb.u_aut_det.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10198_ (.CLK(clknet_leaf_77_wbm_clk_i),
    .D(_00009_),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10199_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(_00010_),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10200_ (.CLK(clknet_leaf_77_wbm_clk_i),
    .D(_00011_),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10201_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(_00012_),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10202_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(_00001_),
    .RESET_B(net280),
    .Q(\u_uart2wb.u_aut_det.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10203_ (.CLK(clknet_leaf_77_wbm_clk_i),
    .D(_00013_),
    .RESET_B(net284),
    .Q(\u_uart2wb.u_aut_det.state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10204_ (.CLK(clknet_leaf_75_wbm_clk_i),
    .D(_00014_),
    .RESET_B(net278),
    .Q(\u_uart2wb.u_aut_det.state[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10205_ (.CLK(clknet_leaf_92_wbm_clk_i),
    .D(_00806_),
    .RESET_B(net285),
    .Q(\u_uart2wb.u_async_reg_bus.out_flag ));
 sky130_fd_sc_hd__dfrtp_1 _10206_ (.CLK(clknet_leaf_68_wbm_clk_i),
    .D(_00807_),
    .RESET_B(net282),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10207_ (.CLK(clknet_leaf_66_wbm_clk_i),
    .D(_00808_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10208_ (.CLK(clknet_leaf_64_wbm_clk_i),
    .D(_00809_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10209_ (.CLK(clknet_leaf_66_wbm_clk_i),
    .D(_00810_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10210_ (.CLK(clknet_leaf_65_wbm_clk_i),
    .D(_00811_),
    .RESET_B(net282),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10211_ (.CLK(clknet_leaf_65_wbm_clk_i),
    .D(_00812_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10212_ (.CLK(clknet_leaf_65_wbm_clk_i),
    .D(_00813_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10213_ (.CLK(clknet_leaf_65_wbm_clk_i),
    .D(_00814_),
    .RESET_B(net281),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10214_ (.CLK(clknet_leaf_65_wbm_clk_i),
    .D(_00815_),
    .RESET_B(net282),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10215_ (.CLK(clknet_leaf_79_wbm_clk_i),
    .D(_00816_),
    .RESET_B(net280),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10216_ (.CLK(clknet_leaf_67_wbm_clk_i),
    .D(_00817_),
    .RESET_B(net282),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10217_ (.CLK(clknet_leaf_79_wbm_clk_i),
    .D(_00818_),
    .RESET_B(net283),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10218_ (.CLK(clknet_leaf_77_wbm_clk_i),
    .D(_00819_),
    .RESET_B(net280),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10219_ (.CLK(clknet_leaf_67_wbm_clk_i),
    .D(_00820_),
    .RESET_B(net284),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10220_ (.CLK(clknet_leaf_67_wbm_clk_i),
    .D(_00821_),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10221_ (.CLK(clknet_leaf_67_wbm_clk_i),
    .D(_00822_),
    .RESET_B(net282),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10222_ (.CLK(clknet_leaf_67_wbm_clk_i),
    .D(_00823_),
    .RESET_B(net279),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10223_ (.CLK(clknet_leaf_66_wbm_clk_i),
    .D(_00824_),
    .RESET_B(net282),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10224_ (.CLK(clknet_leaf_66_wbm_clk_i),
    .D(_00825_),
    .RESET_B(net282),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10225_ (.CLK(clknet_leaf_66_wbm_clk_i),
    .D(_00826_),
    .RESET_B(net282),
    .Q(\u_uart2wb.u_aut_det.clk_cnt[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10226_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00827_),
    .RESET_B(net276),
    .Q(\u_uart2wb.auto_baud_16x[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10227_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00828_),
    .RESET_B(net277),
    .Q(\u_uart2wb.auto_baud_16x[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10228_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00829_),
    .RESET_B(net276),
    .Q(\u_uart2wb.auto_baud_16x[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10229_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00830_),
    .RESET_B(net277),
    .Q(\u_uart2wb.auto_baud_16x[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10230_ (.CLK(clknet_leaf_82_wbm_clk_i),
    .D(_00831_),
    .RESET_B(net276),
    .Q(\u_uart2wb.auto_baud_16x[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10231_ (.CLK(clknet_leaf_82_wbm_clk_i),
    .D(_00832_),
    .RESET_B(net276),
    .Q(\u_uart2wb.auto_baud_16x[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10232_ (.CLK(clknet_leaf_82_wbm_clk_i),
    .D(_00833_),
    .RESET_B(net277),
    .Q(\u_uart2wb.auto_baud_16x[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10233_ (.CLK(clknet_leaf_82_wbm_clk_i),
    .D(_00834_),
    .RESET_B(net276),
    .Q(\u_uart2wb.auto_baud_16x[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10234_ (.CLK(clknet_leaf_82_wbm_clk_i),
    .D(_00835_),
    .RESET_B(net276),
    .Q(\u_uart2wb.auto_baud_16x[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10235_ (.CLK(clknet_leaf_87_wbm_clk_i),
    .D(_00836_),
    .RESET_B(net276),
    .Q(\u_uart2wb.auto_baud_16x[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10236_ (.CLK(clknet_leaf_87_wbm_clk_i),
    .D(_00837_),
    .RESET_B(net276),
    .Q(\u_uart2wb.auto_baud_16x[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10237_ (.CLK(clknet_leaf_82_wbm_clk_i),
    .D(_00838_),
    .RESET_B(net276),
    .Q(\u_uart2wb.auto_baud_16x[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10238_ (.CLK(\clknet_leaf_12_u_uart2wb.baud_clk_16x ),
    .D(_00032_),
    .RESET_B(net250),
    .Q(\u_uart2wb.u_core.u_txfsm.divcnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10239_ (.CLK(\clknet_leaf_12_u_uart2wb.baud_clk_16x ),
    .D(_00033_),
    .RESET_B(net250),
    .Q(\u_uart2wb.u_core.u_txfsm.divcnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10240_ (.CLK(\clknet_leaf_12_u_uart2wb.baud_clk_16x ),
    .D(_00034_),
    .RESET_B(net249),
    .Q(\u_uart2wb.u_core.u_txfsm.divcnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10241_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_00035_),
    .RESET_B(net250),
    .Q(\u_uart2wb.u_core.u_txfsm.divcnt[3] ));
 sky130_fd_sc_hd__dfstp_2 _10242_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00839_),
    .SET_B(net246),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _10243_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_00840_),
    .RESET_B(net248),
    .Q(\u_uart2wb.tx_rd ));
 sky130_fd_sc_hd__dfrtp_1 _10244_ (.CLK(\clknet_leaf_21_u_uart2wb.baud_clk_16x ),
    .D(_00841_),
    .RESET_B(net244),
    .Q(\u_uart2wb.u_core.u_rxfsm.rxstate[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10245_ (.CLK(\clknet_leaf_21_u_uart2wb.baud_clk_16x ),
    .D(_00842_),
    .RESET_B(net243),
    .Q(\u_uart2wb.u_core.u_rxfsm.rxstate[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10246_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00843_),
    .RESET_B(net244),
    .Q(\u_uart2wb.u_core.u_rxfsm.rxstate[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10247_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00844_),
    .RESET_B(net244),
    .Q(\u_uart2wb.u_core.u_rxfsm.rxpos[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10248_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00845_),
    .RESET_B(net243),
    .Q(\u_uart2wb.u_core.u_rxfsm.rxpos[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10249_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00846_),
    .RESET_B(net248),
    .Q(\u_uart2wb.u_core.u_rxfsm.rxpos[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10250_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00847_),
    .RESET_B(net248),
    .Q(\u_uart2wb.u_core.u_rxfsm.rxpos[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10251_ (.CLK(\clknet_leaf_21_u_uart2wb.baud_clk_16x ),
    .D(_00848_),
    .RESET_B(net243),
    .Q(\u_uart2wb.rx_wr ));
 sky130_fd_sc_hd__dfrtp_1 _10252_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00028_),
    .RESET_B(net244),
    .Q(\u_uart2wb.u_core.u_rxfsm.offset[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10253_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00029_),
    .RESET_B(net244),
    .Q(\u_uart2wb.u_core.u_rxfsm.offset[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10254_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00030_),
    .RESET_B(net248),
    .Q(\u_uart2wb.u_core.u_rxfsm.offset[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10255_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00031_),
    .RESET_B(net248),
    .Q(\u_uart2wb.u_core.u_rxfsm.offset[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10256_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_00849_),
    .RESET_B(net238),
    .Q(\u_uart2wb.u_core.u_rxfsm.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10257_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_00850_),
    .RESET_B(net238),
    .Q(\u_uart2wb.u_core.u_rxfsm.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10258_ (.CLK(\clknet_leaf_21_u_uart2wb.baud_clk_16x ),
    .D(_00851_),
    .RESET_B(net243),
    .Q(\u_uart2wb.u_core.u_rxfsm.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10259_ (.CLK(\clknet_leaf_24_u_uart2wb.baud_clk_16x ),
    .D(_00852_),
    .RESET_B(net238),
    .Q(\u_uart2wb.rx_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10260_ (.CLK(\clknet_leaf_24_u_uart2wb.baud_clk_16x ),
    .D(_00853_),
    .RESET_B(net238),
    .Q(\u_uart2wb.rx_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10261_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_00854_),
    .RESET_B(net238),
    .Q(\u_uart2wb.rx_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10262_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_00855_),
    .RESET_B(net237),
    .Q(\u_uart2wb.rx_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10263_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_00856_),
    .RESET_B(net238),
    .Q(\u_uart2wb.rx_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10264_ (.CLK(\clknet_leaf_24_u_uart2wb.baud_clk_16x ),
    .D(_00857_),
    .RESET_B(net238),
    .Q(\u_uart2wb.rx_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10265_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_00858_),
    .RESET_B(net238),
    .Q(\u_uart2wb.rx_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10266_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_00859_),
    .RESET_B(net237),
    .Q(\u_uart2wb.rx_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10267_ (.CLK(clknet_leaf_82_wbm_clk_i),
    .D(_00860_),
    .RESET_B(net299),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10268_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00861_),
    .RESET_B(net299),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10269_ (.CLK(clknet_leaf_82_wbm_clk_i),
    .D(_00862_),
    .RESET_B(net299),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10270_ (.CLK(clknet_leaf_85_wbm_clk_i),
    .D(_00863_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10271_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00864_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10272_ (.CLK(clknet_leaf_85_wbm_clk_i),
    .D(_00865_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10273_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00866_),
    .RESET_B(net297),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10274_ (.CLK(clknet_leaf_86_wbm_clk_i),
    .D(_00867_),
    .RESET_B(net298),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10275_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00868_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10276_ (.CLK(clknet_leaf_85_wbm_clk_i),
    .D(_00869_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10277_ (.CLK(clknet_leaf_86_wbm_clk_i),
    .D(_00870_),
    .RESET_B(net298),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10278_ (.CLK(clknet_leaf_85_wbm_clk_i),
    .D(_00871_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.low_count[11] ));
 sky130_fd_sc_hd__dfstp_1 _10279_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(net345),
    .SET_B(net246),
    .Q(\u_uart2wb.u_core.si_ss ));
 sky130_fd_sc_hd__dfstp_1 _10280_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(net366),
    .SET_B(net246),
    .Q(\u_uart2wb.u_core.u_rxd_sync.in_data_2s ));
 sky130_fd_sc_hd__dfstp_1 _10281_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(uartm_rxd),
    .SET_B(net247),
    .Q(\u_uart2wb.u_core.u_rxd_sync.in_data_s ));
 sky130_fd_sc_hd__dfrtp_1 _10282_ (.CLK(\clknet_leaf_12_u_uart2wb.baud_clk_16x ),
    .D(net359),
    .RESET_B(net300),
    .Q(\u_uart2wb.u_core.u_line_rst.in_data_2s ));
 sky130_fd_sc_hd__dfrtp_1 _10283_ (.CLK(\clknet_leaf_11_u_uart2wb.baud_clk_16x ),
    .D(net315),
    .RESET_B(net301),
    .Q(\u_uart2wb.u_core.u_line_rst.in_data_s ));
 sky130_fd_sc_hd__conb_1 _10283__315 (.HI(net315));
 sky130_fd_sc_hd__dfrtp_1 _10284_ (.CLK(clknet_leaf_86_wbm_clk_i),
    .D(_00021_),
    .RESET_B(net298),
    .Q(\u_uart2wb.u_core.line_clk_16x ));
 sky130_fd_sc_hd__dfrtp_1 _10285_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00872_),
    .RESET_B(net297),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10286_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00873_),
    .RESET_B(net299),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10287_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00874_),
    .RESET_B(net299),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10288_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00875_),
    .RESET_B(net299),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10289_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00876_),
    .RESET_B(net297),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10290_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00877_),
    .RESET_B(net297),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10291_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00878_),
    .RESET_B(net297),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10292_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00879_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10293_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00880_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10294_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00881_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10295_ (.CLK(clknet_leaf_84_wbm_clk_i),
    .D(_00882_),
    .RESET_B(net296),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10296_ (.CLK(clknet_leaf_85_wbm_clk_i),
    .D(_00883_),
    .RESET_B(net298),
    .Q(\u_uart2wb.u_core.u_clk_ctl.high_count[11] ));
 sky130_fd_sc_hd__dfxtp_1 _10297_ (.CLK(clknet_leaf_64_wbm_clk_i),
    .D(_00884_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _10298_ (.CLK(clknet_leaf_64_wbm_clk_i),
    .D(_00885_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10299_ (.CLK(clknet_leaf_64_wbm_clk_i),
    .D(_00886_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10300_ (.CLK(clknet_leaf_64_wbm_clk_i),
    .D(_00887_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _10301_ (.CLK(clknet_leaf_79_wbm_clk_i),
    .D(_00888_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _10302_ (.CLK(clknet_leaf_79_wbm_clk_i),
    .D(_00889_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _10303_ (.CLK(clknet_leaf_79_wbm_clk_i),
    .D(_00890_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 _10304_ (.CLK(clknet_leaf_79_wbm_clk_i),
    .D(_00891_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 _10305_ (.CLK(clknet_leaf_80_wbm_clk_i),
    .D(_00892_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[8] ));
 sky130_fd_sc_hd__dfxtp_1 _10306_ (.CLK(clknet_leaf_83_wbm_clk_i),
    .D(_00893_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[9] ));
 sky130_fd_sc_hd__dfxtp_1 _10307_ (.CLK(clknet_leaf_81_wbm_clk_i),
    .D(_00894_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[10] ));
 sky130_fd_sc_hd__dfxtp_1 _10308_ (.CLK(clknet_leaf_82_wbm_clk_i),
    .D(_00895_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[11] ));
 sky130_fd_sc_hd__dfxtp_2 _10309_ (.CLK(clknet_leaf_81_wbm_clk_i),
    .D(_00896_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[12] ));
 sky130_fd_sc_hd__dfxtp_1 _10310_ (.CLK(clknet_leaf_75_wbm_clk_i),
    .D(_00897_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[13] ));
 sky130_fd_sc_hd__dfxtp_1 _10311_ (.CLK(clknet_leaf_75_wbm_clk_i),
    .D(_00898_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[14] ));
 sky130_fd_sc_hd__dfxtp_1 _10312_ (.CLK(clknet_leaf_75_wbm_clk_i),
    .D(_00899_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[15] ));
 sky130_fd_sc_hd__dfxtp_1 _10313_ (.CLK(clknet_leaf_78_wbm_clk_i),
    .D(_00900_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[16] ));
 sky130_fd_sc_hd__dfxtp_1 _10314_ (.CLK(clknet_leaf_76_wbm_clk_i),
    .D(_00901_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[17] ));
 sky130_fd_sc_hd__dfxtp_1 _10315_ (.CLK(clknet_leaf_78_wbm_clk_i),
    .D(_00902_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[18] ));
 sky130_fd_sc_hd__dfxtp_1 _10316_ (.CLK(clknet_leaf_78_wbm_clk_i),
    .D(_00903_),
    .Q(\u_uart2wb.u_aut_det.ref2_cnt[19] ));
 sky130_fd_sc_hd__dfxtp_1 _10317_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_00904_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[5] ));
 sky130_fd_sc_hd__dfxtp_1 _10318_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_00905_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[13] ));
 sky130_fd_sc_hd__dfxtp_1 _10319_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00906_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[18] ));
 sky130_fd_sc_hd__dfxtp_1 _10320_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00907_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[17] ));
 sky130_fd_sc_hd__dfxtp_1 _10321_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00908_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[20] ));
 sky130_fd_sc_hd__dfxtp_1 _10322_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_00909_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[21] ));
 sky130_fd_sc_hd__dfxtp_1 _10323_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00910_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[12] ));
 sky130_fd_sc_hd__dfxtp_1 _10324_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_00911_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[24] ));
 sky130_fd_sc_hd__dfxtp_1 _10325_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00912_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[26] ));
 sky130_fd_sc_hd__dfxtp_1 _10326_ (.CLK(\clknet_leaf_19_u_uart2wb.baud_clk_16x ),
    .D(_00913_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[25] ));
 sky130_fd_sc_hd__dfxtp_1 _10327_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00914_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[28] ));
 sky130_fd_sc_hd__dfxtp_1 _10328_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_00915_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[29] ));
 sky130_fd_sc_hd__dfxtp_1 _10329_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00916_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[11] ));
 sky130_fd_sc_hd__dfxtp_1 _10330_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00917_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[32] ));
 sky130_fd_sc_hd__dfxtp_1 _10331_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00918_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[33] ));
 sky130_fd_sc_hd__dfxtp_1 _10332_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00919_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[34] ));
 sky130_fd_sc_hd__dfxtp_1 _10333_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00920_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[35] ));
 sky130_fd_sc_hd__dfxtp_1 _10334_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_00921_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[36] ));
 sky130_fd_sc_hd__dfxtp_1 _10335_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_00922_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[37] ));
 sky130_fd_sc_hd__dfxtp_1 _10336_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00923_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[38] ));
 sky130_fd_sc_hd__dfxtp_1 _10337_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00924_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[40] ));
 sky130_fd_sc_hd__dfxtp_1 _10338_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_00925_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[41] ));
 sky130_fd_sc_hd__dfxtp_1 _10339_ (.CLK(\clknet_leaf_20_u_uart2wb.baud_clk_16x ),
    .D(_00926_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[42] ));
 sky130_fd_sc_hd__dfxtp_1 _10340_ (.CLK(\clknet_leaf_18_u_uart2wb.baud_clk_16x ),
    .D(_00927_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[43] ));
 sky130_fd_sc_hd__dfxtp_1 _10341_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_00928_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[44] ));
 sky130_fd_sc_hd__dfxtp_1 _10342_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_00929_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[45] ));
 sky130_fd_sc_hd__dfxtp_1 _10343_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_00930_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[46] ));
 sky130_fd_sc_hd__dfxtp_1 _10344_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_00931_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[48] ));
 sky130_fd_sc_hd__dfxtp_1 _10345_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_00932_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[49] ));
 sky130_fd_sc_hd__dfxtp_1 _10346_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_00933_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[50] ));
 sky130_fd_sc_hd__dfxtp_1 _10347_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_00934_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[51] ));
 sky130_fd_sc_hd__dfxtp_1 _10348_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_00935_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[52] ));
 sky130_fd_sc_hd__dfxtp_1 _10349_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_00936_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[53] ));
 sky130_fd_sc_hd__dfxtp_1 _10350_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_00937_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[54] ));
 sky130_fd_sc_hd__dfxtp_1 _10351_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00938_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _10352_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00939_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _10353_ (.CLK(clknet_leaf_38_wbm_clk_i),
    .D(_00940_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _10354_ (.CLK(clknet_leaf_51_wbm_clk_i),
    .D(_00941_),
    .Q(net25));
 sky130_fd_sc_hd__dfstp_1 _10355_ (.CLK(clknet_leaf_42_wbm_clk_i),
    .D(_00942_),
    .SET_B(net268),
    .Q(\u_reg.cfg_glb_ctrl[0] ));
 sky130_fd_sc_hd__dfstp_2 _10356_ (.CLK(clknet_leaf_42_wbm_clk_i),
    .D(_00943_),
    .SET_B(net268),
    .Q(\u_reg.cfg_glb_ctrl[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10357_ (.CLK(clknet_leaf_42_wbm_clk_i),
    .D(_00944_),
    .RESET_B(net268),
    .Q(\u_reg.cfg_glb_ctrl[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10358_ (.CLK(clknet_leaf_42_wbm_clk_i),
    .D(_00945_),
    .RESET_B(net268),
    .Q(\u_reg.cfg_glb_ctrl[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10359_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00946_),
    .RESET_B(net268),
    .Q(\u_reg.cfg_glb_ctrl[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10360_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00947_),
    .RESET_B(net268),
    .Q(\u_reg.cfg_glb_ctrl[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10361_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00948_),
    .RESET_B(net268),
    .Q(\u_reg.cfg_glb_ctrl[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10362_ (.CLK(clknet_leaf_33_wbm_clk_i),
    .D(_00949_),
    .RESET_B(net269),
    .Q(\u_reg.cfg_glb_ctrl[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10363_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_00950_),
    .RESET_B(net247),
    .Q(\u_uart2wb.u_core.u_txfsm.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10364_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_00951_),
    .RESET_B(net247),
    .Q(\u_uart2wb.u_core.u_txfsm.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10365_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_00952_),
    .RESET_B(net248),
    .Q(\u_uart2wb.u_core.u_txfsm.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10366_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(_00953_),
    .RESET_B(net232),
    .Q(\u_uart2wb.reg_wr ));
 sky130_fd_sc_hd__dfrtp_1 _10367_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(_00954_),
    .RESET_B(net232),
    .Q(\u_uart2wb.reg_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10368_ (.CLK(\clknet_leaf_0_u_uart2wb.baud_clk_16x ),
    .D(_00955_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10369_ (.CLK(\clknet_leaf_0_u_uart2wb.baud_clk_16x ),
    .D(_00956_),
    .RESET_B(net231),
    .Q(\u_uart2wb.reg_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10370_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(_00957_),
    .RESET_B(net232),
    .Q(\u_uart2wb.reg_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10371_ (.CLK(\clknet_leaf_0_u_uart2wb.baud_clk_16x ),
    .D(_00958_),
    .RESET_B(net232),
    .Q(\u_uart2wb.reg_addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10372_ (.CLK(\clknet_leaf_0_u_uart2wb.baud_clk_16x ),
    .D(_00959_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10373_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00960_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_addr[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10374_ (.CLK(\clknet_leaf_0_u_uart2wb.baud_clk_16x ),
    .D(_00961_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_addr[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10375_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00962_),
    .RESET_B(net232),
    .Q(\u_uart2wb.reg_addr[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10376_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00963_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_addr[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10377_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00964_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_addr[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10378_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00965_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_addr[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10379_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00966_),
    .RESET_B(net232),
    .Q(\u_uart2wb.reg_addr[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10380_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00967_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_addr[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10381_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00968_),
    .RESET_B(net231),
    .Q(\u_uart2wb.reg_addr[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10382_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00969_),
    .RESET_B(net231),
    .Q(\u_uart2wb.reg_addr[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10383_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00970_),
    .RESET_B(net231),
    .Q(\u_uart2wb.reg_addr[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10384_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00971_),
    .RESET_B(net231),
    .Q(\u_uart2wb.reg_addr[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10385_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00972_),
    .RESET_B(net232),
    .Q(\u_uart2wb.reg_addr[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10386_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_00973_),
    .RESET_B(net232),
    .Q(\u_uart2wb.reg_addr[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10387_ (.CLK(\clknet_leaf_3_u_uart2wb.baud_clk_16x ),
    .D(_00974_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10388_ (.CLK(\clknet_leaf_0_u_uart2wb.baud_clk_16x ),
    .D(_00975_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_wdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10389_ (.CLK(\clknet_leaf_3_u_uart2wb.baud_clk_16x ),
    .D(_00976_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10390_ (.CLK(\clknet_leaf_0_u_uart2wb.baud_clk_16x ),
    .D(_00977_),
    .RESET_B(net230),
    .Q(\u_uart2wb.reg_wdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10391_ (.CLK(\clknet_leaf_3_u_uart2wb.baud_clk_16x ),
    .D(_00978_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10392_ (.CLK(\clknet_leaf_3_u_uart2wb.baud_clk_16x ),
    .D(_00979_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10393_ (.CLK(\clknet_leaf_3_u_uart2wb.baud_clk_16x ),
    .D(_00980_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10394_ (.CLK(\clknet_leaf_3_u_uart2wb.baud_clk_16x ),
    .D(_00981_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10395_ (.CLK(\clknet_leaf_5_u_uart2wb.baud_clk_16x ),
    .D(_00982_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10396_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00983_),
    .RESET_B(net234),
    .Q(\u_uart2wb.reg_wdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10397_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00984_),
    .RESET_B(net234),
    .Q(\u_uart2wb.reg_wdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10398_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00985_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10399_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00986_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10400_ (.CLK(\clknet_leaf_3_u_uart2wb.baud_clk_16x ),
    .D(_00987_),
    .RESET_B(net234),
    .Q(\u_uart2wb.reg_wdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10401_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00988_),
    .RESET_B(net234),
    .Q(\u_uart2wb.reg_wdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10402_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00989_),
    .RESET_B(net234),
    .Q(\u_uart2wb.reg_wdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10403_ (.CLK(\clknet_leaf_5_u_uart2wb.baud_clk_16x ),
    .D(_00990_),
    .RESET_B(net233),
    .Q(\u_uart2wb.reg_wdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10404_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00991_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10405_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00992_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10406_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00993_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10407_ (.CLK(\clknet_leaf_5_u_uart2wb.baud_clk_16x ),
    .D(_00994_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10408_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00995_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10409_ (.CLK(\clknet_leaf_5_u_uart2wb.baud_clk_16x ),
    .D(_00996_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10410_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00997_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10411_ (.CLK(\clknet_leaf_5_u_uart2wb.baud_clk_16x ),
    .D(_00998_),
    .RESET_B(net236),
    .Q(\u_uart2wb.reg_wdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10412_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_00999_),
    .RESET_B(net236),
    .Q(\u_uart2wb.reg_wdata[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10413_ (.CLK(\clknet_leaf_5_u_uart2wb.baud_clk_16x ),
    .D(_01000_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10414_ (.CLK(\clknet_leaf_4_u_uart2wb.baud_clk_16x ),
    .D(_01001_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10415_ (.CLK(\clknet_leaf_5_u_uart2wb.baud_clk_16x ),
    .D(_01002_),
    .RESET_B(net241),
    .Q(\u_uart2wb.reg_wdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10416_ (.CLK(\clknet_leaf_7_u_uart2wb.baud_clk_16x ),
    .D(_01003_),
    .RESET_B(net235),
    .Q(\u_uart2wb.reg_wdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10417_ (.CLK(\clknet_leaf_6_u_uart2wb.baud_clk_16x ),
    .D(_01004_),
    .RESET_B(net241),
    .Q(\u_uart2wb.reg_wdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10418_ (.CLK(\clknet_leaf_5_u_uart2wb.baud_clk_16x ),
    .D(_01005_),
    .RESET_B(net241),
    .Q(\u_uart2wb.reg_wdata[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10419_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_01006_),
    .RESET_B(net239),
    .Q(\u_uart2wb.reg_req ));
 sky130_fd_sc_hd__dfrtp_2 _10420_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_01007_),
    .RESET_B(net243),
    .Q(\u_uart2wb.tx_data_avail ));
 sky130_fd_sc_hd__dfrtp_1 _10421_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_01008_),
    .RESET_B(net248),
    .Q(\u_uart2wb.u_core.u_txfsm.txdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10422_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_01009_),
    .RESET_B(net247),
    .Q(\u_uart2wb.u_core.u_txfsm.txdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10423_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_01010_),
    .RESET_B(net250),
    .Q(\u_uart2wb.u_core.u_txfsm.txdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10424_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_01011_),
    .RESET_B(net250),
    .Q(\u_uart2wb.u_core.u_txfsm.txdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10425_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_01012_),
    .RESET_B(net247),
    .Q(\u_uart2wb.u_core.u_txfsm.txdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10426_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_01013_),
    .RESET_B(net250),
    .Q(\u_uart2wb.u_core.u_txfsm.txdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10427_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_01014_),
    .RESET_B(net250),
    .Q(\u_uart2wb.u_core.u_txfsm.txdata[6] ));
 sky130_fd_sc_hd__dfxtp_1 _10428_ (.CLK(\clknet_leaf_8_u_uart2wb.baud_clk_16x ),
    .D(_01015_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[64] ));
 sky130_fd_sc_hd__dfxtp_1 _10429_ (.CLK(\clknet_leaf_8_u_uart2wb.baud_clk_16x ),
    .D(_01016_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[65] ));
 sky130_fd_sc_hd__dfxtp_1 _10430_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_01017_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[66] ));
 sky130_fd_sc_hd__dfxtp_1 _10431_ (.CLK(\clknet_leaf_8_u_uart2wb.baud_clk_16x ),
    .D(_01018_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[67] ));
 sky130_fd_sc_hd__dfxtp_1 _10432_ (.CLK(\clknet_leaf_14_u_uart2wb.baud_clk_16x ),
    .D(_01019_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[68] ));
 sky130_fd_sc_hd__dfxtp_1 _10433_ (.CLK(\clknet_leaf_2_u_uart2wb.baud_clk_16x ),
    .D(_01020_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[69] ));
 sky130_fd_sc_hd__dfxtp_1 _10434_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_01021_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[70] ));
 sky130_fd_sc_hd__dfxtp_1 _10435_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_01022_),
    .Q(\u_uart2wb.u_msg.TxMsgSize[0] ));
 sky130_fd_sc_hd__dfxtp_1 _10436_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_01023_),
    .Q(\u_uart2wb.u_msg.TxMsgSize[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10437_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_01024_),
    .Q(\u_uart2wb.u_msg.TxMsgSize[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10438_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_01025_),
    .Q(\u_uart2wb.u_msg.TxMsgSize[3] ));
 sky130_fd_sc_hd__dfxtp_1 _10439_ (.CLK(\clknet_leaf_15_u_uart2wb.baud_clk_16x ),
    .D(_01026_),
    .Q(\u_uart2wb.u_msg.TxMsgSize[4] ));
 sky130_fd_sc_hd__dfxtp_1 _10440_ (.CLK(\clknet_leaf_24_u_uart2wb.baud_clk_16x ),
    .D(_01027_),
    .Q(\u_uart2wb.u_msg.RxMsgCnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _10441_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_01028_),
    .Q(\u_uart2wb.u_msg.RxMsgCnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10442_ (.CLK(\clknet_leaf_21_u_uart2wb.baud_clk_16x ),
    .D(_01029_),
    .Q(\u_uart2wb.u_msg.RxMsgCnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10443_ (.CLK(\clknet_leaf_21_u_uart2wb.baud_clk_16x ),
    .D(_01030_),
    .Q(\u_uart2wb.u_msg.RxMsgCnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _10444_ (.CLK(\clknet_leaf_21_u_uart2wb.baud_clk_16x ),
    .D(_01031_),
    .Q(\u_uart2wb.u_msg.RxMsgCnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10445_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_01032_),
    .RESET_B(net239),
    .Q(\u_uart2wb.u_msg.State[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10446_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_01033_),
    .RESET_B(net238),
    .Q(\u_uart2wb.u_msg.State[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10447_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_01034_),
    .RESET_B(net243),
    .Q(\u_uart2wb.u_msg.State[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10448_ (.CLK(\clknet_leaf_22_u_uart2wb.baud_clk_16x ),
    .D(_01035_),
    .RESET_B(net243),
    .Q(\u_uart2wb.u_msg.State[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10449_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_01036_),
    .RESET_B(net238),
    .Q(\u_uart2wb.u_msg.NextState[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10450_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_01037_),
    .RESET_B(net239),
    .Q(\u_uart2wb.u_msg.NextState[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10451_ (.CLK(\clknet_leaf_21_u_uart2wb.baud_clk_16x ),
    .D(_01038_),
    .RESET_B(net243),
    .Q(\u_uart2wb.u_msg.NextState[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10452_ (.CLK(\clknet_leaf_23_u_uart2wb.baud_clk_16x ),
    .D(_01039_),
    .RESET_B(net243),
    .Q(\u_uart2wb.u_msg.NextState[3] ));
 sky130_fd_sc_hd__dfxtp_1 _10453_ (.CLK(\clknet_leaf_24_u_uart2wb.baud_clk_16x ),
    .D(_01040_),
    .Q(\u_uart2wb.u_msg.cmd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _10454_ (.CLK(\clknet_leaf_26_u_uart2wb.baud_clk_16x ),
    .D(_01041_),
    .Q(\u_uart2wb.u_msg.cmd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10455_ (.CLK(\clknet_leaf_26_u_uart2wb.baud_clk_16x ),
    .D(_01042_),
    .Q(\u_uart2wb.u_msg.cmd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10456_ (.CLK(\clknet_leaf_26_u_uart2wb.baud_clk_16x ),
    .D(_01043_),
    .Q(\u_uart2wb.u_msg.cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _10457_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_01044_),
    .Q(\u_uart2wb.u_msg.cmd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _10458_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_01045_),
    .Q(\u_uart2wb.u_msg.cmd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _10459_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_01046_),
    .Q(\u_uart2wb.u_msg.cmd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _10460_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_01047_),
    .Q(\u_uart2wb.u_msg.cmd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _10461_ (.CLK(\clknet_leaf_1_u_uart2wb.baud_clk_16x ),
    .D(_01048_),
    .Q(\u_uart2wb.u_msg.cmd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _10462_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_01049_),
    .Q(\u_uart2wb.u_msg.cmd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _10463_ (.CLK(\clknet_leaf_27_u_uart2wb.baud_clk_16x ),
    .D(_01050_),
    .Q(\u_uart2wb.u_msg.cmd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _10464_ (.CLK(\clknet_leaf_26_u_uart2wb.baud_clk_16x ),
    .D(_01051_),
    .Q(\u_uart2wb.u_msg.cmd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _10465_ (.CLK(\clknet_leaf_26_u_uart2wb.baud_clk_16x ),
    .D(_01052_),
    .Q(\u_uart2wb.u_msg.cmd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _10466_ (.CLK(\clknet_leaf_25_u_uart2wb.baud_clk_16x ),
    .D(_01053_),
    .Q(\u_uart2wb.u_msg.cmd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _10467_ (.CLK(\clknet_leaf_26_u_uart2wb.baud_clk_16x ),
    .D(_01054_),
    .Q(\u_uart2wb.u_msg.cmd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _10468_ (.CLK(\clknet_leaf_26_u_uart2wb.baud_clk_16x ),
    .D(_01055_),
    .Q(\u_uart2wb.u_msg.cmd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _10469_ (.CLK(\clknet_leaf_16_u_uart2wb.baud_clk_16x ),
    .D(_01056_),
    .Q(\u_uart2wb.tx_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _10470_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_01057_),
    .Q(\u_uart2wb.tx_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10471_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_01058_),
    .Q(\u_uart2wb.tx_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10472_ (.CLK(\clknet_leaf_17_u_uart2wb.baud_clk_16x ),
    .D(_01059_),
    .Q(\u_uart2wb.tx_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _10473_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_01060_),
    .Q(\u_uart2wb.tx_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _10474_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_01061_),
    .Q(\u_uart2wb.tx_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _10475_ (.CLK(\clknet_leaf_13_u_uart2wb.baud_clk_16x ),
    .D(_01062_),
    .Q(\u_uart2wb.tx_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _10476_ (.CLK(\clknet_leaf_9_u_uart2wb.baud_clk_16x ),
    .D(_01063_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[88] ));
 sky130_fd_sc_hd__dfxtp_1 _10477_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_01064_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[89] ));
 sky130_fd_sc_hd__dfxtp_1 _10478_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_01065_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[90] ));
 sky130_fd_sc_hd__dfxtp_1 _10479_ (.CLK(\clknet_leaf_10_u_uart2wb.baud_clk_16x ),
    .D(_01066_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[91] ));
 sky130_fd_sc_hd__dfxtp_1 _10480_ (.CLK(\clknet_leaf_8_u_uart2wb.baud_clk_16x ),
    .D(_01067_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[92] ));
 sky130_fd_sc_hd__dfxtp_1 _10481_ (.CLK(\clknet_leaf_9_u_uart2wb.baud_clk_16x ),
    .D(_01068_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[93] ));
 sky130_fd_sc_hd__dfxtp_1 _10482_ (.CLK(\clknet_leaf_8_u_uart2wb.baud_clk_16x ),
    .D(_01069_),
    .Q(\u_uart2wb.u_msg.TxMsgBuf[94] ));
 sky130_fd_sc_hd__dfrtp_4 _10483_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_01070_),
    .RESET_B(net262),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _10484_ (.CLK(clknet_leaf_88_wbm_clk_i),
    .D(_01071_),
    .RESET_B(net262),
    .Q(\u_spi2wb.u_if.RegSdOut[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10485_ (.CLK(clknet_leaf_89_wbm_clk_i),
    .D(_01072_),
    .RESET_B(net262),
    .Q(\u_spi2wb.u_if.RegSdOut[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10486_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_01073_),
    .RESET_B(net262),
    .Q(\u_spi2wb.u_if.RegSdOut[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10487_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_01074_),
    .RESET_B(net262),
    .Q(\u_spi2wb.u_if.RegSdOut[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10488_ (.CLK(clknet_leaf_13_wbm_clk_i),
    .D(_01075_),
    .RESET_B(net263),
    .Q(\u_spi2wb.u_if.RegSdOut[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10489_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_01076_),
    .RESET_B(net263),
    .Q(\u_spi2wb.u_if.RegSdOut[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10490_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_01077_),
    .RESET_B(net263),
    .Q(\u_spi2wb.u_if.RegSdOut[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10491_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_01078_),
    .RESET_B(net261),
    .Q(\u_spi2wb.u_if.RegSdOut[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10492_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_01079_),
    .RESET_B(net261),
    .Q(\u_spi2wb.u_if.RegSdOut[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10493_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_01080_),
    .RESET_B(net261),
    .Q(\u_spi2wb.u_if.RegSdOut[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10494_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_01081_),
    .RESET_B(net261),
    .Q(\u_spi2wb.u_if.RegSdOut[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10495_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_01082_),
    .RESET_B(net261),
    .Q(\u_spi2wb.u_if.RegSdOut[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10496_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_01083_),
    .RESET_B(net261),
    .Q(\u_spi2wb.u_if.RegSdOut[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10497_ (.CLK(clknet_leaf_7_wbm_clk_i),
    .D(_01084_),
    .RESET_B(net258),
    .Q(\u_spi2wb.u_if.RegSdOut[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10498_ (.CLK(clknet_leaf_8_wbm_clk_i),
    .D(_01085_),
    .RESET_B(net258),
    .Q(\u_spi2wb.u_if.RegSdOut[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10499_ (.CLK(clknet_leaf_8_wbm_clk_i),
    .D(_01086_),
    .RESET_B(net259),
    .Q(\u_spi2wb.u_if.RegSdOut[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10500_ (.CLK(clknet_leaf_8_wbm_clk_i),
    .D(_01087_),
    .RESET_B(net259),
    .Q(\u_spi2wb.u_if.RegSdOut[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10501_ (.CLK(clknet_leaf_8_wbm_clk_i),
    .D(_01088_),
    .RESET_B(net259),
    .Q(\u_spi2wb.u_if.RegSdOut[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10502_ (.CLK(clknet_leaf_8_wbm_clk_i),
    .D(_01089_),
    .RESET_B(net262),
    .Q(\u_spi2wb.u_if.RegSdOut[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10503_ (.CLK(clknet_leaf_11_wbm_clk_i),
    .D(_01090_),
    .RESET_B(net262),
    .Q(\u_spi2wb.u_if.RegSdOut[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10504_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_01091_),
    .RESET_B(net262),
    .Q(\u_spi2wb.u_if.RegSdOut[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10505_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_01092_),
    .RESET_B(net260),
    .Q(\u_spi2wb.u_if.RegSdOut[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10506_ (.CLK(clknet_leaf_9_wbm_clk_i),
    .D(_01093_),
    .RESET_B(net260),
    .Q(\u_spi2wb.u_if.RegSdOut[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10507_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_01094_),
    .RESET_B(net260),
    .Q(\u_spi2wb.u_if.RegSdOut[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10508_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_01095_),
    .RESET_B(net260),
    .Q(\u_spi2wb.u_if.RegSdOut[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10509_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_01096_),
    .RESET_B(net260),
    .Q(\u_spi2wb.u_if.RegSdOut[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10510_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_01097_),
    .RESET_B(net261),
    .Q(\u_spi2wb.u_if.RegSdOut[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10511_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_01098_),
    .RESET_B(net261),
    .Q(\u_spi2wb.u_if.RegSdOut[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10512_ (.CLK(clknet_leaf_89_wbm_clk_i),
    .D(_01099_),
    .RESET_B(net263),
    .Q(\u_spi2wb.u_if.RegSdOut[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10513_ (.CLK(clknet_leaf_10_wbm_clk_i),
    .D(_01100_),
    .RESET_B(net261),
    .Q(\u_spi2wb.u_if.RegSdOut[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10514_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_01101_),
    .RESET_B(net262),
    .Q(\u_spi2wb.u_if.RegSdOut[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10515_ (.CLK(clknet_leaf_12_wbm_clk_i),
    .D(_01102_),
    .RESET_B(net263),
    .Q(\u_spi2wb.u_if.RegSdOut[31] ));
 sky130_fd_sc_hd__dfstp_2 _10516_ (.CLK(clknet_leaf_72_wbm_clk_i),
    .D(_01103_),
    .SET_B(net271),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_4 _10517_ (.CLK(clknet_leaf_74_wbm_clk_i),
    .D(_01104_),
    .RESET_B(net271),
    .Q(\u_spi2wb.reg_wr ));
 sky130_fd_sc_hd__buf_6 _10529_ (.A(net176),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_async_wb.u_cmd_if.rd_clk  (.A(\u_async_wb.u_cmd_if.rd_clk ),
    .X(\clknet_0_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_uart2wb.baud_clk_16x  (.A(\u_uart2wb.baud_clk_16x ),
    .X(\clknet_0_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wbm_clk_i (.A(net320),
    .X(clknet_0_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_uart2wb.baud_clk_16x  (.A(\clknet_0_u_uart2wb.baud_clk_16x ),
    .X(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_uart2wb.baud_clk_16x  (.A(\clknet_0_u_uart2wb.baud_clk_16x ),
    .X(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_0__f_u_async_wb.u_cmd_if.rd_clk  (.A(\clknet_0_u_async_wb.u_cmd_if.rd_clk ),
    .X(\clknet_3_0__leaf_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wbm_clk_i (.A(clknet_0_wbm_clk_i),
    .X(clknet_3_0__leaf_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_1__f_u_async_wb.u_cmd_if.rd_clk  (.A(\clknet_0_u_async_wb.u_cmd_if.rd_clk ),
    .X(\clknet_3_1__leaf_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wbm_clk_i (.A(clknet_0_wbm_clk_i),
    .X(clknet_3_1__leaf_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_2__f_u_async_wb.u_cmd_if.rd_clk  (.A(\clknet_0_u_async_wb.u_cmd_if.rd_clk ),
    .X(\clknet_3_2__leaf_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wbm_clk_i (.A(clknet_0_wbm_clk_i),
    .X(clknet_3_2__leaf_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_3__f_u_async_wb.u_cmd_if.rd_clk  (.A(\clknet_0_u_async_wb.u_cmd_if.rd_clk ),
    .X(\clknet_3_3__leaf_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wbm_clk_i (.A(clknet_0_wbm_clk_i),
    .X(clknet_3_3__leaf_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_4__f_u_async_wb.u_cmd_if.rd_clk  (.A(\clknet_0_u_async_wb.u_cmd_if.rd_clk ),
    .X(\clknet_3_4__leaf_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wbm_clk_i (.A(clknet_0_wbm_clk_i),
    .X(clknet_3_4__leaf_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_5__f_u_async_wb.u_cmd_if.rd_clk  (.A(\clknet_0_u_async_wb.u_cmd_if.rd_clk ),
    .X(\clknet_3_5__leaf_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wbm_clk_i (.A(clknet_0_wbm_clk_i),
    .X(clknet_3_5__leaf_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_6__f_u_async_wb.u_cmd_if.rd_clk  (.A(\clknet_0_u_async_wb.u_cmd_if.rd_clk ),
    .X(\clknet_3_6__leaf_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wbm_clk_i (.A(clknet_0_wbm_clk_i),
    .X(clknet_3_6__leaf_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_7__f_u_async_wb.u_cmd_if.rd_clk  (.A(\clknet_0_u_async_wb.u_cmd_if.rd_clk ),
    .X(\clknet_3_7__leaf_u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wbm_clk_i (.A(clknet_0_wbm_clk_i),
    .X(clknet_3_7__leaf_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_0_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_0_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_0_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_10_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_10_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_10_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_11_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_11_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_11_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_12_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_12_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_12_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_13_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_13_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_13_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_14_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_14_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_14_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_15_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_15_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_15_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_16_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_16_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_16_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_17_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_17_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_17_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_18_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_18_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_18_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_19_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_19_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_19_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_1_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_1_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_1_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_20_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_20_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_20_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_21_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_21_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_21_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_22_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_22_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_22_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_23_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_23_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_23_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_24_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_24_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_24_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_25_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_25_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_25_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_26_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_26_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_26_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_27_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_27_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_27_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_28_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_29_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_2_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_2_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_2_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_30_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_31_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_32_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wbm_clk_i (.A(clknet_3_2__leaf_wbm_clk_i),
    .X(clknet_leaf_33_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_34_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_35_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_36_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_37_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_38_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_39_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_3_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_3_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_3_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_40_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_41_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_42_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_43_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_44_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wbm_clk_i (.A(clknet_3_3__leaf_wbm_clk_i),
    .X(clknet_leaf_45_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_46_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_47_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_48_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_49_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_4_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_4_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_4_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_50_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_51_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_52_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_53_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_54_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_wbm_clk_i (.A(clknet_3_6__leaf_wbm_clk_i),
    .X(clknet_leaf_55_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_wbm_clk_i (.A(clknet_3_7__leaf_wbm_clk_i),
    .X(clknet_leaf_56_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_wbm_clk_i (.A(clknet_3_7__leaf_wbm_clk_i),
    .X(clknet_leaf_57_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_wbm_clk_i (.A(clknet_3_7__leaf_wbm_clk_i),
    .X(clknet_leaf_58_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_wbm_clk_i (.A(clknet_3_7__leaf_wbm_clk_i),
    .X(clknet_leaf_59_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_5_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_5_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_5_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_wbm_clk_i (.A(clknet_3_7__leaf_wbm_clk_i),
    .X(clknet_leaf_60_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_wbm_clk_i (.A(clknet_3_7__leaf_wbm_clk_i),
    .X(clknet_leaf_61_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_wbm_clk_i (.A(clknet_3_7__leaf_wbm_clk_i),
    .X(clknet_leaf_62_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_wbm_clk_i (.A(clknet_3_7__leaf_wbm_clk_i),
    .X(clknet_leaf_63_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_64_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_65_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_66_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_67_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_68_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_69_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_6_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_6_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_6_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_70_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_71_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_72_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_73_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_74_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_75_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_76_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_wbm_clk_i (.A(clknet_3_4__leaf_wbm_clk_i),
    .X(clknet_leaf_77_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_78_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_79_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_7_u_uart2wb.baud_clk_16x  (.A(\clknet_1_0__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_7_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_7_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_80_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_81_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_82_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_83_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_84_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_85_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_86_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_wbm_clk_i (.A(clknet_3_5__leaf_wbm_clk_i),
    .X(clknet_leaf_87_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_88_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_89_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_8_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_8_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_8_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_90_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_91_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_92_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_93_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_wbm_clk_i (.A(clknet_3_0__leaf_wbm_clk_i),
    .X(clknet_leaf_94_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_leaf_9_u_uart2wb.baud_clk_16x  (.A(\clknet_1_1__leaf_u_uart2wb.baud_clk_16x ),
    .X(\clknet_leaf_9_u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wbm_clk_i (.A(clknet_3_1__leaf_wbm_clk_i),
    .X(clknet_leaf_9_wbm_clk_i));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__buf_2 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(net251),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net236),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 fanout234 (.A(net236),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 fanout236 (.A(net251),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 fanout237 (.A(net242),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout238 (.A(net242),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 fanout239 (.A(net242),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_4 fanout240 (.A(net242),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_4 fanout242 (.A(net251),
    .X(net242));
 sky130_fd_sc_hd__buf_4 fanout243 (.A(net245),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(net251),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(net250),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_4 fanout251 (.A(\u_uart2wb.line_reset_n ),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_4 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_4 fanout253 (.A(\u_async_wb.u_cmd_if.rd_reset_n ),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__buf_4 fanout256 (.A(net259),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 fanout259 (.A(net269),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_4 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__buf_4 fanout261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__buf_4 fanout262 (.A(net264),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__buf_2 fanout264 (.A(net269),
    .X(net264));
 sky130_fd_sc_hd__buf_4 fanout265 (.A(net267),
    .X(net265));
 sky130_fd_sc_hd__buf_2 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_4 fanout267 (.A(net269),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_4 fanout268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__buf_4 fanout269 (.A(net68),
    .X(net269));
 sky130_fd_sc_hd__buf_4 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net275),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(net275),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(net68),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 fanout278 (.A(net284),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(net284),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(net283),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_4 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_2 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(\u_uart2wb.arst_ssn ),
    .X(net285));
 sky130_fd_sc_hd__buf_4 fanout286 (.A(net291),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_2 fanout288 (.A(net291),
    .X(net288));
 sky130_fd_sc_hd__buf_4 fanout289 (.A(net291),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 fanout291 (.A(net342),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_4 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_4 fanout295 (.A(net301),
    .X(net295));
 sky130_fd_sc_hd__buf_4 fanout296 (.A(net298),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_2 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__buf_2 fanout299 (.A(net301),
    .X(net299));
 sky130_fd_sc_hd__buf_4 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_2 fanout301 (.A(net70),
    .X(net301));
 sky130_fd_sc_hd__buf_4 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__buf_4 fanout304 (.A(net341),
    .X(net304));
 sky130_fd_sc_hd__buf_4 fanout305 (.A(net341),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\u_async_wb.wbs_ack_f ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_01727_),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\u_async_wb.u_cmd_if.sync_wr_ptr[2] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_01467_),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_01468_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(wbm_rst_i),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\u_async_wb.u_cmd_if.rd_ptr[1] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_01469_),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\u_wbs_rst.in_data_2s ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\u_uart2wb.u_arst_sync.in_data_2s ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\u_async_wb.u_cmd_if.rd_ptr[0] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net70),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net69),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\u_async_wb.u_cmd_if.sync_rd_ptr_0[0] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\u_spi2wb.u_if.sck_l0 ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\u_uart2wb.u_core.u_rxd_sync.in_data_2s ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\u_async_wb.u_resp_if.sync_wr_ptr_0[0] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\u_wbs_rst.in_data_s ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\u_reset_fsm.boot_req_s ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\u_wbm_rst.in_data_2s ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\u_async_wb.u_resp_if.sync_rd_ptr_0[1] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\u_async_wb.u_resp_if.sync_rd_ptr_0[0] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\u_wbm_rst.in_data_s ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\u_async_wb.u_cmd_if.sync_wr_ptr_0[2] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\u_uart2wb.u_arst_sync.in_data_s ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\u_uart2wb.u_aut_det.rxd_sync[0] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\u_async_wb.u_cmd_if.sync_rd_ptr_0[1] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\u_async_wb.u_cmd_if.sync_rd_ptr_0[2] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\u_async_wb.u_resp_if.sync_wr_ptr_0[1] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\u_uart2wb.u_core.u_line_rst.in_data_s ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\u_uart2wb.u_async_reg_bus.out_flag_s ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\u_async_wb.u_cmd_if.sync_wr_ptr_0[1] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\u_async_wb.u_cmd_if.sync_wr_ptr_0[0] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\u_spi2wb.u_if.ssn_l0 ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\u_spi2wb.u_if.sck_l1 ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\u_uart2wb.u_async_reg_bus.in_flag_s ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\u_uart2wb.u_core.u_rxd_sync.in_data_s ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(wbm_stb_i),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\u_spi2wb.u_if.ssn_l1 ),
    .X(net368));
 sky130_fd_sc_hd__buf_2 output1 (.A(net1),
    .X(cfg_clk_skew_ctrl1[0]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(cfg_clk_skew_ctrl1[18]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(system_strap[5]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(system_strap[6]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(system_strap[7]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(system_strap[8]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(system_strap[9]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(uartm_txd));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(wbd_clk_wh));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(wbd_int_rst_n));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(wbd_pll_rst_n));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(wbm_ack_o));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(cfg_clk_skew_ctrl1[19]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(wbm_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(wbm_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(wbm_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(wbm_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(wbm_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(wbm_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(wbm_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(wbm_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(wbm_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(wbm_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(cfg_clk_skew_ctrl1[1]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(wbm_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(wbm_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(wbm_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(wbm_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(wbm_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(wbm_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(wbm_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(wbm_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(wbm_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(wbm_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(cfg_clk_skew_ctrl1[20]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(wbm_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(wbm_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(wbm_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(wbm_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(wbm_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(wbm_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(wbm_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(wbm_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(wbm_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(wbm_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(cfg_clk_skew_ctrl1[21]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(wbm_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(wbm_dat_o[9]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(wbm_err_o));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(wbs_adr_o[0]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(wbs_adr_o[10]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(wbs_adr_o[11]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(wbs_adr_o[12]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(wbs_adr_o[13]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(wbs_adr_o[14]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(wbs_adr_o[15]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(cfg_clk_skew_ctrl1[22]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(wbs_adr_o[16]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(wbs_adr_o[17]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(wbs_adr_o[18]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(wbs_adr_o[19]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(wbs_adr_o[1]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(wbs_adr_o[20]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(wbs_adr_o[21]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(wbs_adr_o[22]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(wbs_adr_o[23]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(wbs_adr_o[24]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(cfg_clk_skew_ctrl1[23]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(wbs_adr_o[25]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(wbs_adr_o[26]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(wbs_adr_o[27]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(wbs_adr_o[28]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(wbs_adr_o[29]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(wbs_adr_o[2]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(wbs_adr_o[30]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(wbs_adr_o[31]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(wbs_adr_o[3]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(wbs_adr_o[4]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(cfg_clk_skew_ctrl1[24]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(wbs_adr_o[5]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(wbs_adr_o[6]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(wbs_adr_o[7]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(wbs_adr_o[8]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(wbs_adr_o[9]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(wbs_clk_out));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(wbs_cyc_o));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(cfg_clk_skew_ctrl1[25]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(cfg_clk_skew_ctrl1[26]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(cfg_clk_skew_ctrl1[10]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(cfg_clk_skew_ctrl1[27]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(wbs_sel_o[0]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(cfg_clk_skew_ctrl1[28]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(wbs_sel_o[1]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(wbs_sel_o[2]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(wbs_sel_o[3]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(wbs_stb_o));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(wbs_we_o));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(cfg_clk_skew_ctrl1[29]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(cfg_clk_skew_ctrl1[2]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(cfg_clk_skew_ctrl1[30]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(cfg_clk_skew_ctrl1[31]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(cfg_clk_skew_ctrl1[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(cfg_clk_skew_ctrl1[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(cfg_clk_skew_ctrl1[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(cfg_clk_skew_ctrl1[6]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(cfg_clk_skew_ctrl1[11]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(cfg_clk_skew_ctrl1[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(cfg_clk_skew_ctrl1[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(cfg_clk_skew_ctrl1[9]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(cfg_clk_skew_ctrl2[0]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(cfg_clk_skew_ctrl2[10]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(cfg_clk_skew_ctrl2[11]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(cfg_clk_skew_ctrl2[12]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(cfg_clk_skew_ctrl2[13]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(cfg_clk_skew_ctrl2[14]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(cfg_clk_skew_ctrl2[15]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(cfg_clk_skew_ctrl1[12]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(cfg_clk_skew_ctrl2[16]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(cfg_clk_skew_ctrl2[17]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(cfg_clk_skew_ctrl2[18]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(cfg_clk_skew_ctrl2[19]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(cfg_clk_skew_ctrl2[1]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(cfg_clk_skew_ctrl2[20]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(cfg_clk_skew_ctrl2[21]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(cfg_clk_skew_ctrl2[22]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(cfg_clk_skew_ctrl2[23]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(cfg_clk_skew_ctrl2[24]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(cfg_clk_skew_ctrl1[13]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(cfg_clk_skew_ctrl2[25]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(cfg_clk_skew_ctrl2[26]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(cfg_clk_skew_ctrl2[27]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(cfg_clk_skew_ctrl2[28]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(cfg_clk_skew_ctrl2[29]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(cfg_clk_skew_ctrl2[2]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(cfg_clk_skew_ctrl2[30]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(cfg_clk_skew_ctrl2[31]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(cfg_clk_skew_ctrl2[3]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(cfg_clk_skew_ctrl2[4]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(cfg_clk_skew_ctrl1[14]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(cfg_clk_skew_ctrl2[5]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(cfg_clk_skew_ctrl2[6]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(cfg_clk_skew_ctrl2[7]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(cfg_clk_skew_ctrl2[8]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(cfg_clk_skew_ctrl2[9]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(cfg_fast_sim));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(cfg_strap_pad_ctrl));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(cpu_clk));
 sky130_fd_sc_hd__buf_2 output68 (.A(net274),
    .X(e_reset_n));
 sky130_fd_sc_hd__buf_2 output69 (.A(net290),
    .X(p_reset_n));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(cfg_clk_skew_ctrl1[15]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net304),
    .X(s_reset_n));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(sdout));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(sdout_oen));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(system_strap[0]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(system_strap[10]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(system_strap[11]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(system_strap[12]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(system_strap[13]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(system_strap[14]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(system_strap[15]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(cfg_clk_skew_ctrl1[16]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(system_strap[16]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(system_strap[17]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(system_strap[18]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(system_strap[19]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(system_strap[1]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(system_strap[20]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(system_strap[21]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(system_strap[22]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(system_strap[23]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(system_strap[24]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(cfg_clk_skew_ctrl1[17]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(system_strap[25]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(system_strap[26]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(system_strap[27]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(system_strap[28]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(system_strap[29]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(system_strap[2]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(system_strap[30]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(system_strap[31]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(system_strap[3]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(system_strap[4]));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(\u_skew_wh.clk_d9 ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(\u_skew_wh.clk_d11 ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(\u_skew_wh.clk_d10 ),
    .X(net323));
 sky130_fd_sc_hd__dlclkp_2 \u_clkgate.u_gate  (.CLK(wbs_clk_i),
    .GATE(net319),
    .GCLK(\u_async_wb.u_cmd_if.rd_clk ));
 sky130_fd_sc_hd__conb_1 \u_clkgate.u_gate_319  (.HI(net319));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \u_delay1_stb0.u_dly  (.A(\u_delay1_stb0.A ),
    .X(\u_delay1_stb0.X ));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \u_delay2_stb1.u_dly  (.A(\u_delay1_stb0.X ),
    .X(\u_delay2_stb1.X ));
 sky130_fd_sc_hd__clkdlybuf4s25_1 \u_delay2_stb2.u_dly  (.A(\u_delay2_stb1.X ),
    .X(\u_delay2_stb2.X ));
 sky130_fd_sc_hd__buf_2 \u_reg.u_buf_pll_rst.u_buf  (.A(\u_reg.u_buf_pll_rst.A ),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 \u_reg.u_buf_wb_rst.u_buf  (.A(\u_reg.u_buf_wb_rst.A ),
    .X(net107));
 sky130_fd_sc_hd__dlclkp_2 \u_reg.u_clkgate_cpu.u_gate  (.CLK(\u_reg.cpu_clk_div ),
    .GATE(\u_reg.clk_enb ),
    .GCLK(net67));
 sky130_fd_sc_hd__dlclkp_1 \u_reg.u_clkgate_wbs.u_gate  (.CLK(\u_reg.u_clkgate_wbs.CLK ),
    .GATE(\u_reg.clk_enb ),
    .GCLK(net175));
 sky130_fd_sc_hd__clkbuf_1 \u_reg.u_cpu_ref_clkbuf.u_buf  (.A(\u_reg.cpu_ref_clk_int ),
    .X(\u_reg.cpu_ref_clk ));
 sky130_fd_sc_hd__buf_4 \u_reg.u_fastsim_buf.u_buf  (.A(\u_reg.cfg_glb_ctrl[8] ),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 \u_reg.u_wbs_ref_clkbuf.u_buf  (.A(\u_reg.u_wbs_ref_clkbuf.A ),
    .X(\u_reg.u_wbclk.mclk ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_1.u_dly0  (.A(\u_skew_wh.clk_inbuf ),
    .X(\u_skew_wh.clkbuf_1.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_1.u_dly1  (.A(\u_skew_wh.clkbuf_1.X1 ),
    .X(\u_skew_wh.clkbuf_1.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_1.u_dly2  (.A(\u_skew_wh.clkbuf_1.X2 ),
    .X(\u_skew_wh.clkbuf_1.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_1.u_dly3  (.A(\u_skew_wh.clkbuf_1.X3 ),
    .X(\u_skew_wh.clk_d1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_10.u_dly0  (.A(\u_skew_wh.clk_d9 ),
    .X(\u_skew_wh.clkbuf_10.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_10.u_dly1  (.A(\u_skew_wh.clkbuf_10.X1 ),
    .X(\u_skew_wh.clkbuf_10.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_10.u_dly2  (.A(\u_skew_wh.clkbuf_10.X2 ),
    .X(\u_skew_wh.clkbuf_10.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_10.u_dly3  (.A(\u_skew_wh.clkbuf_10.X3 ),
    .X(\u_skew_wh.clk_d10 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_11.u_dly0  (.A(\u_skew_wh.clk_d10 ),
    .X(\u_skew_wh.clkbuf_11.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_11.u_dly1  (.A(\u_skew_wh.clkbuf_11.X1 ),
    .X(\u_skew_wh.clkbuf_11.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_11.u_dly2  (.A(\u_skew_wh.clkbuf_11.X2 ),
    .X(\u_skew_wh.clkbuf_11.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_11.u_dly3  (.A(\u_skew_wh.clkbuf_11.X3 ),
    .X(\u_skew_wh.clk_d11 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_12.u_dly0  (.A(\u_skew_wh.clk_d11 ),
    .X(\u_skew_wh.clkbuf_12.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_12.u_dly1  (.A(\u_skew_wh.clkbuf_12.X1 ),
    .X(\u_skew_wh.clkbuf_12.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_12.u_dly2  (.A(\u_skew_wh.clkbuf_12.X2 ),
    .X(\u_skew_wh.clkbuf_12.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_12.u_dly3  (.A(\u_skew_wh.clkbuf_12.X3 ),
    .X(\u_skew_wh.clk_d12 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_13.u_dly0  (.A(\u_skew_wh.clk_d12 ),
    .X(\u_skew_wh.clkbuf_13.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_13.u_dly1  (.A(\u_skew_wh.clkbuf_13.X1 ),
    .X(\u_skew_wh.clkbuf_13.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_13.u_dly2  (.A(\u_skew_wh.clkbuf_13.X2 ),
    .X(\u_skew_wh.clkbuf_13.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_13.u_dly3  (.A(\u_skew_wh.clkbuf_13.X3 ),
    .X(\u_skew_wh.clk_d13 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_14.u_dly0  (.A(\u_skew_wh.clk_d13 ),
    .X(\u_skew_wh.clkbuf_14.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_14.u_dly1  (.A(\u_skew_wh.clkbuf_14.X1 ),
    .X(\u_skew_wh.clkbuf_14.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_14.u_dly2  (.A(\u_skew_wh.clkbuf_14.X2 ),
    .X(\u_skew_wh.clkbuf_14.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_14.u_dly3  (.A(\u_skew_wh.clkbuf_14.X3 ),
    .X(\u_skew_wh.clk_d14 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_15.u_dly0  (.A(\u_skew_wh.clk_d14 ),
    .X(\u_skew_wh.clkbuf_15.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_15.u_dly1  (.A(\u_skew_wh.clkbuf_15.X1 ),
    .X(\u_skew_wh.clkbuf_15.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_15.u_dly2  (.A(\u_skew_wh.clkbuf_15.X2 ),
    .X(\u_skew_wh.clkbuf_15.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_15.u_dly3  (.A(\u_skew_wh.clkbuf_15.X3 ),
    .X(\u_skew_wh.clk_d15 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_2.u_dly0  (.A(\u_skew_wh.clk_d1 ),
    .X(\u_skew_wh.clkbuf_2.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_2.u_dly1  (.A(\u_skew_wh.clkbuf_2.X1 ),
    .X(\u_skew_wh.clkbuf_2.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_2.u_dly2  (.A(\u_skew_wh.clkbuf_2.X2 ),
    .X(\u_skew_wh.clkbuf_2.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_2.u_dly3  (.A(\u_skew_wh.clkbuf_2.X3 ),
    .X(\u_skew_wh.clk_d2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_3.u_dly0  (.A(\u_skew_wh.clk_d2 ),
    .X(\u_skew_wh.clkbuf_3.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_3.u_dly1  (.A(\u_skew_wh.clkbuf_3.X1 ),
    .X(\u_skew_wh.clkbuf_3.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_3.u_dly2  (.A(\u_skew_wh.clkbuf_3.X2 ),
    .X(\u_skew_wh.clkbuf_3.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_3.u_dly3  (.A(\u_skew_wh.clkbuf_3.X3 ),
    .X(\u_skew_wh.clk_d3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_4.u_dly0  (.A(\u_skew_wh.clk_d3 ),
    .X(\u_skew_wh.clkbuf_4.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_4.u_dly1  (.A(\u_skew_wh.clkbuf_4.X1 ),
    .X(\u_skew_wh.clkbuf_4.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_4.u_dly2  (.A(\u_skew_wh.clkbuf_4.X2 ),
    .X(\u_skew_wh.clkbuf_4.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_4.u_dly3  (.A(\u_skew_wh.clkbuf_4.X3 ),
    .X(\u_skew_wh.clk_d4 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_5.u_dly0  (.A(\u_skew_wh.clk_d4 ),
    .X(\u_skew_wh.clkbuf_5.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_5.u_dly1  (.A(\u_skew_wh.clkbuf_5.X1 ),
    .X(\u_skew_wh.clkbuf_5.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_5.u_dly2  (.A(\u_skew_wh.clkbuf_5.X2 ),
    .X(\u_skew_wh.clkbuf_5.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_5.u_dly3  (.A(\u_skew_wh.clkbuf_5.X3 ),
    .X(\u_skew_wh.clk_d5 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_6.u_dly0  (.A(\u_skew_wh.clk_d5 ),
    .X(\u_skew_wh.clkbuf_6.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_6.u_dly1  (.A(\u_skew_wh.clkbuf_6.X1 ),
    .X(\u_skew_wh.clkbuf_6.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_6.u_dly2  (.A(\u_skew_wh.clkbuf_6.X2 ),
    .X(\u_skew_wh.clkbuf_6.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_6.u_dly3  (.A(\u_skew_wh.clkbuf_6.X3 ),
    .X(\u_skew_wh.clk_d6 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_7.u_dly0  (.A(\u_skew_wh.clk_d6 ),
    .X(\u_skew_wh.clkbuf_7.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_7.u_dly1  (.A(\u_skew_wh.clkbuf_7.X1 ),
    .X(\u_skew_wh.clkbuf_7.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_7.u_dly2  (.A(\u_skew_wh.clkbuf_7.X2 ),
    .X(\u_skew_wh.clkbuf_7.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_7.u_dly3  (.A(\u_skew_wh.clkbuf_7.X3 ),
    .X(\u_skew_wh.clk_d7 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_8.u_dly0  (.A(\u_skew_wh.clk_d7 ),
    .X(\u_skew_wh.clkbuf_8.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_8.u_dly1  (.A(\u_skew_wh.clkbuf_8.X1 ),
    .X(\u_skew_wh.clkbuf_8.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_8.u_dly2  (.A(\u_skew_wh.clkbuf_8.X2 ),
    .X(\u_skew_wh.clkbuf_8.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_8.u_dly3  (.A(\u_skew_wh.clkbuf_8.X3 ),
    .X(\u_skew_wh.clk_d8 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_9.u_dly0  (.A(\u_skew_wh.clk_d8 ),
    .X(\u_skew_wh.clkbuf_9.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_9.u_dly1  (.A(\u_skew_wh.clkbuf_9.X1 ),
    .X(\u_skew_wh.clkbuf_9.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_9.u_dly2  (.A(\u_skew_wh.clkbuf_9.X2 ),
    .X(\u_skew_wh.clkbuf_9.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.clkbuf_9.u_dly3  (.A(\u_skew_wh.clkbuf_9.X3 ),
    .X(\u_skew_wh.clk_d9 ));
 sky130_fd_sc_hd__buf_6 \u_skew_wh.u_clkbuf_in.u_buf  (.A(wbd_clk_int),
    .X(\u_skew_wh.clk_inbuf ));
 sky130_fd_sc_hd__clkbuf_2 \u_skew_wh.u_clkbuf_out.u_buf  (.A(\u_skew_wh.d30 ),
    .X(net106));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_00.genblk1.u_mux  (.A0(\u_skew_wh.in0 ),
    .A1(\u_skew_wh.in1 ),
    .S(cfg_cska_wh[0]),
    .X(\u_skew_wh.d00 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_01.genblk1.u_mux  (.A0(\u_skew_wh.in2 ),
    .A1(\u_skew_wh.in3 ),
    .S(cfg_cska_wh[0]),
    .X(\u_skew_wh.d01 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_02.genblk1.u_mux  (.A0(\u_skew_wh.in4 ),
    .A1(\u_skew_wh.in5 ),
    .S(cfg_cska_wh[0]),
    .X(\u_skew_wh.d02 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_03.genblk1.u_mux  (.A0(\u_skew_wh.in6 ),
    .A1(\u_skew_wh.in7 ),
    .S(cfg_cska_wh[0]),
    .X(\u_skew_wh.d03 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_04.genblk1.u_mux  (.A0(\u_skew_wh.in8 ),
    .A1(\u_skew_wh.in9 ),
    .S(cfg_cska_wh[0]),
    .X(\u_skew_wh.d04 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_05.genblk1.u_mux  (.A0(\u_skew_wh.in10 ),
    .A1(\u_skew_wh.in11 ),
    .S(cfg_cska_wh[0]),
    .X(\u_skew_wh.d05 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_06.genblk1.u_mux  (.A0(\u_skew_wh.in12 ),
    .A1(\u_skew_wh.in13 ),
    .S(cfg_cska_wh[0]),
    .X(\u_skew_wh.d06 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_07.genblk1.u_mux  (.A0(\u_skew_wh.in14 ),
    .A1(\u_skew_wh.in15 ),
    .S(cfg_cska_wh[0]),
    .X(\u_skew_wh.d07 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_10.genblk1.u_mux  (.A0(\u_skew_wh.d00 ),
    .A1(\u_skew_wh.d01 ),
    .S(cfg_cska_wh[1]),
    .X(\u_skew_wh.d10 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_11.genblk1.u_mux  (.A0(\u_skew_wh.d02 ),
    .A1(\u_skew_wh.d03 ),
    .S(cfg_cska_wh[1]),
    .X(\u_skew_wh.d11 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_12.genblk1.u_mux  (.A0(\u_skew_wh.d04 ),
    .A1(\u_skew_wh.d05 ),
    .S(cfg_cska_wh[1]),
    .X(\u_skew_wh.d12 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_13.genblk1.u_mux  (.A0(\u_skew_wh.d06 ),
    .A1(\u_skew_wh.d07 ),
    .S(cfg_cska_wh[1]),
    .X(\u_skew_wh.d13 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_20.genblk1.u_mux  (.A0(\u_skew_wh.d10 ),
    .A1(\u_skew_wh.d11 ),
    .S(cfg_cska_wh[2]),
    .X(\u_skew_wh.d20 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_21.genblk1.u_mux  (.A0(\u_skew_wh.d12 ),
    .A1(\u_skew_wh.d13 ),
    .S(cfg_cska_wh[2]),
    .X(\u_skew_wh.d21 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_wh.u_mux_level_30.genblk1.u_mux  (.A0(\u_skew_wh.d20 ),
    .A1(\u_skew_wh.d21 ),
    .S(cfg_cska_wh[3]),
    .X(\u_skew_wh.d30 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_0.u_buf  (.A(\u_skew_wh.clk_inbuf ),
    .X(\u_skew_wh.in0 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_1.u_buf  (.A(\u_skew_wh.clk_d1 ),
    .X(\u_skew_wh.in1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_10.u_buf  (.A(net323),
    .X(\u_skew_wh.in10 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_11.u_buf  (.A(net322),
    .X(\u_skew_wh.in11 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_12.u_buf  (.A(\u_skew_wh.clk_d12 ),
    .X(\u_skew_wh.in12 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_13.u_buf  (.A(\u_skew_wh.clk_d13 ),
    .X(\u_skew_wh.in13 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_14.u_buf  (.A(\u_skew_wh.clk_d14 ),
    .X(\u_skew_wh.in14 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_15.u_buf  (.A(\u_skew_wh.clk_d15 ),
    .X(\u_skew_wh.in15 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_2.u_buf  (.A(\u_skew_wh.clk_d2 ),
    .X(\u_skew_wh.in2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_3.u_buf  (.A(\u_skew_wh.clk_d3 ),
    .X(\u_skew_wh.in3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_4.u_buf  (.A(\u_skew_wh.clk_d4 ),
    .X(\u_skew_wh.in4 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_5.u_buf  (.A(\u_skew_wh.clk_d5 ),
    .X(\u_skew_wh.in5 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_6.u_buf  (.A(\u_skew_wh.clk_d6 ),
    .X(\u_skew_wh.in6 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_7.u_buf  (.A(\u_skew_wh.clk_d7 ),
    .X(\u_skew_wh.in7 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_8.u_buf  (.A(\u_skew_wh.clk_d8 ),
    .X(\u_skew_wh.in8 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_wh.u_tap_9.u_buf  (.A(net321),
    .X(\u_skew_wh.in9 ));
 sky130_fd_sc_hd__mux2_1 \u_uart2wb.u_arst_sync.u_buf.genblk1.u_mux  (.A0(net339),
    .A1(net304),
    .S(net309),
    .X(\u_uart2wb.arst_ssn ));
 sky130_fd_sc_hd__conb_1 \u_uart2wb.u_arst_sync.u_buf.genblk1.u_mux_309  (.LO(net309));
 sky130_fd_sc_hd__mux2_1 \u_uart2wb.u_core.u_line_rst.u_buf.genblk1.u_mux  (.A0(\u_uart2wb.u_core.u_line_rst.in_data_2s ),
    .A1(net301),
    .S(net310),
    .X(\u_uart2wb.line_reset_n ));
 sky130_fd_sc_hd__conb_1 \u_uart2wb.u_core.u_line_rst.u_buf.genblk1.u_mux_310  (.LO(net310));
 sky130_fd_sc_hd__mux2_8 \u_uart2wb.u_core.u_uart_clk.genblk1.u_mux  (.A0(\u_uart2wb.u_core.line_clk_16x ),
    .A1(net311),
    .S(net312),
    .X(\u_uart2wb.baud_clk_16x ));
 sky130_fd_sc_hd__conb_1 \u_uart2wb.u_core.u_uart_clk.genblk1.u_mux_311  (.LO(net311));
 sky130_fd_sc_hd__conb_1 \u_uart2wb.u_core.u_uart_clk.genblk1.u_mux_312  (.LO(net312));
 sky130_fd_sc_hd__mux2_4 \u_wbm_rst.u_buf.genblk1.u_mux  (.A0(net349),
    .A1(\u_wbm_rst.arst_n ),
    .S(net313),
    .X(net68));
 sky130_fd_sc_hd__conb_1 \u_wbm_rst.u_buf.genblk1.u_mux_313  (.LO(net313));
 sky130_fd_sc_hd__mux2_1 \u_wbs_rst.u_buf.genblk1.u_mux  (.A0(net338),
    .A1(net303),
    .S(net314),
    .X(\u_async_wb.u_cmd_if.rd_reset_n ));
 sky130_fd_sc_hd__conb_1 \u_wbs_rst.u_buf.genblk1.u_mux_314  (.LO(net314));
 sky130_fd_sc_hd__buf_2 wire1 (.A(wbm_clk_i),
    .X(net320));
 sky130_fd_sc_hd__buf_4 wire215 (.A(_02257_),
    .X(net215));
 sky130_fd_sc_hd__buf_4 wire216 (.A(_02252_),
    .X(net216));
 sky130_fd_sc_hd__buf_4 wire217 (.A(_02232_),
    .X(net217));
 sky130_fd_sc_hd__buf_4 wire218 (.A(_02226_),
    .X(net218));
 sky130_fd_sc_hd__buf_4 wire219 (.A(_02209_),
    .X(net219));
 sky130_fd_sc_hd__buf_4 wire220 (.A(_02198_),
    .X(net220));
 sky130_fd_sc_hd__buf_4 wire221 (.A(_02190_),
    .X(net221));
 sky130_fd_sc_hd__buf_4 wire222 (.A(_02185_),
    .X(net222));
 sky130_fd_sc_hd__buf_4 wire223 (.A(_02179_),
    .X(net223));
 sky130_fd_sc_hd__buf_4 wire224 (.A(_02153_),
    .X(net224));
 sky130_fd_sc_hd__buf_4 wire225 (.A(_02284_),
    .X(net225));
 sky130_fd_sc_hd__buf_4 wire226 (.A(_02264_),
    .X(net226));
 sky130_fd_sc_hd__buf_4 wire227 (.A(_02244_),
    .X(net227));
 sky130_fd_sc_hd__buf_4 wire228 (.A(_02237_),
    .X(net228));
 sky130_fd_sc_hd__buf_4 wire229 (.A(_02204_),
    .X(net229));
 sky130_fd_sc_hd__buf_4 wire306 (.A(user_clock2),
    .X(net306));
 sky130_fd_sc_hd__buf_6 wire307 (.A(user_clock1),
    .X(net307));
 sky130_fd_sc_hd__buf_4 wire308 (.A(sdin),
    .X(net308));
endmodule

