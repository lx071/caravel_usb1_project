magic
tech sky130A
magscale 1 2
timestamp 1698825809
<< viali >>
rect 218805 9605 218839 9639
rect 221381 9605 221415 9639
rect 225613 9605 225647 9639
rect 340153 9605 340187 9639
rect 342729 9605 342763 9639
rect 345305 9605 345339 9639
rect 352757 9605 352791 9639
rect 354505 9605 354539 9639
rect 366097 9605 366131 9639
rect 368581 9605 368615 9639
rect 384037 9605 384071 9639
rect 183293 9537 183327 9571
rect 184397 9537 184431 9571
rect 190837 9537 190871 9571
rect 195253 9537 195287 9571
rect 195897 9537 195931 9571
rect 198381 9537 198415 9571
rect 202981 9537 203015 9571
rect 203625 9537 203659 9571
rect 205741 9537 205775 9571
rect 206293 9537 206327 9571
rect 210525 9537 210559 9571
rect 211077 9537 211111 9571
rect 213285 9537 213319 9571
rect 213837 9537 213871 9571
rect 218253 9537 218287 9571
rect 220829 9537 220863 9571
rect 224969 9537 225003 9571
rect 228557 9537 228591 9571
rect 232513 9537 232547 9571
rect 236285 9537 236319 9571
rect 239965 9537 239999 9571
rect 244013 9537 244047 9571
rect 339509 9537 339543 9571
rect 342085 9537 342119 9571
rect 344661 9537 344695 9571
rect 346777 9537 346811 9571
rect 347053 9537 347087 9571
rect 347605 9537 347639 9571
rect 349629 9537 349663 9571
rect 352205 9537 352239 9571
rect 354781 9537 354815 9571
rect 357357 9537 357391 9571
rect 358645 9537 358679 9571
rect 358921 9537 358955 9571
rect 359565 9537 359599 9571
rect 361497 9537 361531 9571
rect 363981 9537 364015 9571
rect 366373 9537 366407 9571
rect 368857 9537 368891 9571
rect 371341 9537 371375 9571
rect 373733 9537 373767 9571
rect 376217 9537 376251 9571
rect 378609 9537 378643 9571
rect 381093 9537 381127 9571
rect 383485 9537 383519 9571
rect 182741 9469 182775 9503
rect 190285 9469 190319 9503
rect 194701 9469 194735 9503
rect 197829 9469 197863 9503
rect 202429 9469 202463 9503
rect 205465 9469 205499 9503
rect 210249 9469 210283 9503
rect 213009 9469 213043 9503
rect 217977 9469 218011 9503
rect 220553 9469 220587 9503
rect 224693 9469 224727 9503
rect 228281 9469 228315 9503
rect 232237 9469 232271 9503
rect 236009 9469 236043 9503
rect 236837 9469 236871 9503
rect 239689 9469 239723 9503
rect 243737 9469 243771 9503
rect 338957 9469 338991 9503
rect 341533 9469 341567 9503
rect 344109 9469 344143 9503
rect 349353 9469 349387 9503
rect 351929 9469 351963 9503
rect 357081 9469 357115 9503
rect 361221 9469 361255 9503
rect 362141 9469 362175 9503
rect 363705 9469 363739 9503
rect 364717 9469 364751 9503
rect 371065 9469 371099 9503
rect 373457 9469 373491 9503
rect 375941 9469 375975 9503
rect 378333 9469 378367 9503
rect 380817 9469 380851 9503
rect 383209 9469 383243 9503
rect 233341 9401 233375 9435
rect 381645 9401 381679 9435
rect 191481 9333 191515 9367
rect 199025 9333 199059 9367
rect 229109 9333 229143 9367
rect 244565 9333 244599 9367
rect 350089 9333 350123 9367
rect 355333 9333 355367 9367
rect 357909 9333 357943 9367
rect 367293 9333 367327 9367
rect 369869 9333 369903 9367
rect 374285 9333 374319 9367
rect 376769 9333 376803 9367
rect 379161 9333 379195 9367
rect 240149 8993 240183 9027
rect 152749 8925 152783 8959
rect 160477 8925 160511 8959
rect 161029 8925 161063 8959
rect 168113 8925 168147 8959
rect 172437 8925 172471 8959
rect 173081 8925 173115 8959
rect 175657 8925 175691 8959
rect 176301 8925 176335 8959
rect 179981 8925 180015 8959
rect 180533 8925 180567 8959
rect 187617 8925 187651 8959
rect 321293 8925 321327 8959
rect 321845 8925 321879 8959
rect 322489 8925 322523 8959
rect 326353 8925 326387 8959
rect 326905 8925 326939 8959
rect 331873 8925 331907 8959
rect 332517 8925 332551 8959
rect 336289 8925 336323 8959
rect 336841 8925 336875 8959
rect 337485 8925 337519 8959
rect 152197 8857 152231 8891
rect 160109 8857 160143 8891
rect 167561 8857 167595 8891
rect 171885 8857 171919 8891
rect 175289 8857 175323 8891
rect 179429 8857 179463 8891
rect 187065 8857 187099 8891
rect 331321 8857 331355 8891
rect 153485 8789 153519 8823
rect 168941 8789 168975 8823
rect 188261 8789 188295 8823
rect 327549 8789 327583 8823
rect 371525 8789 371559 8823
rect 302433 8585 302467 8619
rect 307493 8585 307527 8619
rect 312461 8585 312495 8619
rect 144469 8517 144503 8551
rect 145757 8517 145791 8551
rect 164341 8517 164375 8551
rect 142077 8449 142111 8483
rect 145021 8449 145055 8483
rect 149713 8449 149747 8483
rect 157257 8449 157291 8483
rect 157901 8449 157935 8483
rect 164893 8449 164927 8483
rect 165537 8449 165571 8483
rect 301789 8449 301823 8483
rect 306389 8449 306423 8483
rect 306849 8449 306883 8483
rect 311265 8449 311299 8483
rect 311817 8449 311851 8483
rect 316325 8449 316359 8483
rect 316877 8449 316911 8483
rect 317521 8449 317555 8483
rect 141525 8381 141559 8415
rect 142721 8381 142755 8415
rect 149161 8381 149195 8415
rect 156705 8381 156739 8415
rect 301237 8381 301271 8415
rect 101045 8041 101079 8075
rect 122573 8041 122607 8075
rect 277133 8041 277167 8075
rect 282285 8041 282319 8075
rect 287437 8041 287471 8075
rect 292589 8041 292623 8075
rect 276029 7905 276063 7939
rect 91661 7837 91695 7871
rect 92305 7837 92339 7871
rect 96721 7837 96755 7871
rect 114201 7837 114235 7871
rect 121837 7837 121871 7871
rect 126897 7837 126931 7871
rect 131957 7837 131991 7871
rect 137017 7837 137051 7871
rect 138029 7837 138063 7871
rect 149897 7837 149931 7871
rect 276397 7837 276431 7871
rect 281549 7837 281583 7871
rect 286701 7837 286735 7871
rect 291761 7837 291795 7871
rect 296729 7837 296763 7871
rect 297741 7837 297775 7871
rect 92857 7769 92891 7803
rect 113649 7769 113683 7803
rect 121285 7769 121319 7803
rect 126345 7769 126379 7803
rect 131405 7769 131439 7803
rect 136649 7769 136683 7803
rect 280997 7769 281031 7803
rect 286149 7769 286183 7803
rect 291209 7769 291243 7803
rect 296177 7769 296211 7803
rect 94053 7701 94087 7735
rect 95249 7701 95283 7735
rect 97641 7701 97675 7735
rect 114845 7701 114879 7735
rect 127725 7701 127759 7735
rect 132877 7701 132911 7735
rect 251373 7701 251407 7735
rect 252477 7701 252511 7735
rect 256985 7497 257019 7531
rect 262045 7497 262079 7531
rect 267105 7497 267139 7531
rect 272165 7497 272199 7531
rect 96077 7429 96111 7463
rect 97273 7429 97307 7463
rect 98469 7429 98503 7463
rect 101873 7429 101907 7463
rect 250821 7429 250855 7463
rect 91201 7361 91235 7395
rect 91753 7361 91787 7395
rect 92949 7361 92983 7395
rect 93501 7361 93535 7395
rect 94329 7361 94363 7395
rect 95525 7361 95559 7395
rect 96721 7361 96755 7395
rect 97917 7361 97951 7395
rect 99481 7361 99515 7395
rect 100125 7361 100159 7395
rect 100677 7361 100711 7395
rect 101321 7361 101355 7395
rect 250269 7361 250303 7395
rect 251465 7361 251499 7395
rect 252661 7361 252695 7395
rect 254225 7361 254259 7395
rect 254777 7361 254811 7395
rect 256341 7361 256375 7395
rect 260849 7361 260883 7395
rect 261401 7361 261435 7395
rect 266461 7361 266495 7395
rect 270969 7361 271003 7395
rect 271521 7361 271555 7395
rect 94881 7293 94915 7327
rect 252017 7293 252051 7327
rect 253213 7293 253247 7327
rect 255789 7293 255823 7327
rect 265909 7293 265943 7327
rect 90557 7157 90591 7191
rect 92305 7157 92339 7191
rect 103253 7157 103287 7191
rect 113373 7157 113407 7191
rect 249625 7157 249659 7191
rect 124965 6885 124999 6919
rect 102885 6817 102919 6851
rect 104081 6817 104115 6851
rect 105277 6817 105311 6851
rect 108589 6817 108623 6851
rect 112821 6817 112855 6851
rect 115397 6817 115431 6851
rect 258365 6817 258399 6851
rect 259561 6817 259595 6851
rect 91661 6749 91695 6783
rect 92121 6749 92155 6783
rect 93409 6749 93443 6783
rect 93777 6749 93811 6783
rect 94605 6749 94639 6783
rect 95157 6749 95191 6783
rect 96905 6749 96939 6783
rect 97457 6749 97491 6783
rect 99021 6749 99055 6783
rect 102333 6749 102367 6783
rect 103529 6749 103563 6783
rect 104725 6749 104759 6783
rect 108037 6749 108071 6783
rect 110337 6749 110371 6783
rect 112269 6749 112303 6783
rect 113649 6749 113683 6783
rect 114845 6749 114879 6783
rect 117421 6749 117455 6783
rect 251925 6749 251959 6783
rect 255237 6749 255271 6783
rect 256617 6749 256651 6783
rect 257813 6749 257847 6783
rect 259009 6749 259043 6783
rect 260205 6749 260239 6783
rect 99573 6681 99607 6715
rect 107485 6681 107519 6715
rect 110889 6681 110923 6715
rect 114201 6681 114235 6715
rect 117973 6681 118007 6715
rect 251373 6681 251407 6715
rect 255789 6681 255823 6715
rect 257169 6681 257203 6715
rect 260757 6681 260791 6715
rect 90925 6613 90959 6647
rect 92765 6613 92799 6647
rect 98377 6613 98411 6647
rect 101229 6613 101263 6647
rect 109693 6613 109727 6647
rect 111533 6613 111567 6647
rect 116685 6613 116719 6647
rect 120273 6613 120307 6647
rect 121469 6613 121503 6647
rect 252569 6613 252603 6647
rect 253949 6613 253983 6647
rect 254593 6613 254627 6647
rect 99941 6341 99975 6375
rect 101965 6341 101999 6375
rect 106197 6341 106231 6375
rect 107485 6341 107519 6375
rect 110981 6341 111015 6375
rect 122205 6341 122239 6375
rect 124413 6341 124447 6375
rect 261953 6341 261987 6375
rect 266829 6341 266863 6375
rect 99389 6273 99423 6307
rect 101413 6273 101447 6307
rect 103253 6273 103287 6307
rect 105737 6273 105771 6307
rect 106933 6273 106967 6307
rect 108037 6273 108071 6307
rect 110429 6273 110463 6307
rect 112361 6273 112395 6307
rect 112913 6273 112947 6307
rect 113557 6273 113591 6307
rect 118249 6273 118283 6307
rect 120457 6273 120491 6307
rect 121009 6273 121043 6307
rect 121653 6273 121687 6307
rect 123861 6273 123895 6307
rect 125149 6273 125183 6307
rect 125517 6273 125551 6307
rect 127265 6273 127299 6307
rect 127817 6273 127851 6307
rect 128461 6273 128495 6307
rect 261401 6273 261435 6307
rect 262597 6273 262631 6307
rect 264989 6273 265023 6307
rect 266277 6273 266311 6307
rect 103805 6205 103839 6239
rect 114109 6205 114143 6239
rect 118525 6205 118559 6239
rect 129013 6205 129047 6239
rect 263149 6205 263183 6239
rect 265541 6205 265575 6239
rect 98653 6137 98687 6171
rect 94329 6069 94363 6103
rect 96721 6069 96755 6103
rect 100769 6069 100803 6103
rect 102609 6069 102643 6103
rect 104449 6069 104483 6103
rect 105093 6069 105127 6103
rect 109785 6069 109819 6103
rect 111809 6069 111843 6103
rect 114753 6069 114787 6103
rect 117605 6069 117639 6103
rect 123217 6069 123251 6103
rect 126621 6069 126655 6103
rect 131681 6069 131715 6103
rect 256341 6069 256375 6103
rect 257537 6069 257571 6103
rect 259009 6069 259043 6103
rect 259929 6069 259963 6103
rect 260849 6069 260883 6103
rect 264345 6069 264379 6103
rect 107577 5729 107611 5763
rect 116685 5729 116719 5763
rect 121285 5729 121319 5763
rect 124689 5729 124723 5763
rect 135545 5729 135579 5763
rect 264345 5729 264379 5763
rect 269129 5729 269163 5763
rect 106381 5661 106415 5695
rect 107117 5661 107151 5695
rect 109325 5661 109359 5695
rect 109877 5661 109911 5695
rect 116133 5661 116167 5695
rect 117421 5661 117455 5695
rect 117973 5661 118007 5695
rect 119537 5661 119571 5695
rect 120733 5661 120767 5695
rect 122941 5661 122975 5695
rect 123493 5661 123527 5695
rect 124137 5661 124171 5695
rect 130669 5661 130703 5695
rect 130945 5661 130979 5695
rect 131773 5661 131807 5695
rect 132049 5661 132083 5695
rect 134165 5661 134199 5695
rect 134441 5661 134475 5695
rect 135269 5661 135303 5695
rect 138765 5661 138799 5695
rect 263793 5661 263827 5695
rect 266829 5661 266863 5695
rect 267473 5661 267507 5695
rect 268669 5661 268703 5695
rect 269957 5661 269991 5695
rect 120089 5593 120123 5627
rect 139041 5593 139075 5627
rect 268025 5593 268059 5627
rect 270509 5593 270543 5627
rect 108681 5525 108715 5559
rect 113281 5525 113315 5559
rect 115489 5525 115523 5559
rect 118893 5525 118927 5559
rect 128185 5525 128219 5559
rect 130117 5525 130151 5559
rect 133613 5525 133647 5559
rect 138213 5525 138247 5559
rect 141985 5525 142019 5559
rect 262321 5525 262355 5559
rect 263149 5525 263183 5559
rect 266001 5525 266035 5559
rect 126897 5253 126931 5287
rect 134625 5253 134659 5287
rect 126345 5185 126379 5219
rect 127541 5185 127575 5219
rect 130301 5185 130335 5219
rect 131405 5185 131439 5219
rect 133245 5185 133279 5219
rect 134349 5185 134383 5219
rect 137569 5185 137603 5219
rect 141065 5185 141099 5219
rect 141341 5185 141375 5219
rect 142169 5185 142203 5219
rect 144561 5185 144595 5219
rect 145665 5185 145699 5219
rect 145941 5185 145975 5219
rect 148057 5185 148091 5219
rect 271153 5185 271187 5219
rect 117145 5117 117179 5151
rect 128093 5117 128127 5151
rect 130853 5117 130887 5151
rect 131681 5117 131715 5151
rect 133521 5117 133555 5151
rect 137845 5117 137879 5151
rect 142445 5117 142479 5151
rect 144837 5117 144871 5151
rect 148333 5117 148367 5151
rect 271705 5117 271739 5151
rect 123861 5049 123895 5083
rect 120457 4981 120491 5015
rect 122757 4981 122791 5015
rect 125701 4981 125735 5015
rect 129565 4981 129599 5015
rect 132693 4981 132727 5015
rect 135361 4981 135395 5015
rect 137017 4981 137051 5015
rect 140513 4981 140547 5015
rect 144009 4981 144043 5015
rect 147505 4981 147539 5015
rect 268393 4981 268427 5015
rect 269681 4981 269715 5015
rect 270601 4981 270635 5015
rect 137017 4641 137051 4675
rect 138213 4641 138247 4675
rect 136741 4573 136775 4607
rect 137937 4573 137971 4607
rect 140237 4573 140271 4607
rect 141341 4573 141375 4607
rect 149161 4573 149195 4607
rect 149437 4573 149471 4607
rect 131221 4505 131255 4539
rect 139685 4505 139719 4539
rect 140513 4505 140547 4539
rect 141617 4505 141651 4539
rect 127633 4437 127667 4471
rect 134165 4437 134199 4471
rect 136189 4437 136223 4471
rect 145481 4437 145515 4471
rect 137753 4097 137787 4131
rect 143733 4097 143767 4131
rect 145665 4097 145699 4131
rect 147229 4097 147263 4131
rect 148425 4097 148459 4131
rect 150817 4097 150851 4131
rect 144009 4029 144043 4063
rect 145941 4029 145975 4063
rect 147505 4029 147539 4063
rect 148701 4029 148735 4063
rect 151093 4029 151127 4063
rect 143181 3961 143215 3995
rect 141157 3893 141191 3927
rect 145021 3893 145055 3927
rect 146677 3893 146711 3927
rect 1869 3689 1903 3723
rect 4445 3689 4479 3723
rect 6837 3689 6871 3723
rect 9597 3689 9631 3723
rect 12173 3689 12207 3723
rect 14749 3689 14783 3723
rect 17325 3689 17359 3723
rect 19901 3689 19935 3723
rect 22477 3689 22511 3723
rect 30205 3689 30239 3723
rect 36093 3689 36127 3723
rect 43821 3689 43855 3723
rect 45661 3689 45695 3723
rect 48237 3689 48271 3723
rect 59277 3689 59311 3723
rect 66269 3689 66303 3723
rect 67005 3689 67039 3723
rect 68845 3689 68879 3723
rect 122941 3689 122975 3723
rect 130853 3689 130887 3723
rect 35357 3621 35391 3655
rect 40509 3621 40543 3655
rect 61117 3621 61151 3655
rect 63693 3621 63727 3655
rect 109969 3621 110003 3655
rect 115121 3621 115155 3655
rect 117697 3621 117731 3655
rect 125425 3621 125459 3655
rect 133429 3621 133463 3655
rect 135821 3621 135855 3655
rect 24869 3553 24903 3587
rect 37749 3553 37783 3587
rect 113373 3553 113407 3587
rect 148241 3553 148275 3587
rect 31953 3485 31987 3519
rect 32873 3485 32907 3519
rect 35541 3485 35575 3519
rect 40693 3485 40727 3519
rect 43269 3485 43303 3519
rect 45845 3485 45879 3519
rect 48421 3485 48455 3519
rect 50997 3485 51031 3519
rect 53573 3485 53607 3519
rect 56149 3485 56183 3519
rect 58725 3485 58759 3519
rect 61301 3485 61335 3519
rect 63877 3485 63911 3519
rect 66453 3485 66487 3519
rect 69029 3485 69063 3519
rect 71605 3485 71639 3519
rect 74181 3485 74215 3519
rect 74733 3485 74767 3519
rect 81909 3485 81943 3519
rect 89637 3485 89671 3519
rect 90189 3485 90223 3519
rect 97365 3485 97399 3519
rect 105093 3485 105127 3519
rect 112821 3485 112855 3519
rect 120549 3485 120583 3519
rect 128277 3485 128311 3519
rect 130669 3485 130703 3519
rect 131313 3485 131347 3519
rect 133245 3485 133279 3519
rect 133889 3485 133923 3519
rect 136005 3485 136039 3519
rect 136557 3485 136591 3519
rect 1961 3417 1995 3451
rect 4537 3417 4571 3451
rect 7113 3417 7147 3451
rect 9689 3417 9723 3451
rect 12265 3417 12299 3451
rect 14841 3417 14875 3451
rect 17417 3417 17451 3451
rect 19993 3417 20027 3451
rect 22569 3417 22603 3451
rect 25145 3417 25179 3451
rect 26893 3417 26927 3451
rect 27721 3417 27755 3451
rect 30297 3417 30331 3451
rect 37105 3417 37139 3451
rect 38025 3417 38059 3451
rect 47593 3417 47627 3451
rect 76481 3417 76515 3451
rect 76665 3417 76699 3451
rect 79057 3417 79091 3451
rect 79241 3417 79275 3451
rect 82461 3417 82495 3451
rect 84393 3417 84427 3451
rect 86969 3417 87003 3451
rect 92121 3417 92155 3451
rect 94697 3417 94731 3451
rect 99849 3417 99883 3451
rect 102425 3417 102459 3451
rect 105645 3417 105679 3451
rect 107577 3417 107611 3451
rect 110153 3417 110187 3451
rect 115305 3417 115339 3451
rect 117881 3417 117915 3451
rect 123033 3417 123067 3451
rect 125609 3417 125643 3451
rect 128829 3417 128863 3451
rect 6193 3349 6227 3383
rect 11345 3349 11379 3383
rect 16589 3349 16623 3383
rect 21649 3349 21683 3383
rect 27629 3349 27663 3383
rect 32781 3349 32815 3383
rect 43085 3349 43119 3383
rect 50813 3349 50847 3383
rect 51549 3349 51583 3383
rect 52745 3349 52779 3383
rect 53389 3349 53423 3383
rect 55965 3349 55999 3383
rect 58541 3349 58575 3383
rect 63049 3349 63083 3383
rect 68201 3349 68235 3383
rect 71421 3349 71455 3383
rect 73997 3349 74031 3383
rect 78505 3349 78539 3383
rect 81725 3349 81759 3383
rect 83657 3349 83691 3383
rect 84301 3349 84335 3383
rect 86877 3349 86911 3383
rect 89453 3349 89487 3383
rect 92029 3349 92063 3383
rect 93961 3349 93995 3383
rect 94605 3349 94639 3383
rect 97181 3349 97215 3383
rect 97917 3349 97951 3383
rect 99113 3349 99147 3383
rect 99757 3349 99791 3383
rect 102333 3349 102367 3383
rect 104909 3349 104943 3383
rect 107485 3349 107519 3383
rect 109417 3349 109451 3383
rect 112637 3349 112671 3383
rect 114569 3349 114603 3383
rect 120365 3349 120399 3383
rect 121101 3349 121135 3383
rect 124873 3349 124907 3383
rect 128093 3349 128127 3383
rect 485881 3145 485915 3179
rect 488549 3145 488583 3179
rect 491033 3145 491067 3179
rect 493609 3145 493643 3179
rect 496185 3145 496219 3179
rect 498761 3145 498795 3179
rect 501337 3145 501371 3179
rect 503913 3145 503947 3179
rect 506489 3145 506523 3179
rect 509065 3145 509099 3179
rect 511641 3145 511675 3179
rect 71237 3077 71271 3111
rect 107209 3009 107243 3043
rect 117605 3009 117639 3043
rect 40233 2873 40267 2907
rect 45385 2873 45419 2907
rect 76297 2873 76331 2907
rect 86601 2873 86635 2907
rect 194609 2873 194643 2907
rect 1593 2805 1627 2839
rect 3985 2805 4019 2839
rect 6561 2805 6595 2839
rect 9137 2805 9171 2839
rect 14289 2805 14323 2839
rect 19441 2805 19475 2839
rect 24593 2805 24627 2839
rect 29745 2805 29779 2839
rect 34897 2805 34931 2839
rect 37473 2805 37507 2839
rect 42809 2805 42843 2839
rect 50537 2805 50571 2839
rect 53113 2805 53147 2839
rect 55689 2805 55723 2839
rect 58265 2805 58299 2839
rect 60841 2805 60875 2839
rect 65993 2805 66027 2839
rect 68569 2805 68603 2839
rect 73721 2805 73755 2839
rect 81449 2805 81483 2839
rect 84025 2805 84059 2839
rect 89269 2805 89303 2839
rect 91753 2805 91787 2839
rect 96905 2805 96939 2839
rect 99481 2805 99515 2839
rect 102149 2805 102183 2839
rect 104633 2805 104667 2839
rect 112361 2805 112395 2839
rect 115029 2805 115063 2839
rect 120089 2805 120123 2839
rect 122665 2805 122699 2839
rect 127909 2805 127943 2839
rect 138029 2805 138063 2839
rect 143089 2805 143123 2839
rect 148241 2805 148275 2839
rect 153393 2805 153427 2839
rect 158545 2805 158579 2839
rect 163697 2805 163731 2839
rect 168849 2805 168883 2839
rect 174001 2805 174035 2839
rect 179153 2805 179187 2839
rect 184305 2805 184339 2839
rect 189457 2805 189491 2839
rect 200037 2805 200071 2839
rect 205097 2805 205131 2839
rect 210249 2805 210283 2839
rect 215401 2805 215435 2839
rect 220553 2805 220587 2839
rect 225797 2805 225831 2839
rect 514217 2805 514251 2839
rect 5181 2601 5215 2635
rect 9597 2601 9631 2635
rect 61117 2601 61151 2635
rect 68845 2601 68879 2635
rect 73997 2601 74031 2635
rect 76573 2601 76607 2635
rect 81725 2601 81759 2635
rect 87613 2601 87647 2635
rect 92029 2601 92063 2635
rect 97181 2601 97215 2635
rect 102333 2601 102367 2635
rect 103069 2601 103103 2635
rect 110061 2601 110095 2635
rect 110797 2601 110831 2635
rect 112637 2601 112671 2635
rect 141709 2601 141743 2635
rect 192493 2601 192527 2635
rect 193229 2601 193263 2635
rect 205373 2601 205407 2635
rect 208593 2601 208627 2635
rect 210525 2601 210559 2635
rect 224141 2601 224175 2635
rect 229201 2601 229235 2635
rect 231869 2601 231903 2635
rect 234445 2601 234479 2635
rect 237021 2601 237055 2635
rect 242173 2601 242207 2635
rect 244749 2601 244783 2635
rect 247233 2601 247267 2635
rect 249901 2601 249935 2635
rect 257629 2601 257663 2635
rect 260205 2601 260239 2635
rect 265357 2601 265391 2635
rect 270509 2601 270543 2635
rect 273085 2601 273119 2635
rect 275661 2601 275695 2635
rect 280813 2601 280847 2635
rect 283389 2601 283423 2635
rect 285965 2601 285999 2635
rect 288541 2601 288575 2635
rect 291117 2601 291151 2635
rect 293693 2601 293727 2635
rect 296269 2601 296303 2635
rect 298845 2601 298879 2635
rect 301421 2601 301455 2635
rect 303261 2601 303295 2635
rect 303997 2601 304031 2635
rect 306573 2601 306607 2635
rect 309149 2601 309183 2635
rect 316877 2601 316911 2635
rect 322029 2601 322063 2635
rect 327181 2601 327215 2635
rect 360669 2601 360703 2635
rect 365085 2601 365119 2635
rect 365821 2601 365855 2635
rect 370237 2601 370271 2635
rect 376125 2601 376159 2635
rect 378701 2601 378735 2635
rect 385693 2601 385727 2635
rect 390845 2601 390879 2635
rect 399309 2601 399343 2635
rect 412189 2601 412223 2635
rect 450829 2601 450863 2635
rect 453405 2601 453439 2635
rect 466285 2601 466319 2635
rect 484317 2601 484351 2635
rect 12909 2533 12943 2567
rect 18061 2533 18095 2567
rect 19809 2533 19843 2567
rect 43085 2533 43119 2567
rect 45661 2533 45695 2567
rect 107393 2533 107427 2567
rect 117789 2533 117823 2567
rect 118525 2533 118559 2567
rect 177773 2533 177807 2567
rect 182925 2533 182959 2567
rect 184673 2533 184707 2567
rect 290381 2533 290415 2567
rect 295533 2533 295567 2567
rect 300685 2533 300719 2567
rect 308413 2533 308447 2567
rect 313565 2533 313599 2567
rect 334909 2533 334943 2567
rect 347789 2533 347823 2567
rect 349629 2533 349663 2567
rect 355517 2533 355551 2567
rect 367661 2533 367695 2567
rect 375389 2533 375423 2567
rect 388269 2533 388303 2567
rect 393421 2533 393455 2567
rect 395997 2533 396031 2567
rect 398573 2533 398607 2567
rect 404369 2533 404403 2567
rect 414765 2533 414799 2567
rect 419917 2533 419951 2567
rect 425069 2533 425103 2567
rect 430221 2533 430255 2567
rect 434637 2533 434671 2567
rect 435373 2533 435407 2567
rect 439789 2533 439823 2567
rect 457821 2533 457855 2567
rect 461133 2533 461167 2567
rect 1685 2465 1719 2499
rect 33517 2465 33551 2499
rect 41245 2465 41279 2499
rect 136465 2465 136499 2499
rect 153853 2465 153887 2499
rect 311725 2465 311759 2499
rect 352941 2465 352975 2499
rect 373549 2465 373583 2499
rect 401885 2465 401919 2499
rect 437949 2465 437983 2499
rect 445677 2465 445711 2499
rect 476589 2465 476623 2499
rect 481741 2465 481775 2499
rect 4629 2397 4663 2431
rect 8493 2397 8527 2431
rect 9689 2397 9723 2431
rect 12357 2397 12391 2431
rect 17509 2397 17543 2431
rect 22661 2397 22695 2431
rect 27813 2397 27847 2431
rect 32965 2397 32999 2431
rect 40693 2397 40727 2431
rect 43269 2397 43303 2431
rect 45845 2397 45879 2431
rect 48421 2397 48455 2431
rect 48973 2397 49007 2431
rect 50997 2397 51031 2431
rect 53573 2397 53607 2431
rect 56149 2397 56183 2431
rect 56609 2397 56643 2431
rect 58725 2397 58759 2431
rect 61301 2397 61335 2431
rect 63877 2397 63911 2431
rect 66453 2397 66487 2431
rect 69029 2397 69063 2431
rect 71605 2397 71639 2431
rect 74181 2397 74215 2431
rect 79333 2397 79367 2431
rect 87061 2397 87095 2431
rect 89361 2397 89395 2431
rect 94789 2397 94823 2431
rect 95341 2397 95375 2431
rect 102517 2397 102551 2431
rect 110245 2397 110279 2431
rect 117973 2397 118007 2431
rect 121837 2397 121871 2431
rect 123033 2397 123067 2431
rect 125701 2397 125735 2431
rect 130669 2397 130703 2431
rect 131313 2397 131347 2431
rect 133429 2397 133463 2431
rect 135821 2397 135855 2431
rect 138581 2397 138615 2431
rect 141157 2397 141191 2431
rect 143733 2397 143767 2431
rect 146309 2397 146343 2431
rect 148885 2397 148919 2431
rect 151461 2397 151495 2431
rect 154037 2397 154071 2431
rect 156613 2397 156647 2431
rect 158913 2397 158947 2431
rect 159189 2397 159223 2431
rect 161765 2397 161799 2431
rect 166917 2397 166951 2431
rect 172069 2397 172103 2431
rect 177221 2397 177255 2431
rect 179705 2397 179739 2431
rect 182373 2397 182407 2431
rect 187525 2397 187559 2431
rect 188077 2397 188111 2431
rect 192677 2397 192711 2431
rect 195161 2397 195195 2431
rect 197829 2397 197863 2431
rect 198289 2397 198323 2431
rect 200405 2397 200439 2431
rect 202981 2397 203015 2431
rect 203441 2397 203475 2431
rect 205557 2397 205591 2431
rect 208133 2397 208167 2431
rect 210709 2397 210743 2431
rect 213285 2397 213319 2431
rect 213745 2397 213779 2431
rect 215861 2397 215895 2431
rect 218437 2397 218471 2431
rect 218897 2397 218931 2431
rect 221013 2397 221047 2431
rect 223589 2397 223623 2431
rect 228741 2397 228775 2431
rect 231317 2397 231351 2431
rect 233893 2397 233927 2431
rect 236469 2397 236503 2431
rect 239045 2397 239079 2431
rect 239505 2397 239539 2431
rect 241621 2397 241655 2431
rect 244197 2397 244231 2431
rect 246773 2397 246807 2431
rect 249349 2397 249383 2431
rect 251925 2397 251959 2431
rect 252385 2397 252419 2431
rect 254501 2397 254535 2431
rect 257077 2397 257111 2431
rect 259653 2397 259687 2431
rect 262229 2397 262263 2431
rect 262689 2397 262723 2431
rect 264805 2397 264839 2431
rect 267381 2397 267415 2431
rect 269957 2397 269991 2431
rect 272533 2397 272567 2431
rect 275109 2397 275143 2431
rect 277685 2397 277719 2431
rect 280261 2397 280295 2431
rect 282837 2397 282871 2431
rect 285413 2397 285447 2431
rect 287989 2397 288023 2431
rect 290565 2397 290599 2431
rect 293141 2397 293175 2431
rect 295717 2397 295751 2431
rect 298293 2397 298327 2431
rect 300869 2397 300903 2431
rect 303445 2397 303479 2431
rect 306021 2397 306055 2431
rect 308597 2397 308631 2431
rect 311173 2397 311207 2431
rect 313749 2397 313783 2431
rect 316325 2397 316359 2431
rect 318901 2397 318935 2431
rect 321477 2397 321511 2431
rect 324053 2397 324087 2431
rect 326629 2397 326663 2431
rect 329205 2397 329239 2431
rect 331781 2397 331815 2431
rect 334357 2397 334391 2431
rect 336933 2397 336967 2431
rect 339509 2397 339543 2431
rect 342085 2397 342119 2431
rect 344661 2397 344695 2431
rect 347237 2397 347271 2431
rect 349813 2397 349847 2431
rect 352389 2397 352423 2431
rect 354965 2397 354999 2431
rect 357541 2397 357575 2431
rect 360117 2397 360151 2431
rect 362693 2397 362727 2431
rect 365269 2397 365303 2431
rect 367845 2397 367879 2431
rect 370421 2397 370455 2431
rect 372997 2397 373031 2431
rect 375573 2397 375607 2431
rect 378149 2397 378183 2431
rect 380725 2397 380759 2431
rect 383301 2397 383335 2431
rect 385877 2397 385911 2431
rect 388453 2397 388487 2431
rect 391029 2397 391063 2431
rect 393605 2397 393639 2431
rect 394157 2397 394191 2431
rect 396181 2397 396215 2431
rect 396733 2397 396767 2431
rect 398757 2397 398791 2431
rect 401333 2397 401367 2431
rect 403909 2397 403943 2431
rect 406485 2397 406519 2431
rect 409061 2397 409095 2431
rect 411637 2397 411671 2431
rect 414213 2397 414247 2431
rect 416789 2397 416823 2431
rect 419365 2397 419399 2431
rect 421941 2397 421975 2431
rect 424517 2397 424551 2431
rect 427093 2397 427127 2431
rect 429669 2397 429703 2431
rect 432245 2397 432279 2431
rect 434821 2397 434855 2431
rect 437397 2397 437431 2431
rect 439973 2397 440007 2431
rect 442549 2397 442583 2431
rect 445125 2397 445159 2431
rect 447701 2397 447735 2431
rect 450277 2397 450311 2431
rect 452853 2397 452887 2431
rect 455429 2397 455463 2431
rect 455981 2397 456015 2431
rect 458005 2397 458039 2431
rect 460581 2397 460615 2431
rect 463157 2397 463191 2431
rect 465733 2397 465767 2431
rect 468309 2397 468343 2431
rect 470885 2397 470919 2431
rect 473461 2397 473495 2431
rect 476037 2397 476071 2431
rect 478613 2397 478647 2431
rect 481189 2397 481223 2431
rect 483765 2397 483799 2431
rect 486341 2397 486375 2431
rect 488917 2397 488951 2431
rect 491493 2397 491527 2431
rect 494069 2397 494103 2431
rect 496645 2397 496679 2431
rect 499221 2397 499255 2431
rect 501797 2397 501831 2431
rect 504373 2397 504407 2431
rect 506949 2397 506983 2431
rect 509525 2397 509559 2431
rect 512101 2397 512135 2431
rect 514677 2397 514711 2431
rect 1961 2329 1995 2363
rect 2513 2329 2547 2363
rect 7113 2329 7147 2363
rect 13645 2329 13679 2363
rect 14841 2329 14875 2363
rect 18797 2329 18831 2363
rect 19993 2329 20027 2363
rect 23213 2329 23247 2363
rect 25145 2329 25179 2363
rect 28365 2329 28399 2363
rect 30297 2329 30331 2363
rect 35449 2329 35483 2363
rect 38025 2329 38059 2363
rect 60013 2329 60047 2363
rect 76665 2329 76699 2363
rect 81817 2329 81851 2363
rect 84393 2329 84427 2363
rect 89545 2329 89579 2363
rect 91017 2329 91051 2363
rect 92121 2329 92155 2363
rect 97273 2329 97307 2363
rect 99849 2329 99883 2363
rect 105001 2329 105035 2363
rect 107577 2329 107611 2363
rect 112729 2329 112763 2363
rect 115305 2329 115339 2363
rect 120457 2329 120491 2363
rect 128185 2329 128219 2363
rect 138305 2329 138339 2363
rect 143457 2329 143491 2363
rect 146861 2329 146895 2363
rect 148609 2329 148643 2363
rect 164249 2329 164283 2363
rect 169401 2329 169435 2363
rect 174553 2329 174587 2363
rect 184857 2329 184891 2363
rect 190009 2329 190043 2363
rect 226073 2329 226107 2363
rect 350365 2329 350399 2363
rect 363245 2329 363279 2363
rect 458557 2329 458591 2363
rect 479165 2329 479199 2363
rect 4445 2261 4479 2295
rect 7021 2261 7055 2295
rect 12173 2261 12207 2295
rect 14749 2261 14783 2295
rect 17325 2261 17359 2295
rect 22477 2261 22511 2295
rect 23949 2261 23983 2295
rect 25053 2261 25087 2295
rect 27629 2261 27663 2295
rect 29101 2261 29135 2295
rect 30205 2261 30239 2295
rect 32781 2261 32815 2295
rect 35357 2261 35391 2295
rect 37933 2261 37967 2295
rect 40509 2261 40543 2295
rect 44557 2261 44591 2295
rect 48237 2261 48271 2295
rect 50813 2261 50847 2295
rect 53389 2261 53423 2295
rect 55965 2261 55999 2295
rect 58541 2261 58575 2295
rect 63693 2261 63727 2295
rect 64429 2261 64463 2295
rect 66269 2261 66303 2295
rect 71421 2261 71455 2295
rect 72157 2261 72191 2295
rect 75469 2261 75503 2295
rect 79149 2261 79183 2295
rect 79885 2261 79919 2295
rect 84301 2261 84335 2295
rect 86877 2261 86911 2295
rect 94605 2261 94639 2295
rect 99757 2261 99791 2295
rect 104909 2261 104943 2295
rect 106381 2261 106415 2295
rect 115213 2261 115247 2295
rect 120365 2261 120399 2295
rect 122941 2261 122975 2295
rect 125517 2261 125551 2295
rect 126253 2261 126287 2295
rect 128093 2261 128127 2295
rect 130853 2261 130887 2295
rect 133245 2261 133279 2295
rect 133981 2261 134015 2295
rect 136005 2261 136039 2295
rect 140973 2261 141007 2295
rect 146125 2261 146159 2295
rect 151277 2261 151311 2295
rect 152013 2261 152047 2295
rect 156429 2261 156463 2295
rect 157165 2261 157199 2295
rect 161581 2261 161615 2295
rect 162317 2261 162351 2295
rect 164157 2261 164191 2295
rect 166733 2261 166767 2295
rect 167469 2261 167503 2295
rect 169309 2261 169343 2295
rect 171885 2261 171919 2295
rect 172621 2261 172655 2295
rect 174461 2261 174495 2295
rect 177037 2261 177071 2295
rect 179613 2261 179647 2295
rect 182189 2261 182223 2295
rect 187341 2261 187375 2295
rect 189917 2261 189951 2295
rect 195069 2261 195103 2295
rect 197645 2261 197679 2295
rect 200221 2261 200255 2295
rect 202797 2261 202831 2295
rect 207949 2261 207983 2295
rect 213101 2261 213135 2295
rect 215677 2261 215711 2295
rect 218253 2261 218287 2295
rect 220829 2261 220863 2295
rect 223405 2261 223439 2295
rect 225981 2261 226015 2295
rect 228557 2261 228591 2295
rect 231133 2261 231167 2295
rect 233709 2261 233743 2295
rect 236285 2261 236319 2295
rect 238861 2261 238895 2295
rect 241437 2261 241471 2295
rect 244013 2261 244047 2295
rect 246589 2261 246623 2295
rect 249165 2261 249199 2295
rect 251741 2261 251775 2295
rect 254317 2261 254351 2295
rect 255053 2261 255087 2295
rect 256893 2261 256927 2295
rect 259469 2261 259503 2295
rect 262045 2261 262079 2295
rect 264621 2261 264655 2295
rect 267197 2261 267231 2295
rect 267933 2261 267967 2295
rect 269773 2261 269807 2295
rect 272349 2261 272383 2295
rect 274925 2261 274959 2295
rect 277501 2261 277535 2295
rect 278237 2261 278271 2295
rect 280077 2261 280111 2295
rect 282653 2261 282687 2295
rect 285229 2261 285263 2295
rect 287805 2261 287839 2295
rect 292957 2261 292991 2295
rect 298109 2261 298143 2295
rect 305837 2261 305871 2295
rect 310989 2261 311023 2295
rect 314301 2261 314335 2295
rect 316141 2261 316175 2295
rect 318717 2261 318751 2295
rect 319453 2261 319487 2295
rect 321293 2261 321327 2295
rect 323869 2261 323903 2295
rect 324605 2261 324639 2295
rect 326445 2261 326479 2295
rect 329021 2261 329055 2295
rect 329757 2261 329791 2295
rect 331597 2261 331631 2295
rect 332333 2261 332367 2295
rect 334173 2261 334207 2295
rect 336749 2261 336783 2295
rect 337485 2261 337519 2295
rect 339325 2261 339359 2295
rect 340061 2261 340095 2295
rect 341901 2261 341935 2295
rect 342637 2261 342671 2295
rect 344477 2261 344511 2295
rect 345213 2261 345247 2295
rect 347053 2261 347087 2295
rect 352205 2261 352239 2295
rect 354781 2261 354815 2295
rect 357357 2261 357391 2295
rect 358093 2261 358127 2295
rect 359933 2261 359967 2295
rect 362509 2261 362543 2295
rect 368397 2261 368431 2295
rect 370973 2261 371007 2295
rect 372813 2261 372847 2295
rect 377965 2261 377999 2295
rect 380541 2261 380575 2295
rect 381277 2261 381311 2295
rect 383117 2261 383151 2295
rect 383853 2261 383887 2295
rect 386429 2261 386463 2295
rect 389005 2261 389039 2295
rect 391581 2261 391615 2295
rect 401149 2261 401183 2295
rect 403725 2261 403759 2295
rect 406301 2261 406335 2295
rect 407037 2261 407071 2295
rect 408877 2261 408911 2295
rect 409613 2261 409647 2295
rect 411453 2261 411487 2295
rect 414029 2261 414063 2295
rect 416605 2261 416639 2295
rect 417341 2261 417375 2295
rect 419181 2261 419215 2295
rect 421757 2261 421791 2295
rect 422493 2261 422527 2295
rect 424333 2261 424367 2295
rect 426909 2261 426943 2295
rect 427645 2261 427679 2295
rect 429485 2261 429519 2295
rect 432061 2261 432095 2295
rect 432797 2261 432831 2295
rect 437213 2261 437247 2295
rect 440525 2261 440559 2295
rect 442365 2261 442399 2295
rect 443101 2261 443135 2295
rect 444941 2261 444975 2295
rect 447517 2261 447551 2295
rect 448253 2261 448287 2295
rect 450093 2261 450127 2295
rect 452669 2261 452703 2295
rect 455245 2261 455279 2295
rect 460397 2261 460431 2295
rect 462973 2261 463007 2295
rect 463709 2261 463743 2295
rect 465549 2261 465583 2295
rect 468125 2261 468159 2295
rect 468861 2261 468895 2295
rect 470701 2261 470735 2295
rect 471437 2261 471471 2295
rect 473277 2261 473311 2295
rect 473921 2261 473955 2295
rect 475853 2261 475887 2295
rect 478429 2261 478463 2295
rect 481005 2261 481039 2295
rect 483581 2261 483615 2295
rect 486157 2261 486191 2295
rect 488733 2261 488767 2295
rect 491309 2261 491343 2295
rect 493885 2261 493919 2295
rect 496461 2261 496495 2295
rect 499037 2261 499071 2295
rect 501613 2261 501647 2295
rect 504189 2261 504223 2295
rect 506765 2261 506799 2295
rect 509341 2261 509375 2295
rect 511917 2261 511951 2295
rect 514493 2261 514527 2295
<< metal1 >>
rect 92198 11908 92204 11960
rect 92256 11948 92262 11960
rect 199930 11948 199936 11960
rect 92256 11920 199936 11948
rect 92256 11908 92262 11920
rect 199930 11908 199936 11920
rect 199988 11908 199994 11960
rect 100662 11840 100668 11892
rect 100720 11880 100726 11892
rect 199194 11880 199200 11892
rect 100720 11852 199200 11880
rect 100720 11840 100726 11852
rect 199194 11840 199200 11852
rect 199252 11840 199258 11892
rect 175458 11772 175464 11824
rect 175516 11812 175522 11824
rect 195238 11812 195244 11824
rect 175516 11784 195244 11812
rect 175516 11772 175522 11784
rect 195238 11772 195244 11784
rect 195296 11772 195302 11824
rect 107562 11704 107568 11756
rect 107620 11744 107626 11756
rect 194962 11744 194968 11756
rect 107620 11716 194968 11744
rect 107620 11704 107626 11716
rect 194962 11704 194968 11716
rect 195020 11704 195026 11756
rect 99926 11636 99932 11688
rect 99984 11676 99990 11688
rect 199378 11676 199384 11688
rect 99984 11648 199384 11676
rect 99984 11636 99990 11648
rect 199378 11636 199384 11648
rect 199436 11636 199442 11688
rect 184382 11568 184388 11620
rect 184440 11608 184446 11620
rect 195606 11608 195612 11620
rect 184440 11580 195612 11608
rect 184440 11568 184446 11580
rect 195606 11568 195612 11580
rect 195664 11568 195670 11620
rect 157886 11500 157892 11552
rect 157944 11540 157950 11552
rect 199838 11540 199844 11552
rect 157944 11512 199844 11540
rect 157944 11500 157950 11512
rect 199838 11500 199844 11512
rect 199896 11500 199902 11552
rect 97442 11432 97448 11484
rect 97500 11472 97506 11484
rect 195514 11472 195520 11484
rect 97500 11444 195520 11472
rect 97500 11432 97506 11444
rect 195514 11432 195520 11444
rect 195572 11432 195578 11484
rect 195882 11432 195888 11484
rect 195940 11472 195946 11484
rect 199286 11472 199292 11484
rect 195940 11444 199292 11472
rect 195940 11432 195946 11444
rect 199286 11432 199292 11444
rect 199344 11432 199350 11484
rect 195054 11364 195060 11416
rect 195112 11404 195118 11416
rect 200062 11404 200118 12000
rect 200390 11840 200396 11892
rect 200448 11880 200454 11892
rect 200606 11880 200662 12000
rect 200448 11852 200662 11880
rect 200448 11840 200454 11852
rect 195112 11376 200118 11404
rect 195112 11364 195118 11376
rect 186682 11296 186688 11348
rect 186740 11336 186746 11348
rect 199378 11336 199384 11348
rect 186740 11308 199384 11336
rect 186740 11296 186746 11308
rect 199378 11296 199384 11308
rect 199436 11296 199442 11348
rect 92842 11228 92848 11280
rect 92900 11268 92906 11280
rect 92900 11240 198596 11268
rect 92900 11228 92906 11240
rect 123110 11160 123116 11212
rect 123168 11200 123174 11212
rect 184198 11200 184204 11212
rect 123168 11172 184204 11200
rect 123168 11160 123174 11172
rect 184198 11160 184204 11172
rect 184256 11160 184262 11212
rect 195238 11160 195244 11212
rect 195296 11200 195302 11212
rect 198458 11200 198464 11212
rect 195296 11172 198464 11200
rect 195296 11160 195302 11172
rect 198458 11160 198464 11172
rect 198516 11160 198522 11212
rect 198568 11200 198596 11240
rect 199930 11200 199936 11212
rect 198568 11172 199936 11200
rect 199930 11160 199936 11172
rect 199988 11160 199994 11212
rect 200062 11200 200118 11376
rect 200606 11200 200662 11852
rect 200850 11228 200856 11280
rect 200908 11268 200914 11280
rect 201150 11268 201206 12000
rect 200908 11240 201206 11268
rect 200908 11228 200914 11240
rect 201150 11200 201206 11240
rect 201310 11228 201316 11280
rect 201368 11268 201374 11280
rect 201694 11268 201750 12000
rect 201368 11240 201750 11268
rect 201368 11228 201374 11240
rect 201694 11200 201750 11240
rect 201954 11228 201960 11280
rect 202012 11268 202018 11280
rect 202238 11268 202294 12000
rect 202012 11240 202294 11268
rect 202012 11228 202018 11240
rect 202238 11200 202294 11240
rect 202506 11228 202512 11280
rect 202564 11268 202570 11280
rect 202782 11268 202838 12000
rect 202564 11240 202838 11268
rect 202564 11228 202570 11240
rect 202782 11200 202838 11240
rect 202966 11228 202972 11280
rect 203024 11268 203030 11280
rect 203326 11268 203382 12000
rect 203024 11240 203382 11268
rect 203024 11228 203030 11240
rect 203326 11200 203382 11240
rect 203426 11228 203432 11280
rect 203484 11268 203490 11280
rect 203870 11268 203926 12000
rect 204414 11268 204470 12000
rect 204958 11268 205014 12000
rect 203484 11240 203926 11268
rect 203484 11228 203490 11240
rect 203870 11200 203926 11240
rect 204088 11240 204470 11268
rect 203978 11160 203984 11212
rect 204036 11200 204042 11212
rect 204088 11200 204116 11240
rect 204414 11200 204470 11240
rect 204640 11240 205014 11268
rect 204036 11172 204116 11200
rect 204036 11160 204042 11172
rect 204530 11160 204536 11212
rect 204588 11200 204594 11212
rect 204640 11200 204668 11240
rect 204958 11200 205014 11240
rect 205082 11228 205088 11280
rect 205140 11268 205146 11280
rect 205502 11268 205558 12000
rect 205634 11568 205640 11620
rect 205692 11608 205698 11620
rect 206046 11608 206102 12000
rect 205692 11580 206102 11608
rect 205692 11568 205698 11580
rect 205140 11240 205558 11268
rect 205140 11228 205146 11240
rect 205502 11200 205558 11240
rect 206046 11200 206102 11580
rect 206186 11228 206192 11280
rect 206244 11268 206250 11280
rect 206590 11268 206646 12000
rect 207134 11268 207190 12000
rect 206244 11240 206646 11268
rect 206244 11228 206250 11240
rect 206590 11200 206646 11240
rect 207032 11240 207190 11268
rect 204588 11172 204668 11200
rect 204588 11160 204594 11172
rect 98454 11092 98460 11144
rect 98512 11132 98518 11144
rect 195330 11132 195336 11144
rect 98512 11104 195336 11132
rect 98512 11092 98518 11104
rect 195330 11092 195336 11104
rect 195388 11092 195394 11144
rect 199838 11092 199844 11144
rect 199896 11132 199902 11144
rect 207032 11132 207060 11240
rect 207134 11200 207190 11240
rect 207474 11228 207480 11280
rect 207532 11268 207538 11280
rect 207678 11268 207734 12000
rect 207532 11240 207734 11268
rect 207532 11228 207538 11240
rect 207678 11200 207734 11240
rect 208118 11228 208124 11280
rect 208176 11268 208182 11280
rect 208222 11268 208278 12000
rect 208176 11240 208278 11268
rect 208176 11228 208182 11240
rect 208222 11200 208278 11240
rect 208578 11228 208584 11280
rect 208636 11268 208642 11280
rect 208766 11268 208822 12000
rect 209310 11268 209366 12000
rect 208636 11240 208822 11268
rect 208636 11228 208642 11240
rect 208766 11200 208822 11240
rect 209056 11240 209366 11268
rect 209056 11200 209084 11240
rect 209310 11200 209366 11240
rect 209854 11268 209910 12000
rect 209958 11268 209964 11280
rect 209854 11240 209964 11268
rect 209854 11200 209910 11240
rect 209958 11228 209964 11240
rect 210016 11228 210022 11280
rect 210398 11268 210454 12000
rect 210160 11240 210454 11268
rect 208872 11172 209084 11200
rect 199896 11104 205772 11132
rect 207032 11104 207152 11132
rect 199896 11092 199902 11104
rect 104066 11024 104072 11076
rect 104124 11064 104130 11076
rect 195238 11064 195244 11076
rect 104124 11036 195244 11064
rect 104124 11024 104130 11036
rect 195238 11024 195244 11036
rect 195296 11024 195302 11076
rect 195606 11024 195612 11076
rect 195664 11064 195670 11076
rect 195664 11036 199056 11064
rect 195664 11024 195670 11036
rect 180766 10968 195468 10996
rect 97258 10888 97264 10940
rect 97316 10928 97322 10940
rect 180766 10928 180794 10968
rect 97316 10900 180794 10928
rect 195440 10928 195468 10968
rect 195514 10956 195520 11008
rect 195572 10996 195578 11008
rect 198550 10996 198556 11008
rect 195572 10968 198556 10996
rect 195572 10956 195578 10968
rect 198550 10956 198556 10968
rect 198608 10956 198614 11008
rect 198642 10928 198648 10940
rect 195440 10900 198648 10928
rect 97316 10888 97322 10900
rect 198642 10888 198648 10900
rect 198700 10888 198706 10940
rect 199028 10928 199056 11036
rect 199194 11024 199200 11076
rect 199252 11064 199258 11076
rect 205450 11064 205456 11076
rect 199252 11036 205456 11064
rect 199252 11024 199258 11036
rect 205450 11024 205456 11036
rect 205508 11024 205514 11076
rect 205542 11024 205548 11076
rect 205600 11064 205606 11076
rect 205634 11064 205640 11076
rect 205600 11036 205640 11064
rect 205600 11024 205606 11036
rect 205634 11024 205640 11036
rect 205692 11024 205698 11076
rect 205744 11064 205772 11104
rect 207014 11064 207020 11076
rect 205744 11036 207020 11064
rect 207014 11024 207020 11036
rect 207072 11024 207078 11076
rect 207124 11064 207152 11104
rect 207290 11092 207296 11144
rect 207348 11132 207354 11144
rect 208872 11132 208900 11172
rect 210050 11160 210056 11212
rect 210108 11200 210114 11212
rect 210160 11200 210188 11240
rect 210398 11200 210454 11240
rect 210694 11228 210700 11280
rect 210752 11268 210758 11280
rect 210942 11268 210998 12000
rect 210752 11240 210998 11268
rect 210752 11228 210758 11240
rect 210942 11200 210998 11240
rect 211154 11228 211160 11280
rect 211212 11268 211218 11280
rect 211486 11268 211542 12000
rect 211212 11240 211542 11268
rect 211212 11228 211218 11240
rect 211486 11200 211542 11240
rect 211798 11228 211804 11280
rect 211856 11268 211862 11280
rect 212030 11268 212086 12000
rect 211856 11240 212086 11268
rect 211856 11228 211862 11240
rect 212030 11200 212086 11240
rect 212574 11268 212630 12000
rect 212902 11364 212908 11416
rect 212960 11404 212966 11416
rect 213118 11404 213174 12000
rect 212960 11376 213174 11404
rect 212960 11364 212966 11376
rect 212718 11268 212724 11280
rect 212574 11240 212724 11268
rect 212574 11200 212630 11240
rect 212718 11228 212724 11240
rect 212776 11228 212782 11280
rect 213118 11200 213174 11376
rect 213662 11268 213718 12000
rect 213822 11268 213828 11280
rect 213662 11240 213828 11268
rect 213662 11200 213718 11240
rect 213822 11228 213828 11240
rect 213880 11228 213886 11280
rect 213914 11228 213920 11280
rect 213972 11268 213978 11280
rect 214206 11268 214262 12000
rect 214374 11432 214380 11484
rect 214432 11472 214438 11484
rect 214750 11472 214806 12000
rect 214432 11444 214806 11472
rect 214432 11432 214438 11444
rect 213972 11240 214262 11268
rect 213972 11228 213978 11240
rect 214206 11200 214262 11240
rect 214750 11200 214806 11444
rect 215294 11268 215350 12000
rect 215386 11268 215392 11280
rect 215294 11240 215392 11268
rect 215294 11200 215350 11240
rect 215386 11228 215392 11240
rect 215444 11228 215450 11280
rect 215570 11228 215576 11280
rect 215628 11268 215634 11280
rect 215838 11268 215894 12000
rect 216382 11268 216438 12000
rect 215628 11240 215894 11268
rect 215628 11228 215634 11240
rect 215838 11200 215894 11240
rect 215956 11240 216438 11268
rect 210108 11172 210188 11200
rect 210108 11160 210114 11172
rect 213638 11132 213644 11144
rect 207348 11104 208900 11132
rect 208964 11104 213644 11132
rect 207348 11092 207354 11104
rect 207124 11036 207176 11064
rect 199930 10956 199936 11008
rect 199988 10996 199994 11008
rect 201310 10996 201316 11008
rect 199988 10968 201316 10996
rect 199988 10956 199994 10968
rect 201310 10956 201316 10968
rect 201368 10956 201374 11008
rect 201402 10956 201408 11008
rect 201460 10996 201466 11008
rect 207148 10996 207176 11036
rect 207382 11024 207388 11076
rect 207440 11064 207446 11076
rect 208964 11064 208992 11104
rect 213638 11092 213644 11104
rect 213696 11092 213702 11144
rect 214006 11092 214012 11144
rect 214064 11132 214070 11144
rect 215956 11132 215984 11240
rect 216382 11200 216438 11240
rect 216926 11268 216982 12000
rect 217042 11268 217048 11280
rect 216926 11240 217048 11268
rect 216926 11200 216982 11240
rect 217042 11228 217048 11240
rect 217100 11228 217106 11280
rect 217226 11228 217232 11280
rect 217284 11268 217290 11280
rect 217470 11268 217526 12000
rect 217284 11240 217526 11268
rect 217284 11228 217290 11240
rect 217470 11200 217526 11240
rect 217594 11228 217600 11280
rect 217652 11268 217658 11280
rect 218014 11268 218070 12000
rect 217652 11240 218070 11268
rect 217652 11228 217658 11240
rect 218014 11200 218070 11240
rect 218330 11228 218336 11280
rect 218388 11268 218394 11280
rect 218558 11268 218614 12000
rect 218388 11240 218614 11268
rect 218388 11228 218394 11240
rect 218558 11200 218614 11240
rect 219102 11336 219158 12000
rect 219250 11336 219256 11348
rect 219102 11308 219256 11336
rect 219102 11200 219158 11308
rect 219250 11296 219256 11308
rect 219308 11296 219314 11348
rect 219434 11228 219440 11280
rect 219492 11268 219498 11280
rect 219646 11268 219702 12000
rect 220190 11268 220246 12000
rect 219492 11240 219702 11268
rect 219492 11228 219498 11240
rect 219646 11200 219702 11240
rect 219912 11240 220246 11268
rect 219912 11212 219940 11240
rect 219894 11160 219900 11212
rect 219952 11160 219958 11212
rect 220190 11200 220246 11240
rect 220354 11228 220360 11280
rect 220412 11268 220418 11280
rect 220734 11268 220790 12000
rect 220412 11240 220790 11268
rect 220412 11228 220418 11240
rect 220734 11200 220790 11240
rect 220906 11228 220912 11280
rect 220964 11268 220970 11280
rect 221278 11268 221334 12000
rect 220964 11240 221334 11268
rect 220964 11228 220970 11240
rect 221278 11200 221334 11240
rect 221642 11228 221648 11280
rect 221700 11268 221706 11280
rect 221822 11268 221878 12000
rect 221700 11240 221878 11268
rect 221700 11228 221706 11240
rect 221822 11200 221878 11240
rect 222194 11228 222200 11280
rect 222252 11268 222258 11280
rect 222366 11268 222422 12000
rect 222252 11240 222422 11268
rect 222252 11228 222258 11240
rect 222366 11200 222422 11240
rect 222470 11228 222476 11280
rect 222528 11268 222534 11280
rect 222910 11268 222966 12000
rect 222528 11240 222966 11268
rect 222528 11228 222534 11240
rect 222910 11200 222966 11240
rect 223206 11228 223212 11280
rect 223264 11268 223270 11280
rect 223454 11268 223510 12000
rect 223264 11240 223510 11268
rect 223264 11228 223270 11240
rect 223454 11200 223510 11240
rect 223758 11228 223764 11280
rect 223816 11268 223822 11280
rect 223998 11268 224054 12000
rect 224542 11336 224598 12000
rect 223816 11240 224054 11268
rect 223816 11228 223822 11240
rect 223998 11200 224054 11240
rect 224236 11308 224598 11336
rect 214064 11104 215984 11132
rect 214064 11092 214070 11104
rect 216766 11092 216772 11144
rect 216824 11132 216830 11144
rect 224236 11132 224264 11308
rect 224542 11200 224598 11308
rect 224954 11228 224960 11280
rect 225012 11268 225018 11280
rect 225086 11268 225142 12000
rect 225012 11240 225142 11268
rect 225012 11228 225018 11240
rect 225086 11200 225142 11240
rect 225414 11228 225420 11280
rect 225472 11268 225478 11280
rect 225630 11268 225686 12000
rect 225472 11240 225686 11268
rect 225472 11228 225478 11240
rect 225630 11200 225686 11240
rect 225782 11228 225788 11280
rect 225840 11268 225846 11280
rect 226174 11268 226230 12000
rect 225840 11240 226230 11268
rect 225840 11228 225846 11240
rect 226174 11200 226230 11240
rect 226426 11228 226432 11280
rect 226484 11268 226490 11280
rect 226718 11268 226774 12000
rect 226484 11240 226774 11268
rect 226484 11228 226490 11240
rect 226718 11200 226774 11240
rect 226978 11228 226984 11280
rect 227036 11268 227042 11280
rect 227262 11268 227318 12000
rect 227036 11240 227318 11268
rect 227036 11228 227042 11240
rect 227262 11200 227318 11240
rect 227346 11228 227352 11280
rect 227404 11268 227410 11280
rect 227806 11268 227862 12000
rect 227404 11240 227862 11268
rect 227404 11228 227410 11240
rect 227806 11200 227862 11240
rect 228082 11228 228088 11280
rect 228140 11268 228146 11280
rect 228350 11268 228406 12000
rect 228140 11240 228406 11268
rect 228140 11228 228146 11240
rect 228350 11200 228406 11240
rect 228450 11228 228456 11280
rect 228508 11268 228514 11280
rect 228894 11268 228950 12000
rect 228508 11240 228950 11268
rect 228508 11228 228514 11240
rect 228894 11200 228950 11240
rect 229186 11228 229192 11280
rect 229244 11268 229250 11280
rect 229438 11268 229494 12000
rect 229244 11240 229494 11268
rect 229244 11228 229250 11240
rect 229438 11200 229494 11240
rect 229830 11228 229836 11280
rect 229888 11268 229894 11280
rect 229982 11268 230038 12000
rect 229888 11240 230038 11268
rect 229888 11228 229894 11240
rect 229982 11200 230038 11240
rect 230382 11228 230388 11280
rect 230440 11268 230446 11280
rect 230526 11268 230582 12000
rect 230440 11240 230582 11268
rect 230440 11228 230446 11240
rect 230526 11200 230582 11240
rect 230842 11228 230848 11280
rect 230900 11268 230906 11280
rect 231070 11268 231126 12000
rect 230900 11240 231126 11268
rect 230900 11228 230906 11240
rect 231070 11200 231126 11240
rect 231394 11228 231400 11280
rect 231452 11268 231458 11280
rect 231614 11268 231670 12000
rect 231452 11240 231670 11268
rect 231452 11228 231458 11240
rect 231614 11200 231670 11240
rect 231854 11228 231860 11280
rect 231912 11268 231918 11280
rect 232158 11268 232214 12000
rect 231912 11240 232214 11268
rect 231912 11228 231918 11240
rect 232158 11200 232214 11240
rect 232314 11228 232320 11280
rect 232372 11268 232378 11280
rect 232702 11268 232758 12000
rect 232372 11240 232758 11268
rect 232372 11228 232378 11240
rect 232702 11200 232758 11240
rect 233246 11268 233302 12000
rect 233418 11268 233424 11280
rect 233246 11240 233424 11268
rect 233246 11200 233302 11240
rect 233418 11228 233424 11240
rect 233476 11228 233482 11280
rect 233602 11228 233608 11280
rect 233660 11268 233666 11280
rect 233790 11268 233846 12000
rect 233660 11240 233846 11268
rect 233660 11228 233666 11240
rect 233790 11200 233846 11240
rect 233878 11228 233884 11280
rect 233936 11268 233942 11280
rect 234334 11268 234390 12000
rect 233936 11240 234390 11268
rect 233936 11228 233942 11240
rect 234334 11200 234390 11240
rect 234706 11228 234712 11280
rect 234764 11268 234770 11280
rect 234878 11268 234934 12000
rect 234764 11240 234934 11268
rect 234764 11228 234770 11240
rect 234878 11200 234934 11240
rect 234982 11228 234988 11280
rect 235040 11268 235046 11280
rect 235422 11268 235478 12000
rect 235040 11240 235478 11268
rect 235040 11228 235046 11240
rect 235422 11200 235478 11240
rect 235718 11228 235724 11280
rect 235776 11268 235782 11280
rect 235966 11268 236022 12000
rect 235776 11240 236022 11268
rect 235776 11228 235782 11240
rect 235966 11200 236022 11240
rect 236270 11228 236276 11280
rect 236328 11268 236334 11280
rect 236510 11268 236566 12000
rect 236328 11240 236566 11268
rect 236328 11228 236334 11240
rect 236510 11200 236566 11240
rect 236914 11228 236920 11280
rect 236972 11268 236978 11280
rect 237054 11268 237110 12000
rect 236972 11240 237110 11268
rect 236972 11228 236978 11240
rect 237054 11200 237110 11240
rect 237374 11228 237380 11280
rect 237432 11268 237438 11280
rect 237598 11268 237654 12000
rect 237432 11240 237654 11268
rect 237432 11228 237438 11240
rect 237598 11200 237654 11240
rect 237926 11228 237932 11280
rect 237984 11268 237990 11280
rect 238142 11268 238198 12000
rect 237984 11240 238198 11268
rect 237984 11228 237990 11240
rect 238142 11200 238198 11240
rect 238294 11228 238300 11280
rect 238352 11268 238358 11280
rect 238686 11268 238742 12000
rect 238352 11240 238742 11268
rect 238352 11228 238358 11240
rect 238686 11200 238742 11240
rect 238938 11228 238944 11280
rect 238996 11268 239002 11280
rect 239230 11268 239286 12000
rect 238996 11240 239286 11268
rect 238996 11228 239002 11240
rect 239230 11200 239286 11240
rect 239490 11228 239496 11280
rect 239548 11268 239554 11280
rect 239774 11268 239830 12000
rect 239548 11240 239830 11268
rect 239548 11228 239554 11240
rect 239774 11200 239830 11240
rect 240134 11228 240140 11280
rect 240192 11268 240198 11280
rect 240318 11268 240374 12000
rect 240192 11240 240374 11268
rect 240192 11228 240198 11240
rect 240318 11200 240374 11240
rect 240410 11228 240416 11280
rect 240468 11268 240474 11280
rect 240862 11268 240918 12000
rect 240468 11240 240918 11268
rect 240468 11228 240474 11240
rect 240862 11200 240918 11240
rect 241146 11228 241152 11280
rect 241204 11268 241210 11280
rect 241406 11268 241462 12000
rect 241204 11240 241462 11268
rect 241204 11228 241210 11240
rect 241406 11200 241462 11240
rect 241606 11228 241612 11280
rect 241664 11268 241670 11280
rect 241950 11268 242006 12000
rect 241664 11240 242006 11268
rect 241664 11228 241670 11240
rect 241950 11200 242006 11240
rect 242494 11268 242550 12000
rect 242494 11200 242572 11268
rect 242894 11228 242900 11280
rect 242952 11268 242958 11280
rect 243038 11268 243094 12000
rect 242952 11240 243094 11268
rect 242952 11228 242958 11240
rect 243038 11200 243094 11240
rect 243354 11228 243360 11280
rect 243412 11268 243418 11280
rect 243582 11268 243638 12000
rect 244126 11268 244182 12000
rect 243412 11240 243638 11268
rect 243412 11228 243418 11240
rect 243582 11200 243638 11240
rect 242498 11172 242572 11200
rect 244108 11172 244182 11268
rect 244458 11228 244464 11280
rect 244516 11268 244522 11280
rect 244670 11268 244726 12000
rect 244516 11240 244726 11268
rect 244516 11228 244522 11240
rect 244670 11200 244726 11240
rect 245010 11228 245016 11280
rect 245068 11268 245074 11280
rect 245214 11268 245270 12000
rect 245068 11240 245270 11268
rect 245068 11228 245074 11240
rect 245214 11200 245270 11240
rect 245378 11228 245384 11280
rect 245436 11268 245442 11280
rect 245758 11268 245814 12000
rect 245436 11240 245814 11268
rect 245436 11228 245442 11240
rect 245758 11200 245814 11240
rect 246114 11228 246120 11280
rect 246172 11268 246178 11280
rect 246302 11268 246358 12000
rect 246172 11240 246358 11268
rect 246172 11228 246178 11240
rect 246302 11200 246358 11240
rect 246666 11228 246672 11280
rect 246724 11268 246730 11280
rect 246846 11268 246902 12000
rect 246724 11240 246902 11268
rect 246724 11228 246730 11240
rect 246846 11200 246902 11240
rect 246942 11228 246948 11280
rect 247000 11268 247006 11280
rect 247390 11268 247446 12000
rect 247000 11240 247446 11268
rect 247000 11228 247006 11240
rect 247390 11200 247446 11240
rect 247678 11228 247684 11280
rect 247736 11268 247742 11280
rect 247934 11268 247990 12000
rect 247736 11240 247990 11268
rect 247736 11228 247742 11240
rect 247934 11200 247990 11240
rect 248478 11268 248534 12000
rect 248478 11200 248552 11268
rect 248598 11228 248604 11280
rect 248656 11268 248662 11280
rect 249022 11268 249078 12000
rect 248656 11240 249078 11268
rect 248656 11228 248662 11240
rect 249022 11200 249078 11240
rect 249334 11228 249340 11280
rect 249392 11268 249398 11280
rect 249566 11268 249622 12000
rect 249392 11240 249622 11268
rect 249392 11228 249398 11240
rect 249566 11200 249622 11240
rect 249978 11228 249984 11280
rect 250036 11268 250042 11280
rect 250110 11268 250166 12000
rect 250036 11240 250166 11268
rect 250036 11228 250042 11240
rect 250110 11200 250166 11240
rect 250254 11228 250260 11280
rect 250312 11268 250318 11280
rect 250654 11268 250710 12000
rect 250312 11240 250710 11268
rect 250312 11228 250318 11240
rect 250654 11200 250710 11240
rect 251198 11268 251254 12000
rect 251198 11240 251312 11268
rect 251198 11200 251254 11240
rect 216824 11104 224264 11132
rect 216824 11092 216830 11104
rect 224770 11092 224776 11144
rect 224828 11132 224834 11144
rect 226886 11132 226892 11144
rect 224828 11104 226892 11132
rect 224828 11092 224834 11104
rect 226886 11092 226892 11104
rect 226944 11092 226950 11144
rect 242498 11132 242526 11172
rect 226996 11104 242526 11132
rect 207440 11036 208992 11064
rect 207440 11024 207446 11036
rect 211062 11024 211068 11076
rect 211120 11064 211126 11076
rect 226996 11064 227024 11104
rect 211120 11036 227024 11064
rect 211120 11024 211126 11036
rect 229278 11024 229284 11076
rect 229336 11064 229342 11076
rect 236638 11064 236644 11076
rect 229336 11036 236644 11064
rect 229336 11024 229342 11036
rect 236638 11024 236644 11036
rect 236696 11024 236702 11076
rect 239398 11024 239404 11076
rect 239456 11064 239462 11076
rect 244154 11064 244182 11172
rect 248524 11144 248552 11200
rect 251284 11144 251312 11240
rect 251542 11228 251548 11280
rect 251600 11268 251606 11280
rect 251742 11268 251798 12000
rect 251600 11240 251798 11268
rect 251600 11228 251606 11240
rect 251742 11200 251798 11240
rect 251910 11228 251916 11280
rect 251968 11268 251974 11280
rect 252286 11268 252342 12000
rect 251968 11240 252342 11268
rect 251968 11228 251974 11240
rect 252286 11200 252342 11240
rect 252738 11228 252744 11280
rect 252796 11268 252802 11280
rect 252830 11268 252886 12000
rect 252796 11240 252886 11268
rect 252796 11228 252802 11240
rect 252830 11200 252886 11240
rect 253106 11228 253112 11280
rect 253164 11268 253170 11280
rect 253374 11268 253430 12000
rect 253164 11240 253430 11268
rect 253164 11228 253170 11240
rect 253374 11200 253430 11240
rect 253918 11268 253974 12000
rect 254210 11296 254216 11348
rect 254268 11336 254274 11348
rect 254462 11336 254518 12000
rect 254268 11308 254518 11336
rect 254268 11296 254274 11308
rect 254026 11268 254032 11280
rect 253918 11240 254032 11268
rect 253918 11200 253974 11240
rect 254026 11228 254032 11240
rect 254084 11228 254090 11280
rect 254462 11200 254518 11308
rect 255006 11268 255062 12000
rect 255006 11200 255084 11268
rect 255314 11228 255320 11280
rect 255372 11268 255378 11280
rect 255550 11268 255606 12000
rect 255372 11240 255606 11268
rect 255372 11228 255378 11240
rect 255550 11200 255606 11240
rect 255866 11228 255872 11280
rect 255924 11268 255930 11280
rect 256094 11268 256150 12000
rect 255924 11240 256150 11268
rect 255924 11228 255930 11240
rect 256094 11200 256150 11240
rect 256418 11228 256424 11280
rect 256476 11268 256482 11280
rect 256638 11268 256694 12000
rect 257182 11268 257238 12000
rect 277118 11636 277124 11688
rect 277176 11676 277182 11688
rect 359734 11676 359740 11688
rect 277176 11648 359740 11676
rect 277176 11636 277182 11648
rect 359734 11636 359740 11648
rect 359792 11636 359798 11688
rect 359918 11608 359924 11620
rect 256476 11240 256694 11268
rect 256476 11228 256482 11240
rect 256638 11200 256694 11240
rect 256804 11240 257238 11268
rect 255010 11172 255084 11200
rect 248506 11092 248512 11144
rect 248564 11092 248570 11144
rect 251266 11092 251272 11144
rect 251324 11092 251330 11144
rect 239456 11036 244182 11064
rect 239456 11024 239462 11036
rect 255010 11008 255038 11172
rect 255682 11092 255688 11144
rect 255740 11132 255746 11144
rect 256804 11132 256832 11240
rect 257182 11200 257238 11240
rect 258460 11580 359924 11608
rect 255740 11104 256832 11132
rect 255740 11092 255746 11104
rect 255222 11024 255228 11076
rect 255280 11064 255286 11076
rect 258460 11064 258488 11580
rect 359918 11568 359924 11580
rect 359976 11568 359982 11620
rect 258718 11500 258724 11552
rect 258776 11540 258782 11552
rect 354398 11540 354404 11552
rect 258776 11512 354404 11540
rect 258776 11500 258782 11512
rect 354398 11500 354404 11512
rect 354456 11500 354462 11552
rect 258626 11432 258632 11484
rect 258684 11472 258690 11484
rect 358630 11472 358636 11484
rect 258684 11444 358636 11472
rect 258684 11432 258690 11444
rect 358630 11432 358636 11444
rect 358688 11432 358694 11484
rect 258534 11364 258540 11416
rect 258592 11404 258598 11416
rect 311250 11404 311256 11416
rect 258592 11376 311256 11404
rect 258592 11364 258598 11376
rect 311250 11364 311256 11376
rect 311308 11364 311314 11416
rect 346762 11336 346768 11348
rect 255280 11036 258488 11064
rect 258552 11308 346768 11336
rect 255280 11024 255286 11036
rect 201460 10968 207176 10996
rect 201460 10956 201466 10968
rect 207290 10956 207296 11008
rect 207348 10996 207354 11008
rect 212074 10996 212080 11008
rect 207348 10968 212080 10996
rect 207348 10956 207354 10968
rect 212074 10956 212080 10968
rect 212132 10956 212138 11008
rect 212166 10956 212172 11008
rect 212224 10996 212230 11008
rect 224770 10996 224776 11008
rect 212224 10968 224776 10996
rect 212224 10956 212230 10968
rect 224770 10956 224776 10968
rect 224828 10956 224834 11008
rect 229646 10956 229652 11008
rect 229704 10996 229710 11008
rect 239214 10996 239220 11008
rect 229704 10968 239220 10996
rect 229704 10956 229710 10968
rect 239214 10956 239220 10968
rect 239272 10956 239278 11008
rect 254946 10956 254952 11008
rect 255004 10968 255038 11008
rect 258552 10996 258580 11308
rect 346762 11296 346768 11308
rect 346820 11296 346826 11348
rect 347590 11296 347596 11348
rect 347648 11336 347654 11348
rect 355778 11336 355784 11348
rect 347648 11308 355784 11336
rect 347648 11296 347654 11308
rect 355778 11296 355784 11308
rect 355836 11296 355842 11348
rect 360066 11268 360122 12000
rect 357406 11240 360122 11268
rect 336274 11200 336280 11212
rect 258460 10968 258580 10996
rect 258736 11172 336280 11200
rect 255004 10956 255010 10968
rect 199028 10900 201356 10928
rect 102870 10820 102876 10872
rect 102928 10860 102934 10872
rect 102928 10832 195284 10860
rect 102928 10820 102934 10832
rect 96062 10752 96068 10804
rect 96120 10792 96126 10804
rect 195146 10792 195152 10804
rect 96120 10764 195152 10792
rect 96120 10752 96126 10764
rect 195146 10752 195152 10764
rect 195204 10752 195210 10804
rect 195256 10792 195284 10832
rect 195330 10820 195336 10872
rect 195388 10860 195394 10872
rect 201218 10860 201224 10872
rect 195388 10832 201224 10860
rect 195388 10820 195394 10832
rect 201218 10820 201224 10832
rect 201276 10820 201282 10872
rect 201328 10860 201356 10900
rect 201494 10888 201500 10940
rect 201552 10928 201558 10940
rect 216766 10928 216772 10940
rect 201552 10900 216772 10928
rect 201552 10888 201558 10900
rect 216766 10888 216772 10900
rect 216824 10888 216830 10940
rect 235718 10928 235724 10940
rect 229112 10900 235724 10928
rect 220170 10860 220176 10872
rect 201328 10832 220176 10860
rect 220170 10820 220176 10832
rect 220228 10820 220234 10872
rect 221366 10820 221372 10872
rect 221424 10860 221430 10872
rect 221424 10832 225184 10860
rect 221424 10820 221430 10832
rect 206922 10792 206928 10804
rect 195256 10764 206928 10792
rect 206922 10752 206928 10764
rect 206980 10752 206986 10804
rect 207014 10752 207020 10804
rect 207072 10792 207078 10804
rect 207072 10764 212304 10792
rect 207072 10752 207078 10764
rect 101950 10684 101956 10736
rect 102008 10724 102014 10736
rect 205634 10724 205640 10736
rect 102008 10696 205640 10724
rect 102008 10684 102014 10696
rect 205634 10684 205640 10696
rect 205692 10684 205698 10736
rect 205726 10684 205732 10736
rect 205784 10724 205790 10736
rect 212166 10724 212172 10736
rect 205784 10696 212172 10724
rect 205784 10684 205790 10696
rect 212166 10684 212172 10696
rect 212224 10684 212230 10736
rect 212276 10724 212304 10764
rect 212350 10752 212356 10804
rect 212408 10792 212414 10804
rect 225046 10792 225052 10804
rect 212408 10764 225052 10792
rect 212408 10752 212414 10764
rect 225046 10752 225052 10764
rect 225104 10752 225110 10804
rect 225156 10792 225184 10832
rect 226886 10820 226892 10872
rect 226944 10860 226950 10872
rect 229112 10860 229140 10900
rect 235718 10888 235724 10900
rect 235776 10888 235782 10940
rect 236638 10888 236644 10940
rect 236696 10928 236702 10940
rect 248690 10928 248696 10940
rect 236696 10900 248696 10928
rect 236696 10888 236702 10900
rect 248690 10888 248696 10900
rect 248748 10888 248754 10940
rect 249058 10888 249064 10940
rect 249116 10928 249122 10940
rect 258460 10928 258488 10968
rect 249116 10900 258488 10928
rect 249116 10888 249122 10900
rect 226944 10832 229140 10860
rect 226944 10820 226950 10832
rect 229738 10820 229744 10872
rect 229796 10860 229802 10872
rect 239398 10860 239404 10872
rect 229796 10832 239404 10860
rect 229796 10820 229802 10832
rect 239398 10820 239404 10832
rect 239456 10820 239462 10872
rect 258534 10860 258540 10872
rect 241486 10832 258540 10860
rect 238846 10792 238852 10804
rect 225156 10764 238852 10792
rect 238846 10752 238852 10764
rect 238904 10752 238910 10804
rect 219434 10724 219440 10736
rect 212276 10696 219440 10724
rect 219434 10684 219440 10696
rect 219492 10684 219498 10736
rect 220078 10684 220084 10736
rect 220136 10724 220142 10736
rect 241486 10724 241514 10832
rect 258534 10820 258540 10832
rect 258592 10820 258598 10872
rect 248690 10752 248696 10804
rect 248748 10792 248754 10804
rect 258736 10792 258764 11172
rect 336274 11160 336280 11172
rect 336332 11160 336338 11212
rect 342714 11160 342720 11212
rect 342772 11200 342778 11212
rect 355410 11200 355416 11212
rect 342772 11172 355416 11200
rect 342772 11160 342778 11172
rect 355410 11160 355416 11172
rect 355468 11160 355474 11212
rect 357406 11200 357434 11240
rect 360066 11200 360122 11240
rect 360610 11268 360666 12000
rect 360746 11268 360752 11280
rect 360610 11240 360752 11268
rect 360610 11200 360666 11240
rect 360746 11228 360752 11240
rect 360804 11228 360810 11280
rect 360930 11228 360936 11280
rect 360988 11268 360994 11280
rect 361154 11268 361210 12000
rect 360988 11240 361210 11268
rect 360988 11228 360994 11240
rect 361154 11200 361210 11240
rect 361298 11228 361304 11280
rect 361356 11268 361362 11280
rect 361698 11268 361754 12000
rect 361356 11240 361754 11268
rect 361356 11228 361362 11240
rect 361698 11200 361754 11240
rect 362034 11228 362040 11280
rect 362092 11268 362098 11280
rect 362242 11268 362298 12000
rect 362092 11240 362298 11268
rect 362092 11228 362098 11240
rect 362242 11200 362298 11240
rect 362402 11228 362408 11280
rect 362460 11268 362466 11280
rect 362786 11268 362842 12000
rect 363138 11432 363144 11484
rect 363196 11472 363202 11484
rect 363330 11472 363386 12000
rect 363196 11444 363386 11472
rect 363196 11432 363202 11444
rect 362460 11240 362842 11268
rect 362460 11228 362466 11240
rect 362786 11200 362842 11240
rect 363330 11200 363386 11444
rect 363690 11228 363696 11280
rect 363748 11268 363754 11280
rect 363874 11268 363930 12000
rect 363748 11240 363930 11268
rect 363748 11228 363754 11240
rect 363874 11200 363930 11240
rect 364242 11228 364248 11280
rect 364300 11268 364306 11280
rect 364418 11268 364474 12000
rect 364962 11268 365018 12000
rect 364300 11240 364474 11268
rect 364300 11228 364306 11240
rect 364418 11200 364474 11240
rect 364720 11240 365018 11268
rect 355520 11172 357434 11200
rect 258810 11092 258816 11144
rect 258868 11132 258874 11144
rect 355520 11132 355548 11172
rect 364518 11160 364524 11212
rect 364576 11200 364582 11212
rect 364720 11200 364748 11240
rect 364962 11200 365018 11240
rect 365254 11228 365260 11280
rect 365312 11268 365318 11280
rect 365506 11268 365562 12000
rect 365312 11240 365562 11268
rect 365312 11228 365318 11240
rect 365506 11200 365562 11240
rect 365806 11228 365812 11280
rect 365864 11268 365870 11280
rect 366050 11268 366106 12000
rect 365864 11240 366106 11268
rect 365864 11228 365870 11240
rect 366050 11200 366106 11240
rect 366358 11228 366364 11280
rect 366416 11268 366422 11280
rect 366594 11268 366650 12000
rect 366416 11240 366650 11268
rect 366416 11228 366422 11240
rect 366594 11200 366650 11240
rect 366726 11228 366732 11280
rect 366784 11268 366790 11280
rect 367138 11268 367194 12000
rect 366784 11240 367194 11268
rect 366784 11228 366790 11240
rect 367138 11200 367194 11240
rect 367462 11228 367468 11280
rect 367520 11268 367526 11280
rect 367682 11268 367738 12000
rect 367520 11240 367738 11268
rect 367520 11228 367526 11240
rect 367682 11200 367738 11240
rect 368014 11228 368020 11280
rect 368072 11268 368078 11280
rect 368226 11268 368282 12000
rect 368072 11240 368282 11268
rect 368072 11228 368078 11240
rect 368226 11200 368282 11240
rect 368658 11228 368664 11280
rect 368716 11268 368722 11280
rect 368770 11268 368826 12000
rect 369314 11268 369370 12000
rect 368716 11240 368826 11268
rect 368716 11228 368722 11240
rect 368770 11200 368826 11240
rect 368952 11240 369370 11268
rect 368952 11212 368980 11240
rect 364576 11172 364748 11200
rect 364576 11160 364582 11172
rect 368934 11160 368940 11212
rect 368992 11160 368998 11212
rect 369314 11200 369370 11240
rect 369762 11228 369768 11280
rect 369820 11268 369826 11280
rect 369858 11268 369914 12000
rect 369820 11240 369914 11268
rect 369820 11228 369826 11240
rect 369858 11200 369914 11240
rect 370130 11228 370136 11280
rect 370188 11268 370194 11280
rect 370402 11268 370458 12000
rect 370188 11240 370458 11268
rect 370188 11228 370194 11240
rect 370402 11200 370458 11240
rect 370682 11228 370688 11280
rect 370740 11268 370746 11280
rect 370946 11268 371002 12000
rect 370740 11240 371002 11268
rect 370740 11228 370746 11240
rect 370946 11200 371002 11240
rect 371050 11228 371056 11280
rect 371108 11268 371114 11280
rect 371490 11268 371546 12000
rect 371108 11240 371546 11268
rect 371108 11228 371114 11240
rect 371490 11200 371546 11240
rect 371786 11228 371792 11280
rect 371844 11268 371850 11280
rect 372034 11268 372090 12000
rect 371844 11240 372090 11268
rect 371844 11228 371850 11240
rect 372034 11200 372090 11240
rect 372154 11228 372160 11280
rect 372212 11268 372218 11280
rect 372578 11268 372634 12000
rect 372212 11240 372634 11268
rect 372212 11228 372218 11240
rect 372578 11200 372634 11240
rect 372890 11228 372896 11280
rect 372948 11268 372954 11280
rect 373122 11268 373178 12000
rect 372948 11240 373178 11268
rect 372948 11228 372954 11240
rect 373122 11200 373178 11240
rect 373258 11228 373264 11280
rect 373316 11268 373322 11280
rect 373666 11268 373722 12000
rect 373316 11240 373722 11268
rect 373316 11228 373322 11240
rect 373666 11200 373722 11240
rect 373994 11228 374000 11280
rect 374052 11268 374058 11280
rect 374210 11268 374266 12000
rect 374052 11240 374266 11268
rect 374052 11228 374058 11240
rect 374210 11200 374266 11240
rect 374362 11228 374368 11280
rect 374420 11268 374426 11280
rect 374754 11268 374810 12000
rect 374420 11240 374810 11268
rect 374420 11228 374426 11240
rect 374754 11200 374810 11240
rect 375098 11228 375104 11280
rect 375156 11268 375162 11280
rect 375298 11268 375354 12000
rect 375156 11240 375354 11268
rect 375156 11228 375162 11240
rect 375298 11200 375354 11240
rect 375466 11228 375472 11280
rect 375524 11268 375530 11280
rect 375842 11268 375898 12000
rect 375524 11240 375898 11268
rect 375524 11228 375530 11240
rect 375842 11200 375898 11240
rect 376202 11228 376208 11280
rect 376260 11268 376266 11280
rect 376386 11268 376442 12000
rect 376260 11240 376442 11268
rect 376260 11228 376266 11240
rect 376386 11200 376442 11240
rect 376930 11268 376986 12000
rect 377030 11268 377036 11280
rect 376930 11240 377036 11268
rect 376930 11200 376986 11240
rect 377030 11228 377036 11240
rect 377088 11228 377094 11280
rect 377306 11228 377312 11280
rect 377364 11268 377370 11280
rect 377474 11268 377530 12000
rect 377364 11240 377530 11268
rect 377364 11228 377370 11240
rect 377474 11200 377530 11240
rect 377582 11228 377588 11280
rect 377640 11268 377646 11280
rect 378018 11268 378074 12000
rect 377640 11240 378074 11268
rect 377640 11228 377646 11240
rect 378018 11200 378074 11240
rect 378410 11228 378416 11280
rect 378468 11268 378474 11280
rect 378562 11268 378618 12000
rect 378468 11240 378618 11268
rect 378468 11228 378474 11240
rect 378562 11200 378618 11240
rect 378686 11228 378692 11280
rect 378744 11268 378750 11280
rect 379106 11268 379162 12000
rect 378744 11240 379162 11268
rect 378744 11228 378750 11240
rect 379106 11200 379162 11240
rect 379422 11228 379428 11280
rect 379480 11268 379486 11280
rect 379650 11268 379706 12000
rect 380194 11268 380250 12000
rect 379480 11240 379706 11268
rect 379480 11228 379486 11240
rect 379650 11200 379706 11240
rect 380176 11200 380250 11268
rect 380342 11228 380348 11280
rect 380400 11268 380406 11280
rect 380738 11268 380794 12000
rect 381282 11268 381338 12000
rect 380400 11240 380794 11268
rect 380400 11228 380406 11240
rect 380738 11200 380794 11240
rect 381188 11240 381338 11268
rect 258868 11104 355548 11132
rect 258868 11092 258874 11104
rect 355778 11092 355784 11144
rect 355836 11132 355842 11144
rect 355836 11104 362540 11132
rect 355836 11092 355842 11104
rect 354490 11064 354496 11076
rect 260944 11036 354496 11064
rect 260834 10792 260840 10804
rect 248748 10764 258764 10792
rect 258828 10764 260840 10792
rect 248748 10752 248754 10764
rect 220136 10696 241514 10724
rect 220136 10684 220142 10696
rect 251174 10684 251180 10736
rect 251232 10724 251238 10736
rect 255314 10724 255320 10736
rect 251232 10696 255320 10724
rect 251232 10684 251238 10696
rect 255314 10684 255320 10696
rect 255372 10684 255378 10736
rect 258828 10724 258856 10764
rect 260834 10752 260840 10764
rect 260892 10752 260898 10804
rect 257356 10696 258856 10724
rect 195238 10616 195244 10668
rect 195296 10656 195302 10668
rect 198642 10656 198648 10668
rect 195296 10628 198648 10656
rect 195296 10616 195302 10628
rect 198642 10616 198648 10628
rect 198700 10616 198706 10668
rect 198734 10616 198740 10668
rect 198792 10656 198798 10668
rect 201494 10656 201500 10668
rect 198792 10628 201500 10656
rect 198792 10616 198798 10628
rect 201494 10616 201500 10628
rect 201552 10616 201558 10668
rect 202874 10616 202880 10668
rect 202932 10656 202938 10668
rect 205082 10656 205088 10668
rect 202932 10628 205088 10656
rect 202932 10616 202938 10628
rect 205082 10616 205088 10628
rect 205140 10616 205146 10668
rect 205174 10616 205180 10668
rect 205232 10656 205238 10668
rect 257356 10656 257384 10696
rect 205232 10628 257384 10656
rect 205232 10616 205238 10628
rect 106182 10548 106188 10600
rect 106240 10588 106246 10600
rect 206002 10588 206008 10600
rect 106240 10560 206008 10588
rect 106240 10548 106246 10560
rect 206002 10548 206008 10560
rect 206060 10548 206066 10600
rect 206094 10548 206100 10600
rect 206152 10588 206158 10600
rect 212718 10588 212724 10600
rect 206152 10560 212724 10588
rect 206152 10548 206158 10560
rect 212718 10548 212724 10560
rect 212776 10548 212782 10600
rect 213270 10548 213276 10600
rect 213328 10588 213334 10600
rect 219986 10588 219992 10600
rect 213328 10560 219992 10588
rect 213328 10548 213334 10560
rect 219986 10548 219992 10560
rect 220044 10548 220050 10600
rect 224926 10560 225092 10588
rect 109862 10480 109868 10532
rect 109920 10520 109926 10532
rect 206830 10520 206836 10532
rect 109920 10492 206836 10520
rect 109920 10480 109926 10492
rect 206830 10480 206836 10492
rect 206888 10480 206894 10532
rect 206922 10480 206928 10532
rect 206980 10520 206986 10532
rect 211154 10520 211160 10532
rect 206980 10492 211160 10520
rect 206980 10480 206986 10492
rect 211154 10480 211160 10492
rect 211212 10480 211218 10532
rect 211246 10480 211252 10532
rect 211304 10520 211310 10532
rect 217870 10520 217876 10532
rect 211304 10492 217876 10520
rect 211304 10480 211310 10492
rect 217870 10480 217876 10492
rect 217928 10480 217934 10532
rect 218790 10480 218796 10532
rect 218848 10520 218854 10532
rect 224926 10520 224954 10560
rect 218848 10492 224954 10520
rect 225064 10520 225092 10560
rect 225138 10548 225144 10600
rect 225196 10588 225202 10600
rect 238938 10588 238944 10600
rect 225196 10560 238944 10588
rect 225196 10548 225202 10560
rect 238938 10548 238944 10560
rect 238996 10548 239002 10600
rect 239398 10548 239404 10600
rect 239456 10588 239462 10600
rect 245378 10588 245384 10600
rect 239456 10560 245384 10588
rect 239456 10548 239462 10560
rect 245378 10548 245384 10560
rect 245436 10548 245442 10600
rect 250806 10548 250812 10600
rect 250864 10588 250870 10600
rect 258810 10588 258816 10600
rect 250864 10560 258816 10588
rect 250864 10548 250870 10560
rect 258810 10548 258816 10560
rect 258868 10548 258874 10600
rect 229738 10520 229744 10532
rect 225064 10492 229744 10520
rect 218848 10480 218854 10492
rect 229738 10480 229744 10492
rect 229796 10480 229802 10532
rect 238846 10480 238852 10532
rect 238904 10520 238910 10532
rect 246942 10520 246948 10532
rect 238904 10492 246948 10520
rect 238904 10480 238910 10492
rect 246942 10480 246948 10492
rect 247000 10480 247006 10532
rect 247218 10480 247224 10532
rect 247276 10520 247282 10532
rect 258718 10520 258724 10532
rect 247276 10492 258724 10520
rect 247276 10480 247282 10492
rect 258718 10480 258724 10492
rect 258776 10480 258782 10532
rect 122558 10412 122564 10464
rect 122616 10452 122622 10464
rect 199286 10452 199292 10464
rect 122616 10424 199292 10452
rect 122616 10412 122622 10424
rect 199286 10412 199292 10424
rect 199344 10412 199350 10464
rect 199378 10412 199384 10464
rect 199436 10452 199442 10464
rect 203426 10452 203432 10464
rect 199436 10424 203432 10452
rect 199436 10412 199442 10424
rect 203426 10412 203432 10424
rect 203484 10412 203490 10464
rect 203518 10412 203524 10464
rect 203576 10452 203582 10464
rect 205174 10452 205180 10464
rect 203576 10424 205180 10452
rect 203576 10412 203582 10424
rect 205174 10412 205180 10424
rect 205232 10412 205238 10464
rect 205634 10412 205640 10464
rect 205692 10452 205698 10464
rect 209958 10452 209964 10464
rect 205692 10424 209964 10452
rect 205692 10412 205698 10424
rect 209958 10412 209964 10424
rect 210016 10412 210022 10464
rect 210234 10412 210240 10464
rect 210292 10452 210298 10464
rect 240410 10452 240416 10464
rect 210292 10424 240416 10452
rect 210292 10412 210298 10424
rect 240410 10412 240416 10424
rect 240468 10412 240474 10464
rect 241514 10412 241520 10464
rect 241572 10452 241578 10464
rect 251910 10452 251916 10464
rect 241572 10424 251916 10452
rect 241572 10412 241578 10424
rect 251910 10412 251916 10424
rect 251968 10412 251974 10464
rect 256970 10412 256976 10464
rect 257028 10452 257034 10464
rect 260944 10452 260972 11036
rect 354490 11024 354496 11036
rect 354548 11024 354554 11076
rect 362402 11064 362408 11076
rect 354600 11036 362408 11064
rect 262030 10956 262036 11008
rect 262088 10996 262094 11008
rect 354600 10996 354628 11036
rect 362402 11024 362408 11036
rect 362460 11024 362466 11076
rect 362512 11064 362540 11104
rect 362586 11092 362592 11144
rect 362644 11132 362650 11144
rect 362644 11104 379514 11132
rect 362644 11092 362650 11104
rect 362512 11036 368152 11064
rect 361390 10996 361396 11008
rect 262088 10968 354628 10996
rect 355336 10968 361396 10996
rect 262088 10956 262094 10968
rect 267090 10888 267096 10940
rect 267148 10928 267154 10940
rect 355336 10928 355364 10968
rect 361390 10956 361396 10968
rect 361448 10956 361454 11008
rect 363414 10956 363420 11008
rect 363472 10996 363478 11008
rect 368014 10996 368020 11008
rect 363472 10968 368020 10996
rect 363472 10956 363478 10968
rect 368014 10956 368020 10968
rect 368072 10956 368078 11008
rect 368124 10996 368152 11036
rect 368124 10968 374776 10996
rect 267148 10900 355364 10928
rect 267148 10888 267154 10900
rect 355410 10888 355416 10940
rect 355468 10928 355474 10940
rect 362586 10928 362592 10940
rect 355468 10900 362592 10928
rect 355468 10888 355474 10900
rect 362586 10888 362592 10900
rect 362644 10888 362650 10940
rect 364978 10888 364984 10940
rect 365036 10928 365042 10940
rect 365036 10900 371004 10928
rect 365036 10888 365042 10900
rect 272150 10820 272156 10872
rect 272208 10860 272214 10872
rect 360286 10860 360292 10872
rect 272208 10832 360292 10860
rect 272208 10820 272214 10832
rect 360286 10820 360292 10832
rect 360344 10820 360350 10872
rect 363322 10820 363328 10872
rect 363380 10860 363386 10872
rect 368934 10860 368940 10872
rect 363380 10832 368940 10860
rect 363380 10820 363386 10832
rect 368934 10820 368940 10832
rect 368992 10820 368998 10872
rect 354490 10752 354496 10804
rect 354548 10792 354554 10804
rect 359550 10792 359556 10804
rect 354548 10764 359556 10792
rect 354548 10752 354554 10764
rect 359550 10752 359556 10764
rect 359608 10752 359614 10804
rect 361390 10752 361396 10804
rect 361448 10792 361454 10804
rect 363690 10792 363696 10804
rect 361448 10764 363696 10792
rect 361448 10752 361454 10764
rect 363690 10752 363696 10764
rect 363748 10752 363754 10804
rect 364150 10752 364156 10804
rect 364208 10792 364214 10804
rect 364208 10764 364656 10792
rect 364208 10752 364214 10764
rect 282270 10684 282276 10736
rect 282328 10724 282334 10736
rect 360102 10724 360108 10736
rect 282328 10696 360108 10724
rect 282328 10684 282334 10696
rect 360102 10684 360108 10696
rect 360160 10684 360166 10736
rect 360654 10684 360660 10736
rect 360712 10724 360718 10736
rect 364518 10724 364524 10736
rect 360712 10696 364524 10724
rect 360712 10684 360718 10696
rect 364518 10684 364524 10696
rect 364576 10684 364582 10736
rect 364628 10724 364656 10764
rect 370976 10724 371004 10900
rect 374748 10860 374776 10968
rect 379486 10928 379514 11104
rect 380176 11064 380204 11200
rect 381188 11132 381216 11240
rect 381282 11200 381338 11240
rect 381538 11228 381544 11280
rect 381596 11268 381602 11280
rect 381826 11268 381882 12000
rect 381596 11240 381882 11268
rect 381596 11228 381602 11240
rect 381826 11200 381882 11240
rect 382090 11228 382096 11280
rect 382148 11268 382154 11280
rect 382370 11268 382426 12000
rect 382148 11240 382426 11268
rect 382148 11228 382154 11240
rect 382370 11200 382426 11240
rect 382458 11228 382464 11280
rect 382516 11268 382522 11280
rect 382914 11268 382970 12000
rect 382516 11240 382970 11268
rect 382516 11228 382522 11240
rect 382914 11200 382970 11240
rect 383194 11228 383200 11280
rect 383252 11268 383258 11280
rect 383458 11268 383514 12000
rect 384002 11268 384058 12000
rect 383252 11240 383514 11268
rect 383252 11228 383258 11240
rect 383458 11200 383514 11240
rect 383672 11240 384058 11268
rect 383672 11132 383700 11240
rect 384002 11200 384058 11240
rect 384546 11268 384602 12000
rect 381188 11104 381324 11132
rect 380176 11036 380250 11064
rect 380222 10928 380250 11036
rect 379486 10900 380250 10928
rect 381296 10860 381324 11104
rect 374748 10832 381324 10860
rect 383028 11104 383700 11132
rect 384546 11172 384620 11268
rect 384666 11228 384672 11280
rect 384724 11268 384730 11280
rect 385090 11268 385146 12000
rect 384724 11240 385146 11268
rect 384724 11228 384730 11240
rect 385090 11200 385146 11240
rect 385218 11228 385224 11280
rect 385276 11268 385282 11280
rect 385634 11268 385690 12000
rect 385276 11240 385690 11268
rect 385276 11228 385282 11240
rect 385634 11200 385690 11240
rect 385954 11228 385960 11280
rect 386012 11268 386018 11280
rect 386178 11268 386234 12000
rect 386012 11240 386234 11268
rect 386012 11228 386018 11240
rect 386178 11200 386234 11240
rect 386506 11228 386512 11280
rect 386564 11268 386570 11280
rect 386722 11268 386778 12000
rect 387266 11268 387322 12000
rect 386564 11240 386778 11268
rect 386564 11228 386570 11240
rect 386722 11200 386778 11240
rect 386984 11240 387322 11268
rect 374454 10752 374460 10804
rect 374512 10792 374518 10804
rect 380342 10792 380348 10804
rect 374512 10764 380348 10792
rect 374512 10752 374518 10764
rect 380342 10752 380348 10764
rect 380400 10752 380406 10804
rect 381538 10724 381544 10736
rect 364628 10696 369854 10724
rect 370976 10696 381544 10724
rect 287422 10616 287428 10668
rect 287480 10656 287486 10668
rect 287480 10628 360516 10656
rect 287480 10616 287486 10628
rect 292574 10548 292580 10600
rect 292632 10588 292638 10600
rect 360194 10588 360200 10600
rect 292632 10560 360200 10588
rect 292632 10548 292638 10560
rect 360194 10548 360200 10560
rect 360252 10548 360258 10600
rect 360488 10588 360516 10628
rect 360562 10616 360568 10668
rect 360620 10656 360626 10668
rect 365806 10656 365812 10668
rect 360620 10628 365812 10656
rect 360620 10616 360626 10628
rect 365806 10616 365812 10628
rect 365864 10616 365870 10668
rect 369826 10656 369854 10696
rect 381538 10684 381544 10696
rect 381596 10684 381602 10736
rect 382458 10656 382464 10668
rect 369826 10628 382464 10656
rect 382458 10616 382464 10628
rect 382516 10616 382522 10668
rect 363414 10588 363420 10600
rect 360488 10560 363420 10588
rect 363414 10548 363420 10560
rect 363472 10548 363478 10600
rect 367094 10548 367100 10600
rect 367152 10588 367158 10600
rect 374454 10588 374460 10600
rect 367152 10560 374460 10588
rect 367152 10548 367158 10560
rect 374454 10548 374460 10560
rect 374512 10548 374518 10600
rect 379974 10548 379980 10600
rect 380032 10588 380038 10600
rect 383028 10588 383056 11104
rect 383562 10956 383568 11008
rect 383620 10996 383626 11008
rect 384546 10996 384574 11172
rect 385862 11092 385868 11144
rect 385920 11132 385926 11144
rect 386984 11132 387012 11240
rect 387266 11200 387322 11240
rect 387810 11268 387866 12000
rect 387978 11268 387984 11280
rect 387810 11240 387984 11268
rect 387810 11200 387866 11240
rect 387978 11228 387984 11240
rect 388036 11228 388042 11280
rect 388354 11268 388410 12000
rect 388898 11336 388954 12000
rect 388088 11240 388410 11268
rect 385920 11104 387012 11132
rect 385920 11092 385926 11104
rect 387058 11092 387064 11144
rect 387116 11132 387122 11144
rect 388088 11132 388116 11240
rect 388354 11200 388410 11240
rect 388640 11308 388954 11336
rect 387116 11104 388116 11132
rect 387116 11092 387122 11104
rect 385770 11024 385776 11076
rect 385828 11064 385834 11076
rect 388640 11064 388668 11308
rect 388898 11200 388954 11308
rect 389442 11268 389498 12000
rect 389146 11240 389498 11268
rect 388990 11160 388996 11212
rect 389048 11200 389054 11212
rect 389146 11200 389174 11240
rect 389442 11200 389498 11240
rect 389818 11228 389824 11280
rect 389876 11268 389882 11280
rect 389986 11268 390042 12000
rect 389876 11240 390042 11268
rect 389876 11228 389882 11240
rect 389986 11200 390042 11240
rect 390530 11268 390586 12000
rect 390646 11268 390652 11280
rect 390530 11240 390652 11268
rect 390530 11200 390586 11240
rect 390646 11228 390652 11240
rect 390704 11228 390710 11280
rect 391074 11268 391130 12000
rect 391074 11200 391152 11268
rect 391382 11228 391388 11280
rect 391440 11268 391446 11280
rect 391618 11268 391674 12000
rect 391440 11240 391674 11268
rect 391440 11228 391446 11240
rect 391618 11200 391674 11240
rect 391934 11228 391940 11280
rect 391992 11268 391998 11280
rect 392162 11268 392218 12000
rect 391992 11240 392218 11268
rect 391992 11228 391998 11240
rect 392162 11200 392218 11240
rect 392486 11228 392492 11280
rect 392544 11268 392550 11280
rect 392706 11268 392762 12000
rect 392544 11240 392762 11268
rect 392544 11228 392550 11240
rect 392706 11200 392762 11240
rect 392854 11228 392860 11280
rect 392912 11268 392918 11280
rect 393250 11268 393306 12000
rect 392912 11240 393306 11268
rect 392912 11228 392918 11240
rect 393250 11200 393306 11240
rect 393498 11228 393504 11280
rect 393556 11268 393562 11280
rect 393794 11268 393850 12000
rect 393556 11240 393850 11268
rect 393556 11228 393562 11240
rect 393794 11200 393850 11240
rect 394050 11228 394056 11280
rect 394108 11268 394114 11280
rect 394338 11268 394394 12000
rect 394108 11240 394394 11268
rect 394108 11228 394114 11240
rect 394338 11200 394394 11240
rect 394694 11228 394700 11280
rect 394752 11268 394758 11280
rect 394882 11268 394938 12000
rect 394752 11240 394938 11268
rect 394752 11228 394758 11240
rect 394882 11200 394938 11240
rect 395154 11228 395160 11280
rect 395212 11268 395218 11280
rect 395426 11268 395482 12000
rect 395212 11240 395482 11268
rect 395212 11228 395218 11240
rect 395426 11200 395482 11240
rect 395522 11228 395528 11280
rect 395580 11268 395586 11280
rect 395970 11268 396026 12000
rect 395580 11240 396026 11268
rect 395580 11228 395586 11240
rect 395970 11200 396026 11240
rect 396258 11228 396264 11280
rect 396316 11268 396322 11280
rect 396514 11268 396570 12000
rect 396316 11240 396570 11268
rect 396316 11228 396322 11240
rect 396514 11200 396570 11240
rect 397058 11268 397114 12000
rect 397602 11268 397658 12000
rect 389048 11172 389174 11200
rect 389048 11160 389054 11172
rect 391124 11132 391152 11200
rect 385828 11036 388668 11064
rect 391078 11104 391152 11132
rect 397058 11172 397132 11268
rect 397602 11200 397684 11268
rect 397914 11228 397920 11280
rect 397972 11268 397978 11280
rect 398146 11268 398202 12000
rect 397972 11240 398202 11268
rect 397972 11228 397978 11240
rect 398146 11200 398202 11240
rect 398466 11228 398472 11280
rect 398524 11268 398530 11280
rect 398690 11268 398746 12000
rect 399234 11268 399290 12000
rect 398524 11240 398746 11268
rect 398524 11228 398530 11240
rect 398690 11200 398746 11240
rect 399128 11240 399290 11268
rect 385828 11024 385834 11036
rect 383620 10968 384574 10996
rect 383620 10956 383626 10968
rect 390554 10956 390560 11008
rect 390612 10996 390618 11008
rect 391078 10996 391106 11104
rect 390612 10968 391106 10996
rect 390612 10956 390618 10968
rect 396074 10956 396080 11008
rect 396132 10996 396138 11008
rect 397058 10996 397086 11172
rect 397656 11132 397684 11200
rect 397610 11104 397684 11132
rect 399128 11132 399156 11240
rect 399234 11200 399290 11240
rect 399778 11268 399834 12000
rect 400322 11268 400378 12000
rect 399778 11240 399892 11268
rect 399778 11200 399834 11240
rect 399864 11144 399892 11240
rect 400232 11240 400378 11268
rect 399294 11132 399300 11144
rect 399128 11104 399300 11132
rect 396132 10968 397086 10996
rect 396132 10956 396138 10968
rect 397454 10956 397460 11008
rect 397512 10996 397518 11008
rect 397610 10996 397638 11104
rect 399294 11092 399300 11104
rect 399352 11092 399358 11144
rect 399846 11092 399852 11144
rect 399904 11092 399910 11144
rect 400232 11132 400260 11240
rect 400322 11200 400378 11240
rect 400674 11228 400680 11280
rect 400732 11268 400738 11280
rect 400866 11268 400922 12000
rect 400732 11240 400922 11268
rect 400732 11228 400738 11240
rect 400866 11200 400922 11240
rect 400950 11228 400956 11280
rect 401008 11268 401014 11280
rect 401410 11268 401466 12000
rect 401954 11268 402010 12000
rect 401008 11240 401466 11268
rect 401008 11228 401014 11240
rect 401410 11200 401466 11240
rect 401888 11240 402010 11268
rect 401888 11132 401916 11240
rect 401954 11200 402010 11240
rect 402330 11228 402336 11280
rect 402388 11268 402394 11280
rect 402498 11268 402554 12000
rect 402388 11240 402554 11268
rect 402388 11228 402394 11240
rect 402498 11200 402554 11240
rect 403042 11268 403098 12000
rect 403586 11268 403642 12000
rect 403042 11240 403204 11268
rect 403042 11200 403098 11240
rect 403176 11132 403204 11240
rect 403586 11200 403664 11268
rect 403894 11228 403900 11280
rect 403952 11268 403958 11280
rect 404130 11268 404186 12000
rect 403952 11240 404186 11268
rect 403952 11228 403958 11240
rect 404130 11200 404186 11240
rect 438854 11228 438860 11280
rect 438912 11268 438918 11280
rect 440034 11268 440090 12000
rect 438912 11240 440090 11268
rect 438912 11228 438918 11240
rect 440034 11200 440090 11240
rect 440142 11228 440148 11280
rect 440200 11268 440206 11280
rect 440306 11268 440362 12000
rect 440200 11240 440362 11268
rect 440200 11228 440206 11240
rect 440306 11200 440362 11240
rect 440418 11228 440424 11280
rect 440476 11268 440482 11280
rect 440578 11268 440634 12000
rect 440476 11240 440634 11268
rect 440476 11228 440482 11240
rect 440578 11200 440634 11240
rect 440694 11228 440700 11280
rect 440752 11268 440758 11280
rect 440850 11268 440906 12000
rect 440752 11240 440906 11268
rect 440752 11228 440758 11240
rect 440850 11200 440906 11240
rect 441122 11268 441178 12000
rect 441394 11268 441450 12000
rect 441666 11336 441722 12000
rect 441586 11308 441722 11336
rect 441122 11200 441200 11268
rect 441394 11200 441476 11268
rect 400232 11104 400352 11132
rect 401888 11104 402008 11132
rect 400324 11008 400352 11104
rect 401980 11008 402008 11104
rect 403056 11104 403204 11132
rect 403590 11172 403664 11200
rect 403056 11008 403084 11104
rect 403590 11008 403618 11172
rect 441172 11132 441200 11200
rect 441448 11132 441476 11200
rect 441126 11104 441200 11132
rect 441402 11104 441476 11132
rect 441586 11132 441614 11308
rect 441666 11200 441722 11308
rect 441798 11296 441804 11348
rect 441856 11336 441862 11348
rect 441938 11336 441994 12000
rect 441856 11308 441994 11336
rect 441856 11296 441862 11308
rect 441938 11200 441994 11308
rect 442210 11268 442266 12000
rect 442482 11268 442538 12000
rect 442754 11268 442810 12000
rect 442902 11296 442908 11348
rect 442960 11336 442966 11348
rect 443026 11336 443082 12000
rect 442960 11308 443082 11336
rect 442960 11296 442966 11308
rect 442184 11200 442266 11268
rect 442460 11200 442538 11268
rect 442184 11172 442258 11200
rect 442460 11172 442534 11200
rect 442736 11172 442810 11268
rect 443026 11200 443082 11308
rect 443178 11228 443184 11280
rect 443236 11268 443242 11280
rect 443298 11268 443354 12000
rect 443236 11240 443354 11268
rect 443236 11228 443242 11240
rect 443298 11200 443354 11240
rect 443454 11228 443460 11280
rect 443512 11268 443518 11280
rect 443570 11268 443626 12000
rect 443512 11240 443626 11268
rect 443512 11228 443518 11240
rect 443570 11200 443626 11240
rect 443842 11268 443898 12000
rect 443842 11240 443960 11268
rect 443842 11200 443898 11240
rect 441586 11104 441706 11132
rect 440326 11024 440332 11076
rect 440384 11064 440390 11076
rect 441126 11064 441154 11104
rect 440384 11036 441154 11064
rect 440384 11024 440390 11036
rect 397512 10968 397638 10996
rect 397512 10956 397518 10968
rect 400306 10956 400312 11008
rect 400364 10956 400370 11008
rect 401962 10956 401968 11008
rect 402020 10956 402026 11008
rect 403056 10968 403072 11008
rect 403066 10956 403072 10968
rect 403124 10956 403130 11008
rect 403590 10968 403624 11008
rect 403618 10956 403624 10968
rect 403676 10956 403682 11008
rect 440234 10956 440240 11008
rect 440292 10996 440298 11008
rect 441402 10996 441430 11104
rect 441678 11008 441706 11104
rect 440292 10968 441430 10996
rect 440292 10956 440298 10968
rect 441614 10956 441620 11008
rect 441672 10968 441706 11008
rect 441672 10956 441678 10968
rect 442074 10956 442080 11008
rect 442132 10996 442138 11008
rect 442230 10996 442258 11172
rect 442132 10968 442258 10996
rect 442132 10956 442138 10968
rect 441706 10888 441712 10940
rect 441764 10928 441770 10940
rect 442506 10928 442534 11172
rect 442626 10956 442632 11008
rect 442684 10996 442690 11008
rect 442782 10996 442810 11172
rect 443932 11132 443960 11240
rect 444006 11228 444012 11280
rect 444064 11268 444070 11280
rect 444114 11268 444170 12000
rect 444064 11240 444170 11268
rect 444064 11228 444070 11240
rect 444114 11200 444170 11240
rect 444386 11268 444442 12000
rect 444386 11240 444512 11268
rect 444386 11200 444442 11240
rect 444484 11132 444512 11240
rect 444558 11228 444564 11280
rect 444616 11268 444622 11280
rect 444658 11268 444714 12000
rect 444616 11240 444714 11268
rect 444616 11228 444622 11240
rect 444658 11200 444714 11240
rect 444742 11228 444748 11280
rect 444800 11268 444806 11280
rect 444930 11268 444986 12000
rect 444800 11240 444986 11268
rect 444800 11228 444806 11240
rect 444930 11200 444986 11240
rect 445018 11228 445024 11280
rect 445076 11268 445082 11280
rect 445202 11268 445258 12000
rect 445076 11240 445258 11268
rect 445076 11228 445082 11240
rect 445202 11200 445258 11240
rect 445294 11228 445300 11280
rect 445352 11268 445358 11280
rect 445474 11268 445530 12000
rect 445352 11240 445530 11268
rect 445352 11228 445358 11240
rect 445474 11200 445530 11240
rect 445746 11404 445802 12000
rect 445846 11404 445852 11416
rect 445746 11376 445852 11404
rect 445746 11200 445802 11376
rect 445846 11364 445852 11376
rect 445904 11364 445910 11416
rect 445846 11228 445852 11280
rect 445904 11268 445910 11280
rect 446018 11268 446074 12000
rect 445904 11240 446074 11268
rect 445904 11228 445910 11240
rect 446018 11200 446074 11240
rect 446122 11228 446128 11280
rect 446180 11268 446186 11280
rect 446290 11268 446346 12000
rect 446180 11240 446346 11268
rect 446180 11228 446186 11240
rect 446290 11200 446346 11240
rect 446562 11540 446618 12000
rect 446674 11540 446680 11552
rect 446562 11512 446680 11540
rect 446562 11200 446618 11512
rect 446674 11500 446680 11512
rect 446732 11500 446738 11552
rect 446674 11296 446680 11348
rect 446732 11336 446738 11348
rect 446834 11336 446890 12000
rect 446732 11308 446890 11336
rect 446732 11296 446738 11308
rect 446834 11200 446890 11308
rect 447106 11268 447162 12000
rect 447378 11268 447434 12000
rect 447650 11268 447706 12000
rect 447778 11296 447784 11348
rect 447836 11336 447842 11348
rect 447922 11336 447978 12000
rect 447836 11308 447978 11336
rect 447836 11296 447842 11308
rect 443856 11104 443960 11132
rect 444392 11104 444512 11132
rect 447106 11172 447180 11268
rect 447378 11200 447456 11268
rect 447650 11200 447732 11268
rect 447922 11200 447978 11308
rect 448054 11296 448060 11348
rect 448112 11336 448118 11348
rect 448194 11336 448250 12000
rect 448112 11308 448250 11336
rect 448112 11296 448118 11308
rect 448194 11200 448250 11308
rect 448466 11268 448522 12000
rect 480018 11268 480074 12000
rect 480290 11268 480346 12000
rect 480562 11268 480618 12000
rect 448440 11200 448522 11268
rect 479996 11200 480074 11268
rect 442684 10968 442810 10996
rect 442684 10956 442690 10968
rect 443086 10956 443092 11008
rect 443144 10996 443150 11008
rect 443856 10996 443884 11104
rect 443144 10968 443884 10996
rect 443144 10956 443150 10968
rect 444392 10940 444420 11104
rect 447106 11008 447134 11172
rect 447428 11132 447456 11200
rect 447382 11104 447456 11132
rect 447658 11172 447732 11200
rect 448440 11172 448514 11200
rect 479996 11172 480070 11200
rect 480272 11172 480346 11268
rect 447106 10968 447140 11008
rect 447134 10956 447140 10968
rect 447192 10956 447198 11008
rect 441764 10900 442534 10928
rect 441764 10888 441770 10900
rect 444374 10888 444380 10940
rect 444432 10888 444438 10940
rect 447226 10888 447232 10940
rect 447284 10928 447290 10940
rect 447382 10928 447410 11104
rect 447658 11008 447686 11172
rect 447658 10968 447692 11008
rect 447686 10956 447692 10968
rect 447744 10956 447750 11008
rect 447284 10900 447410 10928
rect 447284 10888 447290 10900
rect 448330 10888 448336 10940
rect 448388 10928 448394 10940
rect 448486 10928 448514 11172
rect 478874 10956 478880 11008
rect 478932 10996 478938 11008
rect 480042 10996 480070 11172
rect 478932 10968 480070 10996
rect 480318 11008 480346 11172
rect 480456 11240 480618 11268
rect 480456 11132 480484 11240
rect 480562 11200 480618 11240
rect 480714 11228 480720 11280
rect 480772 11268 480778 11280
rect 480834 11268 480890 12000
rect 480772 11240 480890 11268
rect 480772 11228 480778 11240
rect 480834 11200 480890 11240
rect 481106 11268 481162 12000
rect 481106 11240 481220 11268
rect 481106 11200 481162 11240
rect 481192 11144 481220 11240
rect 481266 11228 481272 11280
rect 481324 11268 481330 11280
rect 481378 11268 481434 12000
rect 481324 11240 481434 11268
rect 481324 11228 481330 11240
rect 481378 11200 481434 11240
rect 481650 11268 481706 12000
rect 481818 11296 481824 11348
rect 481876 11336 481882 11348
rect 481922 11336 481978 12000
rect 481876 11308 481978 11336
rect 481876 11296 481882 11308
rect 481650 11240 481772 11268
rect 481650 11200 481706 11240
rect 480456 11104 480604 11132
rect 480318 10968 480352 11008
rect 478932 10956 478938 10968
rect 480346 10956 480352 10968
rect 480404 10956 480410 11008
rect 448388 10900 448514 10928
rect 448388 10888 448394 10900
rect 480254 10888 480260 10940
rect 480312 10928 480318 10940
rect 480576 10928 480604 11104
rect 481174 11092 481180 11144
rect 481232 11092 481238 11144
rect 481744 11132 481772 11240
rect 481922 11200 481978 11308
rect 482094 11228 482100 11280
rect 482152 11268 482158 11280
rect 482194 11268 482250 12000
rect 482152 11240 482250 11268
rect 482152 11228 482158 11240
rect 482194 11200 482250 11240
rect 482278 11228 482284 11280
rect 482336 11268 482342 11280
rect 482466 11268 482522 12000
rect 482336 11240 482522 11268
rect 482336 11228 482342 11240
rect 482466 11200 482522 11240
rect 482738 11336 482794 12000
rect 482830 11336 482836 11348
rect 482738 11308 482836 11336
rect 482738 11200 482794 11308
rect 482830 11296 482836 11308
rect 482888 11296 482894 11348
rect 483010 11268 483066 12000
rect 483106 11296 483112 11348
rect 483164 11336 483170 11348
rect 483282 11336 483338 12000
rect 483164 11308 483338 11336
rect 483164 11296 483170 11308
rect 482986 11200 483066 11268
rect 483282 11200 483338 11308
rect 483554 11404 483610 12000
rect 483658 11404 483664 11416
rect 483554 11376 483664 11404
rect 483554 11200 483610 11376
rect 483658 11364 483664 11376
rect 483716 11364 483722 11416
rect 483658 11228 483664 11280
rect 483716 11268 483722 11280
rect 483826 11268 483882 12000
rect 484098 11336 484154 12000
rect 483716 11240 483882 11268
rect 483716 11228 483722 11240
rect 483826 11200 483882 11240
rect 483952 11308 484154 11336
rect 482986 11172 483152 11200
rect 481652 11104 481772 11132
rect 481652 10940 481680 11104
rect 480312 10900 480604 10928
rect 480312 10888 480318 10900
rect 481634 10888 481640 10940
rect 481692 10888 481698 10940
rect 483014 10888 483020 10940
rect 483072 10928 483078 10940
rect 483124 10928 483152 11172
rect 483952 11132 483980 11308
rect 484098 11200 484154 11308
rect 484210 11228 484216 11280
rect 484268 11268 484274 11280
rect 484370 11268 484426 12000
rect 484486 11296 484492 11348
rect 484544 11336 484550 11348
rect 484642 11336 484698 12000
rect 484544 11308 484698 11336
rect 484544 11296 484550 11308
rect 484268 11240 484426 11268
rect 484268 11228 484274 11240
rect 484370 11200 484426 11240
rect 484642 11200 484698 11308
rect 484914 11268 484970 12000
rect 485186 11268 485242 12000
rect 485458 11336 485514 12000
rect 485730 11336 485786 12000
rect 485332 11308 485514 11336
rect 484914 11200 484992 11268
rect 485186 11200 485268 11268
rect 484918 11172 484992 11200
rect 483952 11104 484140 11132
rect 484112 11008 484140 11104
rect 484918 11008 484946 11172
rect 485240 11132 485268 11200
rect 485194 11104 485268 11132
rect 485332 11132 485360 11308
rect 485458 11200 485514 11308
rect 485608 11308 485786 11336
rect 485608 11132 485636 11308
rect 485730 11200 485786 11308
rect 486002 11336 486058 12000
rect 486142 11336 486148 11348
rect 486002 11308 486148 11336
rect 486002 11200 486058 11308
rect 486142 11296 486148 11308
rect 486200 11296 486206 11348
rect 486274 11268 486330 12000
rect 486546 11336 486602 12000
rect 486694 11336 486700 11348
rect 486546 11308 486700 11336
rect 486418 11268 486424 11280
rect 486274 11240 486424 11268
rect 486274 11200 486330 11240
rect 486418 11228 486424 11240
rect 486476 11228 486482 11280
rect 486546 11200 486602 11308
rect 486694 11296 486700 11308
rect 486752 11296 486758 11348
rect 486818 11336 486874 12000
rect 486970 11336 486976 11348
rect 486818 11308 486976 11336
rect 486818 11200 486874 11308
rect 486970 11296 486976 11308
rect 487028 11296 487034 11348
rect 487090 11268 487146 12000
rect 487246 11268 487252 11280
rect 487090 11240 487252 11268
rect 487090 11200 487146 11240
rect 487246 11228 487252 11240
rect 487304 11228 487310 11280
rect 487362 11268 487418 12000
rect 487522 11268 487528 11280
rect 487362 11240 487528 11268
rect 487362 11200 487418 11240
rect 487522 11228 487528 11240
rect 487580 11228 487586 11280
rect 487634 11268 487690 12000
rect 487798 11268 487804 11280
rect 487634 11240 487804 11268
rect 487634 11200 487690 11240
rect 487798 11228 487804 11240
rect 487856 11228 487862 11280
rect 487906 11268 487962 12000
rect 488074 11268 488080 11280
rect 487906 11240 488080 11268
rect 487906 11200 487962 11240
rect 488074 11228 488080 11240
rect 488132 11228 488138 11280
rect 488178 11268 488234 12000
rect 488450 11336 488506 12000
rect 488534 11336 488540 11348
rect 488450 11308 488540 11336
rect 488350 11268 488356 11280
rect 488178 11240 488356 11268
rect 488178 11200 488234 11240
rect 488350 11228 488356 11240
rect 488408 11228 488414 11280
rect 488450 11200 488506 11308
rect 488534 11296 488540 11308
rect 488592 11296 488598 11348
rect 488722 11336 488778 12000
rect 488810 11336 488816 11348
rect 488722 11308 488816 11336
rect 488722 11200 488778 11308
rect 488810 11296 488816 11308
rect 488868 11296 488874 11348
rect 485774 11132 485780 11144
rect 485332 11104 485498 11132
rect 485608 11104 485780 11132
rect 484112 10968 484124 11008
rect 484118 10956 484124 10968
rect 484176 10956 484182 11008
rect 484918 10968 484952 11008
rect 484946 10956 484952 10968
rect 485004 10956 485010 11008
rect 485038 10956 485044 11008
rect 485096 10996 485102 11008
rect 485194 10996 485222 11104
rect 485096 10968 485222 10996
rect 485096 10956 485102 10968
rect 483072 10900 483152 10928
rect 483072 10888 483078 10900
rect 484302 10888 484308 10940
rect 484360 10928 484366 10940
rect 485470 10928 485498 11104
rect 485774 11092 485780 11104
rect 485832 11092 485838 11144
rect 484360 10900 485498 10928
rect 484360 10888 484366 10900
rect 380032 10560 383056 10588
rect 380032 10548 380038 10560
rect 297726 10480 297732 10532
rect 297784 10520 297790 10532
rect 370130 10520 370136 10532
rect 297784 10492 370136 10520
rect 297784 10480 297790 10492
rect 370130 10480 370136 10492
rect 370188 10480 370194 10532
rect 257028 10424 260972 10452
rect 257028 10412 257034 10424
rect 302418 10412 302424 10464
rect 302476 10452 302482 10464
rect 371050 10452 371056 10464
rect 302476 10424 371056 10452
rect 302476 10412 302482 10424
rect 371050 10412 371056 10424
rect 371108 10412 371114 10464
rect 378134 10412 378140 10464
rect 378192 10452 378198 10464
rect 385218 10452 385224 10464
rect 378192 10424 385224 10452
rect 378192 10412 378198 10424
rect 385218 10412 385224 10424
rect 385276 10412 385282 10464
rect 145742 10344 145748 10396
rect 145800 10384 145806 10396
rect 205818 10384 205824 10396
rect 145800 10356 205824 10384
rect 145800 10344 145806 10356
rect 205818 10344 205824 10356
rect 205876 10344 205882 10396
rect 210326 10344 210332 10396
rect 210384 10384 210390 10396
rect 220078 10384 220084 10396
rect 210384 10356 220084 10384
rect 210384 10344 210390 10356
rect 220078 10344 220084 10356
rect 220136 10344 220142 10396
rect 220170 10344 220176 10396
rect 220228 10384 220234 10396
rect 230842 10384 230848 10396
rect 220228 10356 230848 10384
rect 220228 10344 220234 10356
rect 230842 10344 230848 10356
rect 230900 10344 230906 10396
rect 239030 10344 239036 10396
rect 239088 10384 239094 10396
rect 249058 10384 249064 10396
rect 239088 10356 249064 10384
rect 239088 10344 239094 10356
rect 249058 10344 249064 10356
rect 249116 10344 249122 10396
rect 307478 10344 307484 10396
rect 307536 10384 307542 10396
rect 372154 10384 372160 10396
rect 307536 10356 372160 10384
rect 307536 10344 307542 10356
rect 372154 10344 372160 10356
rect 372212 10344 372218 10396
rect 376846 10344 376852 10396
rect 376904 10384 376910 10396
rect 383194 10384 383200 10396
rect 376904 10356 383200 10384
rect 376904 10344 376910 10356
rect 383194 10344 383200 10356
rect 383252 10344 383258 10396
rect 56594 10276 56600 10328
rect 56652 10316 56658 10328
rect 145834 10316 145840 10328
rect 56652 10288 145840 10316
rect 56652 10276 56658 10288
rect 145834 10276 145840 10288
rect 145892 10276 145898 10328
rect 149698 10276 149704 10328
rect 149756 10316 149762 10328
rect 205634 10316 205640 10328
rect 149756 10288 205640 10316
rect 149756 10276 149762 10288
rect 205634 10276 205640 10288
rect 205692 10276 205698 10328
rect 210142 10276 210148 10328
rect 210200 10316 210206 10328
rect 212350 10316 212356 10328
rect 210200 10288 212356 10316
rect 210200 10276 210206 10288
rect 212350 10276 212356 10288
rect 212408 10276 212414 10328
rect 212442 10276 212448 10328
rect 212500 10316 212506 10328
rect 217594 10316 217600 10328
rect 212500 10288 217600 10316
rect 212500 10276 212506 10288
rect 217594 10276 217600 10288
rect 217652 10276 217658 10328
rect 217870 10276 217876 10328
rect 217928 10316 217934 10328
rect 220906 10316 220912 10328
rect 217928 10288 220912 10316
rect 217928 10276 217934 10288
rect 220906 10276 220912 10288
rect 220964 10276 220970 10328
rect 251910 10276 251916 10328
rect 251968 10316 251974 10328
rect 258626 10316 258632 10328
rect 251968 10288 258632 10316
rect 251968 10276 251974 10288
rect 258626 10276 258632 10288
rect 258684 10276 258690 10328
rect 312446 10276 312452 10328
rect 312504 10316 312510 10328
rect 373258 10316 373264 10328
rect 312504 10288 373264 10316
rect 312504 10276 312510 10288
rect 373258 10276 373264 10288
rect 373316 10276 373322 10328
rect 382182 10276 382188 10328
rect 382240 10316 382246 10328
rect 385954 10316 385960 10328
rect 382240 10288 385960 10316
rect 382240 10276 382246 10288
rect 385954 10276 385960 10288
rect 386012 10276 386018 10328
rect 95142 10208 95148 10260
rect 95200 10248 95206 10260
rect 176654 10248 176660 10260
rect 95200 10220 176660 10248
rect 95200 10208 95206 10220
rect 176654 10208 176660 10220
rect 176712 10208 176718 10260
rect 187878 10208 187884 10260
rect 187936 10248 187942 10260
rect 198458 10248 198464 10260
rect 187936 10220 198464 10248
rect 187936 10208 187942 10220
rect 198458 10208 198464 10220
rect 198516 10208 198522 10260
rect 198642 10208 198648 10260
rect 198700 10248 198706 10260
rect 205358 10248 205364 10260
rect 198700 10220 205364 10248
rect 198700 10208 198706 10220
rect 205358 10208 205364 10220
rect 205416 10208 205422 10260
rect 206002 10208 206008 10260
rect 206060 10248 206066 10260
rect 213914 10248 213920 10260
rect 206060 10220 213920 10248
rect 206060 10208 206066 10220
rect 213914 10208 213920 10220
rect 213972 10208 213978 10260
rect 214098 10208 214104 10260
rect 214156 10248 214162 10260
rect 316310 10248 316316 10260
rect 214156 10220 316316 10248
rect 214156 10208 214162 10220
rect 316310 10208 316316 10220
rect 316368 10208 316374 10260
rect 317506 10208 317512 10260
rect 317564 10248 317570 10260
rect 374362 10248 374368 10260
rect 317564 10220 374368 10248
rect 317564 10208 317570 10220
rect 374362 10208 374368 10220
rect 374420 10208 374426 10260
rect 382918 10208 382924 10260
rect 382976 10248 382982 10260
rect 386506 10248 386512 10260
rect 382976 10220 386512 10248
rect 382976 10208 382982 10220
rect 386506 10208 386512 10220
rect 386564 10208 386570 10260
rect 173066 10140 173072 10192
rect 173124 10180 173130 10192
rect 225782 10180 225788 10192
rect 173124 10152 225788 10180
rect 173124 10140 173130 10152
rect 225782 10140 225788 10152
rect 225840 10140 225846 10192
rect 322474 10140 322480 10192
rect 322532 10180 322538 10192
rect 375466 10180 375472 10192
rect 322532 10152 375472 10180
rect 322532 10140 322538 10152
rect 375466 10140 375472 10152
rect 375524 10140 375530 10192
rect 112806 10072 112812 10124
rect 112864 10112 112870 10124
rect 175366 10112 175372 10124
rect 112864 10084 175372 10112
rect 112864 10072 112870 10084
rect 175366 10072 175372 10084
rect 175424 10072 175430 10124
rect 176286 10072 176292 10124
rect 176344 10112 176350 10124
rect 227346 10112 227352 10124
rect 176344 10084 227352 10112
rect 176344 10072 176350 10084
rect 227346 10072 227352 10084
rect 227404 10072 227410 10124
rect 332502 10072 332508 10124
rect 332560 10112 332566 10124
rect 377582 10112 377588 10124
rect 332560 10084 377588 10112
rect 332560 10072 332566 10084
rect 377582 10072 377588 10084
rect 377640 10072 377646 10124
rect 93762 10004 93768 10056
rect 93820 10044 93826 10056
rect 186222 10044 186228 10056
rect 93820 10016 186228 10044
rect 93820 10004 93826 10016
rect 186222 10004 186228 10016
rect 186280 10004 186286 10056
rect 186314 10004 186320 10056
rect 186372 10044 186378 10056
rect 205634 10044 205640 10056
rect 186372 10016 205640 10044
rect 186372 10004 186378 10016
rect 205634 10004 205640 10016
rect 205692 10004 205698 10056
rect 206738 10044 206744 10056
rect 205744 10016 206744 10044
rect 92106 9936 92112 9988
rect 92164 9976 92170 9988
rect 195054 9976 195060 9988
rect 92164 9948 195060 9976
rect 92164 9936 92170 9948
rect 195054 9936 195060 9948
rect 195112 9936 195118 9988
rect 195146 9936 195152 9988
rect 195204 9976 195210 9988
rect 198366 9976 198372 9988
rect 195204 9948 198372 9976
rect 195204 9936 195210 9948
rect 198366 9936 198372 9948
rect 198424 9936 198430 9988
rect 198550 9936 198556 9988
rect 198608 9976 198614 9988
rect 202874 9976 202880 9988
rect 198608 9948 202880 9976
rect 198608 9936 198614 9948
rect 202874 9936 202880 9948
rect 202932 9936 202938 9988
rect 203610 9936 203616 9988
rect 203668 9976 203674 9988
rect 205744 9976 205772 10016
rect 206738 10004 206744 10016
rect 206796 10004 206802 10056
rect 206830 10004 206836 10056
rect 206888 10044 206894 10056
rect 217226 10044 217232 10056
rect 206888 10016 217232 10044
rect 206888 10004 206894 10016
rect 217226 10004 217232 10016
rect 217284 10004 217290 10056
rect 219986 10004 219992 10056
rect 220044 10044 220050 10056
rect 321278 10044 321284 10056
rect 220044 10016 321284 10044
rect 220044 10004 220050 10016
rect 321278 10004 321284 10016
rect 321336 10004 321342 10056
rect 337470 10004 337476 10056
rect 337528 10044 337534 10056
rect 378686 10044 378692 10056
rect 337528 10016 378692 10044
rect 337528 10004 337534 10016
rect 378686 10004 378692 10016
rect 378744 10004 378750 10056
rect 203668 9948 205772 9976
rect 203668 9936 203674 9948
rect 205818 9936 205824 9988
rect 205876 9976 205882 9988
rect 214006 9976 214012 9988
rect 205876 9948 214012 9976
rect 205876 9936 205882 9948
rect 214006 9936 214012 9948
rect 214064 9936 214070 9988
rect 218422 9936 218428 9988
rect 218480 9976 218486 9988
rect 326338 9976 326344 9988
rect 218480 9948 326344 9976
rect 218480 9936 218486 9948
rect 326338 9936 326344 9948
rect 326396 9936 326402 9988
rect 340138 9936 340144 9988
rect 340196 9976 340202 9988
rect 379422 9976 379428 9988
rect 340196 9948 379428 9976
rect 340196 9936 340202 9948
rect 379422 9936 379428 9948
rect 379480 9936 379486 9988
rect 178034 9868 178040 9920
rect 178092 9908 178098 9920
rect 211246 9908 211252 9920
rect 178092 9880 211252 9908
rect 178092 9868 178098 9880
rect 211246 9868 211252 9880
rect 211304 9868 211310 9920
rect 213822 9868 213828 9920
rect 213880 9908 213886 9920
rect 229646 9908 229652 9920
rect 213880 9880 229652 9908
rect 213880 9868 213886 9880
rect 229646 9868 229652 9880
rect 229704 9868 229710 9920
rect 262398 9868 262404 9920
rect 262456 9908 262462 9920
rect 368566 9908 368572 9920
rect 262456 9880 368572 9908
rect 262456 9868 262462 9880
rect 368566 9868 368572 9880
rect 368624 9868 368630 9920
rect 1104 9818 528816 9840
rect 1104 9766 67574 9818
rect 67626 9766 67638 9818
rect 67690 9766 67702 9818
rect 67754 9766 67766 9818
rect 67818 9766 67830 9818
rect 67882 9766 199502 9818
rect 199554 9766 199566 9818
rect 199618 9766 199630 9818
rect 199682 9766 199694 9818
rect 199746 9766 199758 9818
rect 199810 9766 331430 9818
rect 331482 9766 331494 9818
rect 331546 9766 331558 9818
rect 331610 9766 331622 9818
rect 331674 9766 331686 9818
rect 331738 9766 463358 9818
rect 463410 9766 463422 9818
rect 463474 9766 463486 9818
rect 463538 9766 463550 9818
rect 463602 9766 463614 9818
rect 463666 9766 528816 9818
rect 1104 9744 528816 9766
rect 127802 9664 127808 9716
rect 127860 9704 127866 9716
rect 186590 9704 186596 9716
rect 127860 9676 186596 9704
rect 127860 9664 127866 9676
rect 186590 9664 186596 9676
rect 186648 9664 186654 9716
rect 198458 9664 198464 9716
rect 198516 9704 198522 9716
rect 200850 9704 200856 9716
rect 198516 9676 200856 9704
rect 198516 9664 198522 9676
rect 200850 9664 200856 9676
rect 200908 9664 200914 9716
rect 200942 9664 200948 9716
rect 201000 9704 201006 9716
rect 205266 9704 205272 9716
rect 201000 9676 205272 9704
rect 201000 9664 201006 9676
rect 205266 9664 205272 9676
rect 205324 9664 205330 9716
rect 205542 9664 205548 9716
rect 205600 9704 205606 9716
rect 306374 9704 306380 9716
rect 205600 9676 306380 9704
rect 205600 9664 205606 9676
rect 306374 9664 306380 9676
rect 306432 9664 306438 9716
rect 382090 9704 382096 9716
rect 352760 9676 382096 9704
rect 123386 9596 123392 9648
rect 123444 9636 123450 9648
rect 123444 9608 218100 9636
rect 123444 9596 123450 9608
rect 166966 9540 167316 9568
rect 82446 9460 82452 9512
rect 82504 9500 82510 9512
rect 166966 9500 166994 9540
rect 82504 9472 166994 9500
rect 82504 9460 82510 9472
rect 74718 9392 74724 9444
rect 74776 9432 74782 9444
rect 167086 9432 167092 9444
rect 74776 9404 167092 9432
rect 74776 9392 74782 9404
rect 167086 9392 167092 9404
rect 167144 9392 167150 9444
rect 167288 9432 167316 9540
rect 171778 9528 171784 9580
rect 171836 9568 171842 9580
rect 178034 9568 178040 9580
rect 171836 9540 178040 9568
rect 171836 9528 171842 9540
rect 178034 9528 178040 9540
rect 178092 9528 178098 9580
rect 183281 9571 183339 9577
rect 183281 9537 183293 9571
rect 183327 9568 183339 9571
rect 184382 9568 184388 9580
rect 183327 9540 184388 9568
rect 183327 9537 183339 9540
rect 183281 9531 183339 9537
rect 184382 9528 184388 9540
rect 184440 9528 184446 9580
rect 190825 9571 190883 9577
rect 190825 9537 190837 9571
rect 190871 9568 190883 9571
rect 191466 9568 191472 9580
rect 190871 9540 191472 9568
rect 190871 9537 190883 9540
rect 190825 9531 190883 9537
rect 191466 9528 191472 9540
rect 191524 9528 191530 9580
rect 195241 9571 195299 9577
rect 195241 9537 195253 9571
rect 195287 9568 195299 9571
rect 195882 9568 195888 9580
rect 195287 9540 195888 9568
rect 195287 9537 195299 9540
rect 195241 9531 195299 9537
rect 195882 9528 195888 9540
rect 195940 9528 195946 9580
rect 198369 9571 198427 9577
rect 198369 9537 198381 9571
rect 198415 9568 198427 9571
rect 202969 9571 203027 9577
rect 198415 9540 199056 9568
rect 198415 9537 198427 9540
rect 198369 9531 198427 9537
rect 167362 9460 167368 9512
rect 167420 9500 167426 9512
rect 182729 9503 182787 9509
rect 182729 9500 182741 9503
rect 167420 9472 182741 9500
rect 167420 9460 167426 9472
rect 182729 9469 182741 9472
rect 182775 9469 182787 9503
rect 182729 9463 182787 9469
rect 190273 9503 190331 9509
rect 190273 9469 190285 9503
rect 190319 9469 190331 9503
rect 190273 9463 190331 9469
rect 190288 9432 190316 9463
rect 194686 9460 194692 9512
rect 194744 9460 194750 9512
rect 197817 9503 197875 9509
rect 197817 9500 197829 9503
rect 195946 9472 197829 9500
rect 195946 9432 195974 9472
rect 197817 9469 197829 9472
rect 197863 9469 197875 9503
rect 197817 9463 197875 9469
rect 167288 9404 190316 9432
rect 190426 9404 195974 9432
rect 90174 9324 90180 9376
rect 90232 9364 90238 9376
rect 190426 9364 190454 9404
rect 90232 9336 190454 9364
rect 90232 9324 90238 9336
rect 191466 9324 191472 9376
rect 191524 9324 191530 9376
rect 199028 9373 199056 9540
rect 202969 9537 202981 9571
rect 203015 9568 203027 9571
rect 203610 9568 203616 9580
rect 203015 9540 203616 9568
rect 203015 9537 203027 9540
rect 202969 9531 203027 9537
rect 203610 9528 203616 9540
rect 203668 9528 203674 9580
rect 205729 9571 205787 9577
rect 205729 9537 205741 9571
rect 205775 9568 205787 9571
rect 206278 9568 206284 9580
rect 205775 9540 206284 9568
rect 205775 9537 205787 9540
rect 205729 9531 205787 9537
rect 206278 9528 206284 9540
rect 206336 9528 206342 9580
rect 210513 9571 210571 9577
rect 210513 9537 210525 9571
rect 210559 9568 210571 9571
rect 211062 9568 211068 9580
rect 210559 9540 211068 9568
rect 210559 9537 210571 9540
rect 210513 9531 210571 9537
rect 211062 9528 211068 9540
rect 211120 9528 211126 9580
rect 213273 9571 213331 9577
rect 213273 9537 213285 9571
rect 213319 9568 213331 9571
rect 213822 9568 213828 9580
rect 213319 9540 213828 9568
rect 213319 9537 213331 9540
rect 213273 9531 213331 9537
rect 213822 9528 213828 9540
rect 213880 9528 213886 9580
rect 202414 9460 202420 9512
rect 202472 9460 202478 9512
rect 205450 9460 205456 9512
rect 205508 9460 205514 9512
rect 210234 9460 210240 9512
rect 210292 9460 210298 9512
rect 212534 9460 212540 9512
rect 212592 9500 212598 9512
rect 212997 9503 213055 9509
rect 212997 9500 213009 9503
rect 212592 9472 213009 9500
rect 212592 9460 212598 9472
rect 212997 9469 213009 9472
rect 213043 9469 213055 9503
rect 212997 9463 213055 9469
rect 217962 9460 217968 9512
rect 218020 9460 218026 9512
rect 218072 9500 218100 9608
rect 218790 9596 218796 9648
rect 218848 9596 218854 9648
rect 221366 9636 221372 9648
rect 220832 9608 221372 9636
rect 218241 9571 218299 9577
rect 218241 9537 218253 9571
rect 218287 9568 218299 9571
rect 218808 9568 218836 9596
rect 220832 9577 220860 9608
rect 221366 9596 221372 9608
rect 221424 9596 221430 9648
rect 225601 9639 225659 9645
rect 225601 9605 225613 9639
rect 225647 9636 225659 9639
rect 248598 9636 248604 9648
rect 225647 9608 248604 9636
rect 225647 9605 225659 9608
rect 225601 9599 225659 9605
rect 218287 9540 218836 9568
rect 220817 9571 220875 9577
rect 218287 9537 218299 9540
rect 218241 9531 218299 9537
rect 220817 9537 220829 9571
rect 220863 9537 220875 9571
rect 220817 9531 220875 9537
rect 224957 9571 225015 9577
rect 224957 9537 224969 9571
rect 225003 9568 225015 9571
rect 225616 9568 225644 9599
rect 248598 9596 248604 9608
rect 248656 9596 248662 9648
rect 340138 9636 340144 9648
rect 339512 9608 340144 9636
rect 225003 9540 225644 9568
rect 228545 9571 228603 9577
rect 225003 9537 225015 9540
rect 224957 9531 225015 9537
rect 228545 9537 228557 9571
rect 228591 9568 228603 9571
rect 229094 9568 229100 9580
rect 228591 9540 229100 9568
rect 228591 9537 228603 9540
rect 228545 9531 228603 9537
rect 229094 9528 229100 9540
rect 229152 9528 229158 9580
rect 232501 9571 232559 9577
rect 232501 9537 232513 9571
rect 232547 9568 232559 9571
rect 232547 9540 233372 9568
rect 232547 9537 232559 9540
rect 232501 9531 232559 9537
rect 220354 9500 220360 9512
rect 218072 9472 220360 9500
rect 220354 9460 220360 9472
rect 220412 9460 220418 9512
rect 220538 9460 220544 9512
rect 220596 9460 220602 9512
rect 224678 9460 224684 9512
rect 224736 9460 224742 9512
rect 228266 9460 228272 9512
rect 228324 9460 228330 9512
rect 232038 9460 232044 9512
rect 232096 9500 232102 9512
rect 232225 9503 232283 9509
rect 232225 9500 232237 9503
rect 232096 9472 232237 9500
rect 232096 9460 232102 9472
rect 232225 9469 232237 9472
rect 232271 9469 232283 9503
rect 232225 9463 232283 9469
rect 200758 9392 200764 9444
rect 200816 9432 200822 9444
rect 232314 9432 232320 9444
rect 200816 9404 232320 9432
rect 200816 9392 200822 9404
rect 232314 9392 232320 9404
rect 232372 9392 232378 9444
rect 233344 9441 233372 9540
rect 234430 9528 234436 9580
rect 234488 9568 234494 9580
rect 236273 9571 236331 9577
rect 234488 9540 236224 9568
rect 234488 9528 234494 9540
rect 235994 9460 236000 9512
rect 236052 9460 236058 9512
rect 233329 9435 233387 9441
rect 233329 9401 233341 9435
rect 233375 9432 233387 9435
rect 236196 9432 236224 9540
rect 236273 9537 236285 9571
rect 236319 9568 236331 9571
rect 236319 9540 236868 9568
rect 236319 9537 236331 9540
rect 236273 9531 236331 9537
rect 236840 9512 236868 9540
rect 239950 9528 239956 9580
rect 240008 9528 240014 9580
rect 243998 9528 244004 9580
rect 244056 9528 244062 9580
rect 339512 9577 339540 9608
rect 340138 9596 340144 9608
rect 340196 9596 340202 9648
rect 342714 9636 342720 9648
rect 342088 9608 342720 9636
rect 342088 9577 342116 9608
rect 342714 9596 342720 9608
rect 342772 9596 342778 9648
rect 352760 9645 352788 9676
rect 382090 9664 382096 9676
rect 382148 9664 382154 9716
rect 345293 9639 345351 9645
rect 345293 9636 345305 9639
rect 344986 9608 345305 9636
rect 339497 9571 339555 9577
rect 339497 9537 339509 9571
rect 339543 9537 339555 9571
rect 339497 9531 339555 9537
rect 342073 9571 342131 9577
rect 342073 9537 342085 9571
rect 342119 9537 342131 9571
rect 342073 9531 342131 9537
rect 344649 9571 344707 9577
rect 344649 9537 344661 9571
rect 344695 9568 344707 9571
rect 344986 9568 345014 9608
rect 345293 9605 345305 9608
rect 345339 9636 345351 9639
rect 352745 9639 352803 9645
rect 345339 9608 352144 9636
rect 345339 9605 345351 9608
rect 345293 9599 345351 9605
rect 344695 9540 345014 9568
rect 344695 9537 344707 9540
rect 344649 9531 344707 9537
rect 346762 9528 346768 9580
rect 346820 9528 346826 9580
rect 347041 9571 347099 9577
rect 347041 9537 347053 9571
rect 347087 9568 347099 9571
rect 347590 9568 347596 9580
rect 347087 9540 347596 9568
rect 347087 9537 347099 9540
rect 347041 9531 347099 9537
rect 347590 9528 347596 9540
rect 347648 9528 347654 9580
rect 349617 9571 349675 9577
rect 349617 9537 349629 9571
rect 349663 9568 349675 9571
rect 350074 9568 350080 9580
rect 349663 9540 350080 9568
rect 349663 9537 349675 9540
rect 349617 9531 349675 9537
rect 350074 9528 350080 9540
rect 350132 9528 350138 9580
rect 236822 9460 236828 9512
rect 236880 9460 236886 9512
rect 239674 9460 239680 9512
rect 239732 9460 239738 9512
rect 243722 9460 243728 9512
rect 243780 9460 243786 9512
rect 338942 9460 338948 9512
rect 339000 9460 339006 9512
rect 341521 9503 341579 9509
rect 341521 9469 341533 9503
rect 341567 9469 341579 9503
rect 341521 9463 341579 9469
rect 341536 9432 341564 9463
rect 344094 9460 344100 9512
rect 344152 9460 344158 9512
rect 349338 9460 349344 9512
rect 349396 9460 349402 9512
rect 351914 9460 351920 9512
rect 351972 9460 351978 9512
rect 352116 9500 352144 9608
rect 352745 9605 352757 9639
rect 352791 9605 352803 9639
rect 352745 9599 352803 9605
rect 352193 9571 352251 9577
rect 352193 9537 352205 9571
rect 352239 9568 352251 9571
rect 352760 9568 352788 9599
rect 354398 9596 354404 9648
rect 354456 9636 354462 9648
rect 354493 9639 354551 9645
rect 354493 9636 354505 9639
rect 354456 9608 354505 9636
rect 354456 9596 354462 9608
rect 354493 9605 354505 9608
rect 354539 9605 354551 9639
rect 354493 9599 354551 9605
rect 354582 9596 354588 9648
rect 354640 9636 354646 9648
rect 366085 9639 366143 9645
rect 366085 9636 366097 9639
rect 354640 9608 366097 9636
rect 354640 9596 354646 9608
rect 366085 9605 366097 9608
rect 366131 9605 366143 9639
rect 367278 9636 367284 9648
rect 366085 9599 366143 9605
rect 366376 9608 367284 9636
rect 352239 9540 352788 9568
rect 354769 9571 354827 9577
rect 352239 9537 352251 9540
rect 352193 9531 352251 9537
rect 354769 9537 354781 9571
rect 354815 9568 354827 9571
rect 355318 9568 355324 9580
rect 354815 9540 355324 9568
rect 354815 9537 354827 9540
rect 354769 9531 354827 9537
rect 355318 9528 355324 9540
rect 355376 9528 355382 9580
rect 357345 9571 357403 9577
rect 357345 9537 357357 9571
rect 357391 9568 357403 9571
rect 357894 9568 357900 9580
rect 357391 9540 357900 9568
rect 357391 9537 357403 9540
rect 357345 9531 357403 9537
rect 357894 9528 357900 9540
rect 357952 9528 357958 9580
rect 358630 9528 358636 9580
rect 358688 9528 358694 9580
rect 366376 9577 366404 9608
rect 367278 9596 367284 9608
rect 367336 9596 367342 9648
rect 368566 9596 368572 9648
rect 368624 9596 368630 9648
rect 379238 9636 379244 9648
rect 370884 9608 379244 9636
rect 358909 9571 358967 9577
rect 358909 9537 358921 9571
rect 358955 9568 358967 9571
rect 359553 9571 359611 9577
rect 359553 9568 359565 9571
rect 358955 9540 359565 9568
rect 358955 9537 358967 9540
rect 358909 9531 358967 9537
rect 359553 9537 359565 9540
rect 359599 9568 359611 9571
rect 361485 9571 361543 9577
rect 359599 9540 361344 9568
rect 359599 9537 359611 9540
rect 359553 9531 359611 9537
rect 352116 9472 354720 9500
rect 354582 9432 354588 9444
rect 233375 9404 234614 9432
rect 236196 9404 341564 9432
rect 341628 9404 354588 9432
rect 233375 9401 233387 9404
rect 233329 9395 233387 9401
rect 199013 9367 199071 9373
rect 199013 9333 199025 9367
rect 199059 9364 199071 9367
rect 199194 9364 199200 9376
rect 199059 9336 199200 9364
rect 199059 9333 199071 9336
rect 199013 9327 199071 9333
rect 199194 9324 199200 9336
rect 199252 9324 199258 9376
rect 229094 9324 229100 9376
rect 229152 9324 229158 9376
rect 234586 9364 234614 9404
rect 241514 9364 241520 9376
rect 234586 9336 241520 9364
rect 241514 9324 241520 9336
rect 241572 9324 241578 9376
rect 243998 9324 244004 9376
rect 244056 9364 244062 9376
rect 244553 9367 244611 9373
rect 244553 9364 244565 9367
rect 244056 9336 244565 9364
rect 244056 9324 244062 9336
rect 244553 9333 244565 9336
rect 244599 9364 244611 9367
rect 255682 9364 255688 9376
rect 244599 9336 255688 9364
rect 244599 9333 244611 9336
rect 244553 9327 244611 9333
rect 255682 9324 255688 9336
rect 255740 9324 255746 9376
rect 260190 9324 260196 9376
rect 260248 9364 260254 9376
rect 341628 9364 341656 9404
rect 354582 9392 354588 9404
rect 354640 9392 354646 9444
rect 354692 9432 354720 9472
rect 357066 9460 357072 9512
rect 357124 9460 357130 9512
rect 360194 9460 360200 9512
rect 360252 9500 360258 9512
rect 361209 9503 361267 9509
rect 361209 9500 361221 9503
rect 360252 9472 361221 9500
rect 360252 9460 360258 9472
rect 361209 9469 361221 9472
rect 361255 9469 361267 9503
rect 361209 9463 361267 9469
rect 361316 9432 361344 9540
rect 361485 9537 361497 9571
rect 361531 9568 361543 9571
rect 363969 9571 364027 9577
rect 361531 9540 362172 9568
rect 361531 9537 361543 9540
rect 361485 9531 361543 9537
rect 362144 9512 362172 9540
rect 363969 9537 363981 9571
rect 364015 9537 364027 9571
rect 363969 9531 364027 9537
rect 366361 9571 366419 9577
rect 366361 9537 366373 9571
rect 366407 9537 366419 9571
rect 366361 9531 366419 9537
rect 366468 9540 368796 9568
rect 362126 9460 362132 9512
rect 362184 9460 362190 9512
rect 363690 9460 363696 9512
rect 363748 9460 363754 9512
rect 363984 9500 364012 9531
rect 364705 9503 364763 9509
rect 364705 9500 364717 9503
rect 363984 9472 364717 9500
rect 364705 9469 364717 9472
rect 364751 9500 364763 9503
rect 366468 9500 366496 9540
rect 364751 9472 366496 9500
rect 368768 9500 368796 9540
rect 368842 9528 368848 9580
rect 368900 9528 368906 9580
rect 370884 9500 370912 9608
rect 379238 9596 379244 9608
rect 379296 9596 379302 9648
rect 382182 9636 382188 9648
rect 379486 9608 382188 9636
rect 371326 9528 371332 9580
rect 371384 9528 371390 9580
rect 373721 9571 373779 9577
rect 373721 9537 373733 9571
rect 373767 9568 373779 9571
rect 374270 9568 374276 9580
rect 373767 9540 374276 9568
rect 373767 9537 373779 9540
rect 373721 9531 373779 9537
rect 374270 9528 374276 9540
rect 374328 9528 374334 9580
rect 376205 9571 376263 9577
rect 374380 9540 376064 9568
rect 368768 9472 370912 9500
rect 364751 9469 364763 9472
rect 364705 9463 364763 9469
rect 371050 9460 371056 9512
rect 371108 9460 371114 9512
rect 372706 9460 372712 9512
rect 372764 9500 372770 9512
rect 373445 9503 373503 9509
rect 373445 9500 373457 9503
rect 372764 9472 373457 9500
rect 372764 9460 372770 9472
rect 373445 9469 373457 9472
rect 373491 9469 373503 9503
rect 373445 9463 373503 9469
rect 373534 9460 373540 9512
rect 373592 9500 373598 9512
rect 374380 9500 374408 9540
rect 373592 9472 374408 9500
rect 373592 9460 373598 9472
rect 375926 9460 375932 9512
rect 375984 9460 375990 9512
rect 376036 9500 376064 9540
rect 376205 9537 376217 9571
rect 376251 9568 376263 9571
rect 376754 9568 376760 9580
rect 376251 9540 376760 9568
rect 376251 9537 376263 9540
rect 376205 9531 376263 9537
rect 376754 9528 376760 9540
rect 376812 9528 376818 9580
rect 378597 9571 378655 9577
rect 376864 9540 378456 9568
rect 376864 9500 376892 9540
rect 376036 9472 376892 9500
rect 378318 9460 378324 9512
rect 378376 9460 378382 9512
rect 378428 9500 378456 9540
rect 378597 9537 378609 9571
rect 378643 9568 378655 9571
rect 379146 9568 379152 9580
rect 378643 9540 379152 9568
rect 378643 9537 378655 9540
rect 378597 9531 378655 9537
rect 379146 9528 379152 9540
rect 379204 9528 379210 9580
rect 379486 9568 379514 9608
rect 382182 9596 382188 9608
rect 382240 9596 382246 9648
rect 384025 9639 384083 9645
rect 384025 9605 384037 9639
rect 384071 9636 384083 9639
rect 388990 9636 388996 9648
rect 384071 9608 388996 9636
rect 384071 9605 384083 9608
rect 384025 9599 384083 9605
rect 379256 9540 379514 9568
rect 381081 9571 381139 9577
rect 379256 9500 379284 9540
rect 381081 9537 381093 9571
rect 381127 9568 381139 9571
rect 383473 9571 383531 9577
rect 381127 9540 381676 9568
rect 381127 9537 381139 9540
rect 381081 9531 381139 9537
rect 379974 9500 379980 9512
rect 378428 9472 379284 9500
rect 379486 9472 379980 9500
rect 373626 9432 373632 9444
rect 354692 9404 361252 9432
rect 361316 9404 373632 9432
rect 260248 9336 341656 9364
rect 260248 9324 260254 9336
rect 350074 9324 350080 9376
rect 350132 9324 350138 9376
rect 355318 9324 355324 9376
rect 355376 9324 355382 9376
rect 357894 9324 357900 9376
rect 357952 9324 357958 9376
rect 361224 9364 361252 9404
rect 373626 9392 373632 9404
rect 373684 9392 373690 9444
rect 373810 9392 373816 9444
rect 373868 9432 373874 9444
rect 379486 9432 379514 9472
rect 379974 9460 379980 9472
rect 380032 9460 380038 9512
rect 380802 9460 380808 9512
rect 380860 9460 380866 9512
rect 381648 9441 381676 9540
rect 383473 9537 383485 9571
rect 383519 9568 383531 9571
rect 384040 9568 384068 9599
rect 388990 9596 388996 9608
rect 389048 9596 389054 9648
rect 383519 9540 384068 9568
rect 383519 9537 383531 9540
rect 383473 9531 383531 9537
rect 383010 9460 383016 9512
rect 383068 9500 383074 9512
rect 383197 9503 383255 9509
rect 383197 9500 383209 9503
rect 383068 9472 383209 9500
rect 383068 9460 383074 9472
rect 383197 9469 383209 9472
rect 383243 9469 383255 9503
rect 383197 9463 383255 9469
rect 373868 9404 379514 9432
rect 381633 9435 381691 9441
rect 373868 9392 373874 9404
rect 381633 9401 381645 9435
rect 381679 9432 381691 9435
rect 385770 9432 385776 9444
rect 381679 9404 385776 9432
rect 381679 9401 381691 9404
rect 381633 9395 381691 9401
rect 385770 9392 385776 9404
rect 385828 9392 385834 9444
rect 367094 9364 367100 9376
rect 361224 9336 367100 9364
rect 367094 9324 367100 9336
rect 367152 9324 367158 9376
rect 367278 9324 367284 9376
rect 367336 9324 367342 9376
rect 368842 9324 368848 9376
rect 368900 9364 368906 9376
rect 369857 9367 369915 9373
rect 369857 9364 369869 9367
rect 368900 9336 369869 9364
rect 368900 9324 368906 9336
rect 369857 9333 369869 9336
rect 369903 9364 369915 9367
rect 373534 9364 373540 9376
rect 369903 9336 373540 9364
rect 369903 9333 369915 9336
rect 369857 9327 369915 9333
rect 373534 9324 373540 9336
rect 373592 9324 373598 9376
rect 374270 9324 374276 9376
rect 374328 9324 374334 9376
rect 376754 9324 376760 9376
rect 376812 9324 376818 9376
rect 379146 9324 379152 9376
rect 379204 9324 379210 9376
rect 379238 9324 379244 9376
rect 379296 9364 379302 9376
rect 384666 9364 384672 9376
rect 379296 9336 384672 9364
rect 379296 9324 379302 9336
rect 384666 9324 384672 9336
rect 384724 9324 384730 9376
rect 1104 9274 528816 9296
rect 1104 9222 66914 9274
rect 66966 9222 66978 9274
rect 67030 9222 67042 9274
rect 67094 9222 67106 9274
rect 67158 9222 67170 9274
rect 67222 9222 198842 9274
rect 198894 9222 198906 9274
rect 198958 9222 198970 9274
rect 199022 9222 199034 9274
rect 199086 9222 199098 9274
rect 199150 9222 330770 9274
rect 330822 9222 330834 9274
rect 330886 9222 330898 9274
rect 330950 9222 330962 9274
rect 331014 9222 331026 9274
rect 331078 9222 462698 9274
rect 462750 9222 462762 9274
rect 462814 9222 462826 9274
rect 462878 9222 462890 9274
rect 462942 9222 462954 9274
rect 463006 9222 528816 9274
rect 1104 9200 528816 9222
rect 87598 9120 87604 9172
rect 87656 9160 87662 9172
rect 194686 9160 194692 9172
rect 87656 9132 194692 9160
rect 87656 9120 87662 9132
rect 194686 9120 194692 9132
rect 194744 9120 194750 9172
rect 194962 9120 194968 9172
rect 195020 9160 195026 9172
rect 215386 9160 215392 9172
rect 195020 9132 215392 9160
rect 195020 9120 195026 9132
rect 215386 9120 215392 9132
rect 215444 9120 215450 9172
rect 232866 9120 232872 9172
rect 232924 9160 232930 9172
rect 338942 9160 338948 9172
rect 232924 9132 338948 9160
rect 232924 9120 232930 9132
rect 338942 9120 338948 9132
rect 339000 9120 339006 9172
rect 357434 9120 357440 9172
rect 357492 9160 357498 9172
rect 375926 9160 375932 9172
rect 357492 9132 375932 9160
rect 357492 9120 357498 9132
rect 375926 9120 375932 9132
rect 375984 9120 375990 9172
rect 376754 9120 376760 9172
rect 376812 9160 376818 9172
rect 387978 9160 387984 9172
rect 376812 9132 387984 9160
rect 376812 9120 376818 9132
rect 387978 9120 387984 9132
rect 388036 9120 388042 9172
rect 110782 9052 110788 9104
rect 110840 9092 110846 9104
rect 217962 9092 217968 9104
rect 110840 9064 217968 9092
rect 110840 9052 110846 9064
rect 217962 9052 217968 9064
rect 218020 9052 218026 9104
rect 229094 9052 229100 9104
rect 229152 9092 229158 9104
rect 250254 9092 250260 9104
rect 229152 9064 250260 9092
rect 229152 9052 229158 9064
rect 250254 9052 250260 9064
rect 250312 9052 250318 9104
rect 265342 9052 265348 9104
rect 265400 9092 265406 9104
rect 371050 9092 371056 9104
rect 265400 9064 371056 9092
rect 265400 9052 265406 9064
rect 371050 9052 371056 9064
rect 371108 9052 371114 9104
rect 374270 9052 374276 9104
rect 374328 9092 374334 9104
rect 385862 9092 385868 9104
rect 374328 9064 385868 9092
rect 374328 9052 374334 9064
rect 385862 9052 385868 9064
rect 385920 9052 385926 9104
rect 161446 8996 168696 9024
rect 152737 8959 152795 8965
rect 152737 8925 152749 8959
rect 152783 8956 152795 8959
rect 160465 8959 160523 8965
rect 152783 8928 153516 8956
rect 152783 8925 152795 8928
rect 152737 8919 152795 8925
rect 43806 8848 43812 8900
rect 43864 8888 43870 8900
rect 152185 8891 152243 8897
rect 152185 8888 152197 8891
rect 43864 8860 152197 8888
rect 43864 8848 43870 8860
rect 152185 8857 152197 8860
rect 152231 8857 152243 8891
rect 152185 8851 152243 8857
rect 153488 8829 153516 8928
rect 160465 8925 160477 8959
rect 160511 8956 160523 8959
rect 161017 8959 161075 8965
rect 161017 8956 161029 8959
rect 160511 8928 161029 8956
rect 160511 8925 160523 8928
rect 160465 8919 160523 8925
rect 161017 8925 161029 8928
rect 161063 8956 161075 8959
rect 161446 8956 161474 8996
rect 161063 8928 161474 8956
rect 168101 8959 168159 8965
rect 161063 8925 161075 8928
rect 161017 8919 161075 8925
rect 168101 8925 168113 8959
rect 168147 8925 168159 8959
rect 168668 8956 168696 8996
rect 168742 8984 168748 9036
rect 168800 9024 168806 9036
rect 168800 8996 176654 9024
rect 168800 8984 168806 8996
rect 171778 8956 171784 8968
rect 168668 8928 171784 8956
rect 168101 8919 168159 8925
rect 160094 8848 160100 8900
rect 160152 8848 160158 8900
rect 167546 8848 167552 8900
rect 167604 8848 167610 8900
rect 168116 8888 168144 8919
rect 171778 8916 171784 8928
rect 171836 8916 171842 8968
rect 172425 8959 172483 8965
rect 172425 8925 172437 8959
rect 172471 8956 172483 8959
rect 173066 8956 173072 8968
rect 172471 8928 173072 8956
rect 172471 8925 172483 8928
rect 172425 8919 172483 8925
rect 173066 8916 173072 8928
rect 173124 8916 173130 8968
rect 175645 8959 175703 8965
rect 175645 8925 175657 8959
rect 175691 8956 175703 8959
rect 176286 8956 176292 8968
rect 175691 8928 176292 8956
rect 175691 8925 175703 8928
rect 175645 8919 175703 8925
rect 176286 8916 176292 8928
rect 176344 8916 176350 8968
rect 168116 8860 168880 8888
rect 153473 8823 153531 8829
rect 153473 8789 153485 8823
rect 153519 8820 153531 8823
rect 168742 8820 168748 8832
rect 153519 8792 168748 8820
rect 153519 8789 153531 8792
rect 153473 8783 153531 8789
rect 168742 8780 168748 8792
rect 168800 8780 168806 8832
rect 168852 8820 168880 8860
rect 171226 8848 171232 8900
rect 171284 8888 171290 8900
rect 171873 8891 171931 8897
rect 171873 8888 171885 8891
rect 171284 8860 171885 8888
rect 171284 8848 171290 8860
rect 171873 8857 171885 8860
rect 171919 8857 171931 8891
rect 171873 8851 171931 8857
rect 175274 8848 175280 8900
rect 175332 8848 175338 8900
rect 168929 8823 168987 8829
rect 168929 8820 168941 8823
rect 168852 8792 168941 8820
rect 168929 8789 168941 8792
rect 168975 8820 168987 8823
rect 175458 8820 175464 8832
rect 168975 8792 175464 8820
rect 168975 8789 168987 8792
rect 168929 8783 168987 8789
rect 175458 8780 175464 8792
rect 175516 8780 175522 8832
rect 176626 8820 176654 8996
rect 176746 8984 176752 9036
rect 176804 9024 176810 9036
rect 239674 9024 239680 9036
rect 176804 8996 239680 9024
rect 176804 8984 176810 8996
rect 239674 8984 239680 8996
rect 239732 8984 239738 9036
rect 239950 8984 239956 9036
rect 240008 9024 240014 9036
rect 240137 9027 240195 9033
rect 240137 9024 240149 9027
rect 240008 8996 240149 9024
rect 240008 8984 240014 8996
rect 240137 8993 240149 8996
rect 240183 9024 240195 9027
rect 251174 9024 251180 9036
rect 240183 8996 251180 9024
rect 240183 8993 240195 8996
rect 240137 8987 240195 8993
rect 251174 8984 251180 8996
rect 251232 8984 251238 9036
rect 275646 8984 275652 9036
rect 275704 9024 275710 9036
rect 380802 9024 380808 9036
rect 275704 8996 380808 9024
rect 275704 8984 275710 8996
rect 380802 8984 380808 8996
rect 380860 8984 380866 9036
rect 179969 8959 180027 8965
rect 179969 8925 179981 8959
rect 180015 8956 180027 8959
rect 180521 8959 180579 8965
rect 180521 8956 180533 8959
rect 180015 8928 180533 8956
rect 180015 8925 180027 8928
rect 179969 8919 180027 8925
rect 180521 8925 180533 8928
rect 180567 8956 180579 8959
rect 187510 8956 187516 8968
rect 180567 8928 187516 8956
rect 180567 8925 180579 8928
rect 180521 8919 180579 8925
rect 187510 8916 187516 8928
rect 187568 8916 187574 8968
rect 187605 8959 187663 8965
rect 187605 8925 187617 8959
rect 187651 8925 187663 8959
rect 187605 8919 187663 8925
rect 179414 8848 179420 8900
rect 179472 8848 179478 8900
rect 186406 8848 186412 8900
rect 186464 8888 186470 8900
rect 187053 8891 187111 8897
rect 187053 8888 187065 8891
rect 186464 8860 187065 8888
rect 186464 8848 186470 8860
rect 187053 8857 187065 8860
rect 187099 8857 187111 8891
rect 187620 8888 187648 8919
rect 187694 8916 187700 8968
rect 187752 8956 187758 8968
rect 229186 8956 229192 8968
rect 187752 8928 229192 8956
rect 187752 8916 187758 8928
rect 229186 8916 229192 8928
rect 229244 8916 229250 8968
rect 236822 8916 236828 8968
rect 236880 8956 236886 8968
rect 254026 8956 254032 8968
rect 236880 8928 254032 8956
rect 236880 8916 236886 8928
rect 254026 8916 254032 8928
rect 254084 8916 254090 8968
rect 321278 8916 321284 8968
rect 321336 8916 321342 8968
rect 321833 8959 321891 8965
rect 321833 8925 321845 8959
rect 321879 8956 321891 8959
rect 322474 8956 322480 8968
rect 321879 8928 322480 8956
rect 321879 8925 321891 8928
rect 321833 8919 321891 8925
rect 322474 8916 322480 8928
rect 322532 8916 322538 8968
rect 326338 8916 326344 8968
rect 326396 8916 326402 8968
rect 326893 8959 326951 8965
rect 326893 8925 326905 8959
rect 326939 8956 326951 8959
rect 327534 8956 327540 8968
rect 326939 8928 327540 8956
rect 326939 8925 326951 8928
rect 326893 8919 326951 8925
rect 327534 8916 327540 8928
rect 327592 8916 327598 8968
rect 331861 8959 331919 8965
rect 331861 8925 331873 8959
rect 331907 8956 331919 8959
rect 332502 8956 332508 8968
rect 331907 8928 332508 8956
rect 331907 8925 331919 8928
rect 331861 8919 331919 8925
rect 332502 8916 332508 8928
rect 332560 8916 332566 8968
rect 336274 8916 336280 8968
rect 336332 8916 336338 8968
rect 336829 8959 336887 8965
rect 336829 8925 336841 8959
rect 336875 8956 336887 8959
rect 337470 8956 337476 8968
rect 336875 8928 337476 8956
rect 336875 8925 336887 8928
rect 336829 8919 336887 8925
rect 337470 8916 337476 8928
rect 337528 8916 337534 8968
rect 355318 8916 355324 8968
rect 355376 8956 355382 8968
rect 364150 8956 364156 8968
rect 355376 8928 364156 8956
rect 355376 8916 355382 8928
rect 364150 8916 364156 8928
rect 364208 8916 364214 8968
rect 365806 8916 365812 8968
rect 365864 8956 365870 8968
rect 378318 8956 378324 8968
rect 365864 8928 378324 8956
rect 365864 8916 365870 8928
rect 378318 8916 378324 8928
rect 378376 8916 378382 8968
rect 187620 8860 187740 8888
rect 187053 8851 187111 8857
rect 187510 8820 187516 8832
rect 176626 8792 187516 8820
rect 187510 8780 187516 8792
rect 187568 8780 187574 8832
rect 187712 8820 187740 8860
rect 187786 8848 187792 8900
rect 187844 8888 187850 8900
rect 212442 8888 212448 8900
rect 187844 8860 212448 8888
rect 187844 8848 187850 8860
rect 212442 8848 212448 8860
rect 212500 8848 212506 8900
rect 224126 8848 224132 8900
rect 224184 8888 224190 8900
rect 331309 8891 331367 8897
rect 331309 8888 331321 8891
rect 224184 8860 316034 8888
rect 224184 8848 224190 8860
rect 188249 8823 188307 8829
rect 188249 8820 188261 8823
rect 187712 8792 188261 8820
rect 188249 8789 188261 8792
rect 188295 8820 188307 8823
rect 200758 8820 200764 8832
rect 188295 8792 200764 8820
rect 188295 8789 188307 8792
rect 188249 8783 188307 8789
rect 200758 8780 200764 8792
rect 200816 8780 200822 8832
rect 316006 8820 316034 8860
rect 321388 8860 325694 8888
rect 321388 8820 321416 8860
rect 316006 8792 321416 8820
rect 325666 8820 325694 8860
rect 326724 8860 331321 8888
rect 326724 8820 326752 8860
rect 331309 8857 331321 8860
rect 331355 8857 331367 8891
rect 331309 8851 331367 8857
rect 362126 8848 362132 8900
rect 362184 8888 362190 8900
rect 383562 8888 383568 8900
rect 362184 8860 383568 8888
rect 362184 8848 362190 8860
rect 383562 8848 383568 8860
rect 383620 8848 383626 8900
rect 325666 8792 326752 8820
rect 327534 8780 327540 8832
rect 327592 8780 327598 8832
rect 371326 8780 371332 8832
rect 371384 8820 371390 8832
rect 371513 8823 371571 8829
rect 371513 8820 371525 8823
rect 371384 8792 371525 8820
rect 371384 8780 371390 8792
rect 371513 8789 371525 8792
rect 371559 8820 371571 8823
rect 382918 8820 382924 8832
rect 371559 8792 382924 8820
rect 371559 8789 371571 8792
rect 371513 8783 371571 8789
rect 382918 8780 382924 8792
rect 382976 8780 382982 8832
rect 1104 8730 528816 8752
rect 1104 8678 67574 8730
rect 67626 8678 67638 8730
rect 67690 8678 67702 8730
rect 67754 8678 67766 8730
rect 67818 8678 67830 8730
rect 67882 8678 199502 8730
rect 199554 8678 199566 8730
rect 199618 8678 199630 8730
rect 199682 8678 199694 8730
rect 199746 8678 199758 8730
rect 199810 8678 331430 8730
rect 331482 8678 331494 8730
rect 331546 8678 331558 8730
rect 331610 8678 331622 8730
rect 331674 8678 331686 8730
rect 331738 8678 463358 8730
rect 463410 8678 463422 8730
rect 463474 8678 463486 8730
rect 463538 8678 463550 8730
rect 463602 8678 463614 8730
rect 463666 8678 528816 8730
rect 1104 8656 528816 8678
rect 135254 8576 135260 8628
rect 135312 8616 135318 8628
rect 167546 8616 167552 8628
rect 135312 8588 167552 8616
rect 135312 8576 135318 8588
rect 167546 8576 167552 8588
rect 167604 8576 167610 8628
rect 175366 8576 175372 8628
rect 175424 8616 175430 8628
rect 219894 8616 219900 8628
rect 175424 8588 219900 8616
rect 175424 8576 175430 8588
rect 219894 8576 219900 8588
rect 219952 8576 219958 8628
rect 302418 8576 302424 8628
rect 302476 8576 302482 8628
rect 307478 8576 307484 8628
rect 307536 8576 307542 8628
rect 312446 8576 312452 8628
rect 312504 8576 312510 8628
rect 312906 8576 312912 8628
rect 312964 8616 312970 8628
rect 351914 8616 351920 8628
rect 312964 8588 351920 8616
rect 312964 8576 312970 8588
rect 351914 8576 351920 8588
rect 351972 8576 351978 8628
rect 357894 8576 357900 8628
rect 357952 8616 357958 8628
rect 376846 8616 376852 8628
rect 357952 8588 376852 8616
rect 357952 8576 357958 8588
rect 376846 8576 376852 8588
rect 376904 8576 376910 8628
rect 379146 8576 379152 8628
rect 379204 8616 379210 8628
rect 387058 8616 387064 8628
rect 379204 8588 387064 8616
rect 379204 8576 379210 8588
rect 387058 8576 387064 8588
rect 387116 8576 387122 8628
rect 144457 8551 144515 8557
rect 144457 8548 144469 8551
rect 118666 8520 144469 8548
rect 36078 8372 36084 8424
rect 36136 8412 36142 8424
rect 118666 8412 118694 8520
rect 144457 8517 144469 8520
rect 144503 8517 144515 8551
rect 145742 8548 145748 8560
rect 144457 8511 144515 8517
rect 145024 8520 145748 8548
rect 145024 8489 145052 8520
rect 145742 8508 145748 8520
rect 145800 8508 145806 8560
rect 145834 8508 145840 8560
rect 145892 8548 145898 8560
rect 164329 8551 164387 8557
rect 164329 8548 164341 8551
rect 145892 8520 164341 8548
rect 145892 8508 145898 8520
rect 164329 8517 164341 8520
rect 164375 8517 164387 8551
rect 164329 8511 164387 8517
rect 195606 8508 195612 8560
rect 195664 8548 195670 8560
rect 198642 8548 198648 8560
rect 195664 8520 198648 8548
rect 195664 8508 195670 8520
rect 198642 8508 198648 8520
rect 198700 8508 198706 8560
rect 199194 8508 199200 8560
rect 199252 8548 199258 8560
rect 237374 8548 237380 8560
rect 199252 8520 237380 8548
rect 199252 8508 199258 8520
rect 237374 8508 237380 8520
rect 237432 8508 237438 8560
rect 242158 8508 242164 8560
rect 242216 8548 242222 8560
rect 349338 8548 349344 8560
rect 242216 8520 349344 8548
rect 242216 8508 242222 8520
rect 349338 8508 349344 8520
rect 349396 8508 349402 8560
rect 350074 8508 350080 8560
rect 350132 8548 350138 8560
rect 364978 8548 364984 8560
rect 350132 8520 364984 8548
rect 350132 8508 350138 8520
rect 364978 8508 364984 8520
rect 365036 8508 365042 8560
rect 367278 8508 367284 8560
rect 367336 8548 367342 8560
rect 378134 8548 378140 8560
rect 367336 8520 378140 8548
rect 367336 8508 367342 8520
rect 378134 8508 378140 8520
rect 378192 8508 378198 8560
rect 142065 8483 142123 8489
rect 142065 8449 142077 8483
rect 142111 8449 142123 8483
rect 142065 8443 142123 8449
rect 145009 8483 145067 8489
rect 145009 8449 145021 8483
rect 145055 8449 145067 8483
rect 145009 8443 145067 8449
rect 141513 8415 141571 8421
rect 141513 8412 141525 8415
rect 36136 8384 118694 8412
rect 137986 8384 141525 8412
rect 36136 8372 36142 8384
rect 33502 8304 33508 8356
rect 33560 8344 33566 8356
rect 137986 8344 138014 8384
rect 141513 8381 141525 8384
rect 141559 8381 141571 8415
rect 142080 8412 142108 8443
rect 149698 8440 149704 8492
rect 149756 8440 149762 8492
rect 157245 8483 157303 8489
rect 157245 8449 157257 8483
rect 157291 8480 157303 8483
rect 157886 8480 157892 8492
rect 157291 8452 157892 8480
rect 157291 8449 157303 8452
rect 157245 8443 157303 8449
rect 157886 8440 157892 8452
rect 157944 8440 157950 8492
rect 164881 8483 164939 8489
rect 164881 8449 164893 8483
rect 164927 8480 164939 8483
rect 165525 8483 165583 8489
rect 165525 8480 165537 8483
rect 164927 8452 165537 8480
rect 164927 8449 164939 8452
rect 164881 8443 164939 8449
rect 165525 8449 165537 8452
rect 165571 8480 165583 8483
rect 222470 8480 222476 8492
rect 165571 8452 222476 8480
rect 165571 8449 165583 8452
rect 165525 8443 165583 8449
rect 222470 8440 222476 8452
rect 222528 8440 222534 8492
rect 301777 8483 301835 8489
rect 301777 8449 301789 8483
rect 301823 8480 301835 8483
rect 302418 8480 302424 8492
rect 301823 8452 302424 8480
rect 301823 8449 301835 8452
rect 301777 8443 301835 8449
rect 302418 8440 302424 8452
rect 302476 8440 302482 8492
rect 306374 8440 306380 8492
rect 306432 8440 306438 8492
rect 306837 8483 306895 8489
rect 306837 8449 306849 8483
rect 306883 8480 306895 8483
rect 307478 8480 307484 8492
rect 306883 8452 307484 8480
rect 306883 8449 306895 8452
rect 306837 8443 306895 8449
rect 307478 8440 307484 8452
rect 307536 8440 307542 8492
rect 311250 8440 311256 8492
rect 311308 8440 311314 8492
rect 311805 8483 311863 8489
rect 311805 8449 311817 8483
rect 311851 8480 311863 8483
rect 312446 8480 312452 8492
rect 311851 8452 312452 8480
rect 311851 8449 311863 8452
rect 311805 8443 311863 8449
rect 312446 8440 312452 8452
rect 312504 8440 312510 8492
rect 316310 8440 316316 8492
rect 316368 8440 316374 8492
rect 316865 8483 316923 8489
rect 316865 8449 316877 8483
rect 316911 8480 316923 8483
rect 317506 8480 317512 8492
rect 316911 8452 317512 8480
rect 316911 8449 316923 8452
rect 316865 8443 316923 8449
rect 317506 8440 317512 8452
rect 317564 8440 317570 8492
rect 142709 8415 142767 8421
rect 142709 8412 142721 8415
rect 142080 8384 142721 8412
rect 141513 8375 141571 8381
rect 142709 8381 142721 8384
rect 142755 8412 142767 8415
rect 142755 8384 147674 8412
rect 142755 8381 142767 8384
rect 142709 8375 142767 8381
rect 147646 8344 147674 8384
rect 149054 8372 149060 8424
rect 149112 8412 149118 8424
rect 149149 8415 149207 8421
rect 149149 8412 149161 8415
rect 149112 8384 149161 8412
rect 149112 8372 149118 8384
rect 149149 8381 149161 8384
rect 149195 8381 149207 8415
rect 149149 8375 149207 8381
rect 156690 8372 156696 8424
rect 156748 8372 156754 8424
rect 191466 8372 191472 8424
rect 191524 8412 191530 8424
rect 233878 8412 233884 8424
rect 191524 8384 233884 8412
rect 191524 8372 191530 8384
rect 233878 8372 233884 8384
rect 233936 8372 233942 8424
rect 301222 8372 301228 8424
rect 301280 8372 301286 8424
rect 366266 8372 366272 8424
rect 366324 8412 366330 8424
rect 367462 8412 367468 8424
rect 366324 8384 367468 8412
rect 366324 8372 366330 8384
rect 367462 8372 367468 8384
rect 367520 8372 367526 8424
rect 186314 8344 186320 8356
rect 33560 8316 138014 8344
rect 142540 8316 142752 8344
rect 33560 8304 33566 8316
rect 85574 8236 85580 8288
rect 85632 8276 85638 8288
rect 142540 8276 142568 8316
rect 85632 8248 142568 8276
rect 142724 8276 142752 8316
rect 145576 8316 145788 8344
rect 147646 8316 186320 8344
rect 145576 8276 145604 8316
rect 142724 8248 145604 8276
rect 145760 8276 145788 8316
rect 186314 8304 186320 8316
rect 186372 8304 186378 8356
rect 198734 8304 198740 8356
rect 198792 8344 198798 8356
rect 276014 8344 276020 8356
rect 198792 8316 276020 8344
rect 198792 8304 198798 8316
rect 276014 8304 276020 8316
rect 276072 8304 276078 8356
rect 448330 8344 448336 8356
rect 446968 8316 448336 8344
rect 160094 8276 160100 8288
rect 145760 8248 160100 8276
rect 85632 8236 85638 8248
rect 160094 8236 160100 8248
rect 160152 8236 160158 8288
rect 186498 8236 186504 8288
rect 186556 8276 186562 8288
rect 201954 8276 201960 8288
rect 186556 8248 201960 8276
rect 186556 8236 186562 8248
rect 201954 8236 201960 8248
rect 202012 8236 202018 8288
rect 202046 8236 202052 8288
rect 202104 8276 202110 8288
rect 207474 8276 207480 8288
rect 202104 8248 207480 8276
rect 202104 8236 202110 8248
rect 207474 8236 207480 8248
rect 207532 8236 207538 8288
rect 361482 8236 361488 8288
rect 361540 8276 361546 8288
rect 400950 8276 400956 8288
rect 361540 8248 400956 8276
rect 361540 8236 361546 8248
rect 400950 8236 400956 8248
rect 401008 8236 401014 8288
rect 430206 8236 430212 8288
rect 430264 8276 430270 8288
rect 446968 8276 446996 8316
rect 448330 8304 448336 8316
rect 448388 8304 448394 8356
rect 430264 8248 446996 8276
rect 430264 8236 430270 8248
rect 447042 8236 447048 8288
rect 447100 8276 447106 8288
rect 448054 8276 448060 8288
rect 447100 8248 448060 8276
rect 447100 8236 447106 8248
rect 448054 8236 448060 8248
rect 448112 8236 448118 8288
rect 481818 8236 481824 8288
rect 481876 8276 481882 8288
rect 483106 8276 483112 8288
rect 481876 8248 483112 8276
rect 481876 8236 481882 8248
rect 483106 8236 483112 8248
rect 483164 8236 483170 8288
rect 486142 8236 486148 8288
rect 486200 8276 486206 8288
rect 488534 8276 488540 8288
rect 486200 8248 488540 8276
rect 486200 8236 486206 8248
rect 488534 8236 488540 8248
rect 488592 8236 488598 8288
rect 1104 8186 528816 8208
rect 1104 8134 66914 8186
rect 66966 8134 66978 8186
rect 67030 8134 67042 8186
rect 67094 8134 67106 8186
rect 67158 8134 67170 8186
rect 67222 8134 198842 8186
rect 198894 8134 198906 8186
rect 198958 8134 198970 8186
rect 199022 8134 199034 8186
rect 199086 8134 199098 8186
rect 199150 8134 330770 8186
rect 330822 8134 330834 8186
rect 330886 8134 330898 8186
rect 330950 8134 330962 8186
rect 331014 8134 331026 8186
rect 331078 8134 462698 8186
rect 462750 8134 462762 8186
rect 462814 8134 462826 8186
rect 462878 8134 462890 8186
rect 462942 8134 462954 8186
rect 463006 8134 528816 8186
rect 1104 8112 528816 8134
rect 35894 8032 35900 8084
rect 35952 8072 35958 8084
rect 101033 8075 101091 8081
rect 101033 8072 101045 8075
rect 35952 8044 101045 8072
rect 35952 8032 35958 8044
rect 101033 8041 101045 8044
rect 101079 8072 101091 8075
rect 101306 8072 101312 8084
rect 101079 8044 101312 8072
rect 101079 8041 101091 8044
rect 101033 8035 101091 8041
rect 101306 8032 101312 8044
rect 101364 8032 101370 8084
rect 122558 8032 122564 8084
rect 122616 8032 122622 8084
rect 123294 8032 123300 8084
rect 123352 8072 123358 8084
rect 221642 8072 221648 8084
rect 123352 8044 221648 8072
rect 123352 8032 123358 8044
rect 221642 8032 221648 8044
rect 221700 8032 221706 8084
rect 277118 8032 277124 8084
rect 277176 8032 277182 8084
rect 282270 8032 282276 8084
rect 282328 8032 282334 8084
rect 287146 8032 287152 8084
rect 287204 8072 287210 8084
rect 287422 8072 287428 8084
rect 287204 8044 287428 8072
rect 287204 8032 287210 8044
rect 287422 8032 287428 8044
rect 287480 8032 287486 8084
rect 292574 8032 292580 8084
rect 292632 8032 292638 8084
rect 293862 8032 293868 8084
rect 293920 8072 293926 8084
rect 378410 8072 378416 8084
rect 293920 8044 378416 8072
rect 293920 8032 293926 8044
rect 378410 8032 378416 8044
rect 378468 8032 378474 8084
rect 392118 8032 392124 8084
rect 392176 8072 392182 8084
rect 394694 8072 394700 8084
rect 392176 8044 394700 8072
rect 392176 8032 392182 8044
rect 394694 8032 394700 8044
rect 394752 8032 394758 8084
rect 445570 8032 445576 8084
rect 445628 8072 445634 8084
rect 447042 8072 447048 8084
rect 445628 8044 447048 8072
rect 445628 8032 445634 8044
rect 447042 8032 447048 8044
rect 447100 8032 447106 8084
rect 481726 8032 481732 8084
rect 481784 8072 481790 8084
rect 484486 8072 484492 8084
rect 481784 8044 484492 8072
rect 481784 8032 481790 8044
rect 484486 8032 484492 8044
rect 484544 8032 484550 8084
rect 487522 8032 487528 8084
rect 487580 8072 487586 8084
rect 501322 8072 501328 8084
rect 487580 8044 501328 8072
rect 487580 8032 487586 8044
rect 501322 8032 501328 8044
rect 501380 8032 501386 8084
rect 59262 7964 59268 8016
rect 59320 8004 59326 8016
rect 135254 8004 135260 8016
rect 59320 7976 135260 8004
rect 59320 7964 59326 7976
rect 135254 7964 135260 7976
rect 135312 7964 135318 8016
rect 139026 7964 139032 8016
rect 139084 8004 139090 8016
rect 246114 8004 246120 8016
rect 139084 7976 246120 8004
rect 139084 7964 139090 7976
rect 246114 7964 246120 7976
rect 246172 7964 246178 8016
rect 267642 7964 267648 8016
rect 267700 8004 267706 8016
rect 364242 8004 364248 8016
rect 267700 7976 364248 8004
rect 267700 7964 267706 7976
rect 364242 7964 364248 7976
rect 364300 7964 364306 8016
rect 365714 7964 365720 8016
rect 365772 8004 365778 8016
rect 371786 8004 371792 8016
rect 365772 7976 371792 8004
rect 365772 7964 365778 7976
rect 371786 7964 371792 7976
rect 371844 7964 371850 8016
rect 372522 7964 372528 8016
rect 372580 8004 372586 8016
rect 376202 8004 376208 8016
rect 372580 7976 376208 8004
rect 372580 7964 372586 7976
rect 376202 7964 376208 7976
rect 376260 7964 376266 8016
rect 382274 7964 382280 8016
rect 382332 8004 382338 8016
rect 402330 8004 402336 8016
rect 382332 7976 402336 8004
rect 382332 7964 382338 7976
rect 402330 7964 402336 7976
rect 402388 7964 402394 8016
rect 426158 7964 426164 8016
rect 426216 8004 426222 8016
rect 447778 8004 447784 8016
rect 426216 7976 447784 8004
rect 426216 7964 426222 7976
rect 447778 7964 447784 7976
rect 447836 7964 447842 8016
rect 482002 7964 482008 8016
rect 482060 8004 482066 8016
rect 485038 8004 485044 8016
rect 482060 7976 485044 8004
rect 482060 7964 482066 7976
rect 485038 7964 485044 7976
rect 485096 7964 485102 8016
rect 486970 7964 486976 8016
rect 487028 8004 487034 8016
rect 496170 8004 496176 8016
rect 487028 7976 496176 8004
rect 487028 7964 487034 7976
rect 496170 7964 496176 7976
rect 496228 7964 496234 8016
rect 22462 7896 22468 7948
rect 22520 7936 22526 7948
rect 99466 7936 99472 7948
rect 22520 7908 99472 7936
rect 22520 7896 22526 7908
rect 99466 7896 99472 7908
rect 99524 7896 99530 7948
rect 120994 7896 121000 7948
rect 121052 7936 121058 7948
rect 228450 7936 228456 7948
rect 121052 7908 228456 7936
rect 121052 7896 121058 7908
rect 228450 7896 228456 7908
rect 228508 7896 228514 7948
rect 276014 7896 276020 7948
rect 276072 7896 276078 7948
rect 276124 7908 350534 7936
rect 71038 7828 71044 7880
rect 71096 7868 71102 7880
rect 86310 7868 86316 7880
rect 71096 7840 86316 7868
rect 71096 7828 71102 7840
rect 86310 7828 86316 7840
rect 86368 7828 86374 7880
rect 91370 7868 91376 7880
rect 86420 7840 91376 7868
rect 42978 7760 42984 7812
rect 43036 7800 43042 7812
rect 86420 7800 86448 7840
rect 91370 7828 91376 7840
rect 91428 7828 91434 7880
rect 91649 7871 91707 7877
rect 91649 7868 91661 7871
rect 91480 7840 91661 7868
rect 91278 7800 91284 7812
rect 43036 7772 86448 7800
rect 86512 7772 91284 7800
rect 43036 7760 43042 7772
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 86512 7732 86540 7772
rect 91278 7760 91284 7772
rect 91336 7760 91342 7812
rect 14792 7704 86540 7732
rect 14792 7692 14798 7704
rect 86586 7692 86592 7744
rect 86644 7732 86650 7744
rect 91480 7732 91508 7840
rect 91649 7837 91661 7840
rect 91695 7868 91707 7871
rect 92293 7871 92351 7877
rect 92293 7868 92305 7871
rect 91695 7840 92305 7868
rect 91695 7837 91707 7840
rect 91649 7831 91707 7837
rect 92293 7837 92305 7840
rect 92339 7837 92351 7871
rect 96706 7868 96712 7880
rect 92293 7831 92351 7837
rect 92768 7840 96712 7868
rect 91830 7760 91836 7812
rect 91888 7800 91894 7812
rect 92768 7800 92796 7840
rect 96706 7828 96712 7840
rect 96764 7828 96770 7880
rect 114189 7871 114247 7877
rect 114189 7837 114201 7871
rect 114235 7868 114247 7871
rect 114830 7868 114836 7880
rect 114235 7840 114836 7868
rect 114235 7837 114247 7840
rect 114189 7831 114247 7837
rect 114830 7828 114836 7840
rect 114888 7828 114894 7880
rect 121825 7871 121883 7877
rect 121825 7837 121837 7871
rect 121871 7868 121883 7871
rect 122558 7868 122564 7880
rect 121871 7840 122564 7868
rect 121871 7837 121883 7840
rect 121825 7831 121883 7837
rect 122558 7828 122564 7840
rect 122616 7828 122622 7880
rect 126885 7871 126943 7877
rect 126885 7837 126897 7871
rect 126931 7868 126943 7871
rect 131945 7871 132003 7877
rect 126931 7840 127756 7868
rect 126931 7837 126943 7840
rect 126885 7831 126943 7837
rect 91888 7772 92796 7800
rect 91888 7760 91894 7772
rect 92842 7760 92848 7812
rect 92900 7760 92906 7812
rect 92952 7772 103514 7800
rect 86644 7704 91508 7732
rect 86644 7692 86650 7704
rect 91738 7692 91744 7744
rect 91796 7732 91802 7744
rect 92952 7732 92980 7772
rect 91796 7704 92980 7732
rect 91796 7692 91802 7704
rect 94038 7692 94044 7744
rect 94096 7692 94102 7744
rect 95234 7692 95240 7744
rect 95292 7692 95298 7744
rect 97626 7692 97632 7744
rect 97684 7692 97690 7744
rect 103486 7732 103514 7772
rect 113634 7760 113640 7812
rect 113692 7760 113698 7812
rect 121273 7803 121331 7809
rect 121273 7800 121285 7803
rect 113744 7772 121285 7800
rect 113744 7732 113772 7772
rect 121273 7769 121285 7772
rect 121319 7769 121331 7803
rect 121273 7763 121331 7769
rect 126330 7760 126336 7812
rect 126388 7760 126394 7812
rect 127728 7744 127756 7840
rect 131945 7837 131957 7871
rect 131991 7837 132003 7871
rect 131945 7831 132003 7837
rect 131390 7760 131396 7812
rect 131448 7760 131454 7812
rect 131960 7800 131988 7831
rect 132034 7828 132040 7880
rect 132092 7868 132098 7880
rect 137005 7871 137063 7877
rect 132092 7840 136772 7868
rect 132092 7828 132098 7840
rect 131960 7772 132908 7800
rect 132880 7744 132908 7772
rect 136634 7760 136640 7812
rect 136692 7760 136698 7812
rect 136744 7800 136772 7840
rect 137005 7837 137017 7871
rect 137051 7868 137063 7871
rect 138017 7871 138075 7877
rect 138017 7868 138029 7871
rect 137051 7840 138029 7868
rect 137051 7837 137063 7840
rect 137005 7831 137063 7837
rect 138017 7837 138029 7840
rect 138063 7868 138075 7871
rect 141234 7868 141240 7880
rect 138063 7840 141240 7868
rect 138063 7837 138075 7840
rect 138017 7831 138075 7837
rect 141234 7828 141240 7840
rect 141292 7828 141298 7880
rect 149698 7828 149704 7880
rect 149756 7868 149762 7880
rect 149885 7871 149943 7877
rect 149885 7868 149897 7871
rect 149756 7840 149897 7868
rect 149756 7828 149762 7840
rect 149885 7837 149897 7840
rect 149931 7837 149943 7871
rect 149885 7831 149943 7837
rect 268378 7828 268384 7880
rect 268436 7868 268442 7880
rect 276124 7868 276152 7908
rect 268436 7840 276152 7868
rect 276385 7871 276443 7877
rect 268436 7828 268442 7840
rect 276385 7837 276397 7871
rect 276431 7868 276443 7871
rect 277118 7868 277124 7880
rect 276431 7840 277124 7868
rect 276431 7837 276443 7840
rect 276385 7831 276443 7837
rect 277118 7828 277124 7840
rect 277176 7828 277182 7880
rect 281537 7871 281595 7877
rect 281537 7837 281549 7871
rect 281583 7868 281595 7871
rect 282270 7868 282276 7880
rect 281583 7840 282276 7868
rect 281583 7837 281595 7840
rect 281537 7831 281595 7837
rect 282270 7828 282276 7840
rect 282328 7828 282334 7880
rect 286689 7871 286747 7877
rect 286689 7837 286701 7871
rect 286735 7868 286747 7871
rect 287146 7868 287152 7880
rect 286735 7840 287152 7868
rect 286735 7837 286747 7840
rect 286689 7831 286747 7837
rect 287146 7828 287152 7840
rect 287204 7828 287210 7880
rect 291749 7871 291807 7877
rect 287256 7840 291332 7868
rect 239490 7800 239496 7812
rect 136744 7772 239496 7800
rect 239490 7760 239496 7772
rect 239548 7760 239554 7812
rect 275940 7772 277394 7800
rect 103486 7704 113772 7732
rect 114830 7692 114836 7744
rect 114888 7692 114894 7744
rect 127710 7692 127716 7744
rect 127768 7692 127774 7744
rect 132862 7692 132868 7744
rect 132920 7692 132926 7744
rect 186590 7692 186596 7744
rect 186648 7732 186654 7744
rect 234982 7732 234988 7744
rect 186648 7704 234988 7732
rect 186648 7692 186654 7704
rect 234982 7692 234988 7704
rect 235040 7692 235046 7744
rect 251361 7735 251419 7741
rect 251361 7701 251373 7735
rect 251407 7732 251419 7735
rect 251450 7732 251456 7744
rect 251407 7704 251456 7732
rect 251407 7701 251419 7704
rect 251361 7695 251419 7701
rect 251450 7692 251456 7704
rect 251508 7692 251514 7744
rect 252462 7692 252468 7744
rect 252520 7692 252526 7744
rect 258350 7692 258356 7744
rect 258408 7732 258414 7744
rect 275940 7732 275968 7772
rect 258408 7704 275968 7732
rect 277366 7732 277394 7772
rect 280338 7760 280344 7812
rect 280396 7800 280402 7812
rect 280985 7803 281043 7809
rect 280985 7800 280997 7803
rect 280396 7772 280997 7800
rect 280396 7760 280402 7772
rect 280985 7769 280997 7772
rect 281031 7769 281043 7803
rect 280985 7763 281043 7769
rect 281092 7772 282316 7800
rect 281092 7732 281120 7772
rect 277366 7704 281120 7732
rect 282288 7732 282316 7772
rect 286134 7760 286140 7812
rect 286192 7760 286198 7812
rect 287256 7732 287284 7840
rect 291194 7760 291200 7812
rect 291252 7760 291258 7812
rect 291304 7800 291332 7840
rect 291749 7837 291761 7871
rect 291795 7868 291807 7871
rect 292574 7868 292580 7880
rect 291795 7840 292580 7868
rect 291795 7837 291807 7840
rect 291749 7831 291807 7837
rect 292574 7828 292580 7840
rect 292632 7828 292638 7880
rect 296717 7871 296775 7877
rect 296717 7837 296729 7871
rect 296763 7868 296775 7871
rect 297726 7868 297732 7880
rect 296763 7840 297732 7868
rect 296763 7837 296775 7840
rect 296717 7831 296775 7837
rect 297726 7828 297732 7840
rect 297784 7828 297790 7880
rect 350506 7868 350534 7908
rect 364702 7896 364708 7948
rect 364760 7936 364766 7948
rect 364760 7908 366680 7936
rect 364760 7896 364766 7908
rect 366266 7868 366272 7880
rect 350506 7840 366272 7868
rect 366266 7828 366272 7840
rect 366324 7828 366330 7880
rect 366652 7868 366680 7908
rect 367094 7896 367100 7948
rect 367152 7936 367158 7948
rect 372890 7936 372896 7948
rect 367152 7908 372896 7936
rect 367152 7896 367158 7908
rect 372890 7896 372896 7908
rect 372948 7896 372954 7948
rect 375558 7896 375564 7948
rect 375616 7936 375622 7948
rect 400674 7936 400680 7948
rect 375616 7908 400680 7936
rect 375616 7896 375622 7908
rect 400674 7896 400680 7908
rect 400732 7896 400738 7948
rect 480438 7896 480444 7948
rect 480496 7936 480502 7948
rect 483658 7936 483664 7948
rect 480496 7908 483664 7936
rect 480496 7896 480502 7908
rect 483658 7896 483664 7908
rect 483716 7896 483722 7948
rect 487798 7896 487804 7948
rect 487856 7936 487862 7948
rect 503898 7936 503904 7948
rect 487856 7908 503904 7936
rect 487856 7896 487862 7908
rect 503898 7896 503904 7908
rect 503956 7896 503962 7948
rect 392854 7868 392860 7880
rect 366652 7840 392860 7868
rect 392854 7828 392860 7840
rect 392912 7828 392918 7880
rect 419902 7828 419908 7880
rect 419960 7868 419966 7880
rect 447226 7868 447232 7880
rect 419960 7840 447232 7868
rect 419960 7828 419966 7840
rect 447226 7828 447232 7840
rect 447284 7828 447290 7880
rect 487246 7828 487252 7880
rect 487304 7868 487310 7880
rect 498746 7868 498752 7880
rect 487304 7840 498752 7868
rect 487304 7828 487310 7840
rect 498746 7828 498752 7840
rect 498804 7828 498810 7880
rect 291304 7772 292620 7800
rect 282288 7704 287284 7732
rect 292592 7732 292620 7772
rect 296162 7760 296168 7812
rect 296220 7760 296226 7812
rect 366358 7800 366364 7812
rect 296686 7772 366364 7800
rect 296686 7732 296714 7772
rect 366358 7760 366364 7772
rect 366416 7760 366422 7812
rect 368474 7760 368480 7812
rect 368532 7800 368538 7812
rect 373994 7800 374000 7812
rect 368532 7772 374000 7800
rect 368532 7760 368538 7772
rect 373994 7760 374000 7772
rect 374052 7760 374058 7812
rect 374270 7760 374276 7812
rect 374328 7800 374334 7812
rect 393498 7800 393504 7812
rect 374328 7772 393504 7800
rect 374328 7760 374334 7772
rect 393498 7760 393504 7772
rect 393556 7760 393562 7812
rect 393958 7760 393964 7812
rect 394016 7800 394022 7812
rect 440142 7800 440148 7812
rect 394016 7772 440148 7800
rect 394016 7760 394022 7772
rect 440142 7760 440148 7772
rect 440200 7760 440206 7812
rect 488074 7760 488080 7812
rect 488132 7800 488138 7812
rect 506474 7800 506480 7812
rect 488132 7772 506480 7800
rect 488132 7760 488138 7772
rect 506474 7760 506480 7772
rect 506532 7760 506538 7812
rect 292592 7704 296714 7732
rect 258408 7692 258414 7704
rect 349062 7692 349068 7744
rect 349120 7732 349126 7744
rect 403894 7732 403900 7744
rect 349120 7704 403900 7732
rect 349120 7692 349126 7704
rect 403894 7692 403900 7704
rect 403952 7692 403958 7744
rect 414750 7692 414756 7744
rect 414808 7732 414814 7744
rect 446674 7732 446680 7744
rect 414808 7704 446680 7732
rect 414808 7692 414814 7704
rect 446674 7692 446680 7704
rect 446732 7692 446738 7744
rect 488350 7692 488356 7744
rect 488408 7732 488414 7744
rect 509050 7732 509056 7744
rect 488408 7704 509056 7732
rect 488408 7692 488414 7704
rect 509050 7692 509056 7704
rect 509108 7692 509114 7744
rect 1104 7642 528816 7664
rect 1104 7590 67574 7642
rect 67626 7590 67638 7642
rect 67690 7590 67702 7642
rect 67754 7590 67766 7642
rect 67818 7590 67830 7642
rect 67882 7590 199502 7642
rect 199554 7590 199566 7642
rect 199618 7590 199630 7642
rect 199682 7590 199694 7642
rect 199746 7590 199758 7642
rect 199810 7590 331430 7642
rect 331482 7590 331494 7642
rect 331546 7590 331558 7642
rect 331610 7590 331622 7642
rect 331674 7590 331686 7642
rect 331738 7590 463358 7642
rect 463410 7590 463422 7642
rect 463474 7590 463486 7642
rect 463538 7590 463550 7642
rect 463602 7590 463614 7642
rect 463666 7590 528816 7642
rect 1104 7568 528816 7590
rect 29914 7488 29920 7540
rect 29972 7528 29978 7540
rect 97626 7528 97632 7540
rect 29972 7500 97632 7528
rect 29972 7488 29978 7500
rect 97626 7488 97632 7500
rect 97684 7528 97690 7540
rect 126330 7528 126336 7540
rect 97684 7500 97948 7528
rect 97684 7488 97690 7500
rect 63494 7420 63500 7472
rect 63552 7460 63558 7472
rect 95234 7460 95240 7472
rect 63552 7432 95240 7460
rect 63552 7420 63558 7432
rect 95234 7420 95240 7432
rect 95292 7460 95298 7472
rect 95292 7432 95556 7460
rect 95292 7420 95298 7432
rect 91189 7395 91247 7401
rect 91189 7392 91201 7395
rect 90560 7364 91201 7392
rect 90560 7200 90588 7364
rect 91189 7361 91201 7364
rect 91235 7361 91247 7395
rect 91189 7355 91247 7361
rect 91741 7395 91799 7401
rect 91741 7361 91753 7395
rect 91787 7392 91799 7395
rect 92198 7392 92204 7404
rect 91787 7364 92204 7392
rect 91787 7361 91799 7364
rect 91741 7355 91799 7361
rect 92198 7352 92204 7364
rect 92256 7352 92262 7404
rect 92937 7395 92995 7401
rect 92937 7392 92949 7395
rect 92308 7364 92949 7392
rect 92308 7200 92336 7364
rect 92937 7361 92949 7364
rect 92983 7361 92995 7395
rect 92937 7355 92995 7361
rect 93486 7352 93492 7404
rect 93544 7352 93550 7404
rect 95528 7401 95556 7432
rect 96062 7420 96068 7472
rect 96120 7420 96126 7472
rect 97258 7420 97264 7472
rect 97316 7420 97322 7472
rect 94317 7395 94375 7401
rect 94317 7361 94329 7395
rect 94363 7361 94375 7395
rect 94317 7355 94375 7361
rect 95513 7395 95571 7401
rect 95513 7361 95525 7395
rect 95559 7361 95571 7395
rect 95513 7355 95571 7361
rect 92382 7284 92388 7336
rect 92440 7324 92446 7336
rect 94038 7324 94044 7336
rect 92440 7296 94044 7324
rect 92440 7284 92446 7296
rect 94038 7284 94044 7296
rect 94096 7324 94102 7336
rect 94332 7324 94360 7355
rect 96706 7352 96712 7404
rect 96764 7352 96770 7404
rect 97920 7401 97948 7500
rect 99346 7500 126336 7528
rect 98454 7420 98460 7472
rect 98512 7420 98518 7472
rect 97905 7395 97963 7401
rect 97905 7361 97917 7395
rect 97951 7361 97963 7395
rect 97905 7355 97963 7361
rect 94096 7296 94360 7324
rect 94096 7284 94102 7296
rect 94866 7284 94872 7336
rect 94924 7284 94930 7336
rect 96614 7284 96620 7336
rect 96672 7324 96678 7336
rect 99346 7324 99374 7500
rect 126330 7488 126336 7500
rect 126388 7488 126394 7540
rect 127710 7488 127716 7540
rect 127768 7528 127774 7540
rect 201494 7528 201500 7540
rect 127768 7500 201500 7528
rect 127768 7488 127774 7500
rect 201494 7488 201500 7500
rect 201552 7488 201558 7540
rect 237006 7488 237012 7540
rect 237064 7528 237070 7540
rect 237064 7500 253934 7528
rect 237064 7488 237070 7500
rect 101858 7420 101864 7472
rect 101916 7420 101922 7472
rect 131390 7460 131396 7472
rect 103486 7432 131396 7460
rect 99466 7352 99472 7404
rect 99524 7392 99530 7404
rect 100113 7395 100171 7401
rect 100113 7392 100125 7395
rect 99524 7364 100125 7392
rect 99524 7352 99530 7364
rect 100113 7361 100125 7364
rect 100159 7361 100171 7395
rect 100113 7355 100171 7361
rect 100662 7352 100668 7404
rect 100720 7352 100726 7404
rect 101306 7352 101312 7404
rect 101364 7352 101370 7404
rect 103486 7392 103514 7432
rect 131390 7420 131396 7432
rect 131448 7420 131454 7472
rect 141234 7420 141240 7472
rect 141292 7460 141298 7472
rect 210694 7460 210700 7472
rect 141292 7432 210700 7460
rect 141292 7420 141298 7432
rect 210694 7420 210700 7432
rect 210752 7420 210758 7472
rect 250806 7420 250812 7472
rect 250864 7420 250870 7472
rect 253906 7460 253934 7500
rect 256970 7488 256976 7540
rect 257028 7488 257034 7540
rect 262030 7488 262036 7540
rect 262088 7488 262094 7540
rect 267090 7488 267096 7540
rect 267148 7488 267154 7540
rect 272150 7488 272156 7540
rect 272208 7488 272214 7540
rect 358814 7488 358820 7540
rect 358872 7528 358878 7540
rect 368658 7528 368664 7540
rect 358872 7500 368664 7528
rect 358872 7488 358878 7500
rect 368658 7488 368664 7500
rect 368716 7488 368722 7540
rect 370774 7488 370780 7540
rect 370832 7528 370838 7540
rect 375098 7528 375104 7540
rect 370832 7500 375104 7528
rect 370832 7488 370838 7500
rect 375098 7488 375104 7500
rect 375156 7488 375162 7540
rect 375374 7488 375380 7540
rect 375432 7528 375438 7540
rect 394050 7528 394056 7540
rect 375432 7500 394056 7528
rect 375432 7488 375438 7500
rect 394050 7488 394056 7500
rect 394108 7488 394114 7540
rect 486418 7488 486424 7540
rect 486476 7528 486482 7540
rect 491018 7528 491024 7540
rect 486476 7500 491024 7528
rect 486476 7488 486482 7500
rect 491018 7488 491024 7500
rect 491076 7488 491082 7540
rect 344094 7460 344100 7472
rect 253906 7432 344100 7460
rect 344094 7420 344100 7432
rect 344152 7420 344158 7472
rect 362310 7420 362316 7472
rect 362368 7460 362374 7472
rect 369762 7460 369768 7472
rect 362368 7432 369768 7460
rect 362368 7420 362374 7432
rect 369762 7420 369768 7432
rect 369820 7420 369826 7472
rect 373442 7420 373448 7472
rect 373500 7460 373506 7472
rect 377306 7460 377312 7472
rect 373500 7432 377312 7460
rect 373500 7420 373506 7432
rect 377306 7420 377312 7432
rect 377364 7420 377370 7472
rect 486694 7420 486700 7472
rect 486752 7460 486758 7472
rect 493594 7460 493600 7472
rect 486752 7432 493600 7460
rect 486752 7420 486758 7432
rect 493594 7420 493600 7432
rect 493652 7420 493658 7472
rect 102152 7364 103514 7392
rect 96672 7296 99374 7324
rect 96672 7284 96678 7296
rect 90542 7148 90548 7200
rect 90600 7148 90606 7200
rect 92290 7148 92296 7200
rect 92348 7148 92354 7200
rect 96706 7148 96712 7200
rect 96764 7188 96770 7200
rect 102152 7188 102180 7364
rect 114830 7352 114836 7404
rect 114888 7392 114894 7404
rect 187878 7392 187884 7404
rect 114888 7364 187884 7392
rect 114888 7352 114894 7364
rect 187878 7352 187884 7364
rect 187936 7352 187942 7404
rect 189166 7352 189172 7404
rect 189224 7392 189230 7404
rect 208578 7392 208584 7404
rect 189224 7364 208584 7392
rect 189224 7352 189230 7364
rect 208578 7352 208584 7364
rect 208636 7352 208642 7404
rect 250257 7395 250315 7401
rect 250257 7392 250269 7395
rect 249628 7364 250269 7392
rect 102226 7216 102232 7268
rect 102284 7256 102290 7268
rect 113634 7256 113640 7268
rect 102284 7228 113640 7256
rect 102284 7216 102290 7228
rect 113634 7216 113640 7228
rect 113692 7216 113698 7268
rect 123478 7216 123484 7268
rect 123536 7256 123542 7268
rect 218330 7256 218336 7268
rect 123536 7228 218336 7256
rect 123536 7216 123542 7228
rect 218330 7216 218336 7228
rect 218388 7216 218394 7268
rect 96764 7160 102180 7188
rect 96764 7148 96770 7160
rect 103238 7148 103244 7200
rect 103296 7148 103302 7200
rect 113358 7148 113364 7200
rect 113416 7148 113422 7200
rect 118510 7148 118516 7200
rect 118568 7188 118574 7200
rect 226426 7188 226432 7200
rect 118568 7160 226432 7188
rect 118568 7148 118574 7160
rect 226426 7148 226432 7160
rect 226484 7148 226490 7200
rect 249518 7148 249524 7200
rect 249576 7188 249582 7200
rect 249628 7197 249656 7364
rect 250257 7361 250269 7364
rect 250303 7361 250315 7395
rect 250257 7355 250315 7361
rect 251450 7352 251456 7404
rect 251508 7352 251514 7404
rect 252462 7352 252468 7404
rect 252520 7392 252526 7404
rect 252649 7395 252707 7401
rect 252649 7392 252661 7395
rect 252520 7364 252661 7392
rect 252520 7352 252526 7364
rect 252649 7361 252661 7364
rect 252695 7361 252707 7395
rect 252649 7355 252707 7361
rect 253934 7352 253940 7404
rect 253992 7392 253998 7404
rect 254213 7395 254271 7401
rect 254213 7392 254225 7395
rect 253992 7364 254225 7392
rect 253992 7352 253998 7364
rect 254213 7361 254225 7364
rect 254259 7361 254271 7395
rect 254213 7355 254271 7361
rect 254765 7395 254823 7401
rect 254765 7361 254777 7395
rect 254811 7392 254823 7395
rect 255222 7392 255228 7404
rect 254811 7364 255228 7392
rect 254811 7361 254823 7364
rect 254765 7355 254823 7361
rect 255222 7352 255228 7364
rect 255280 7352 255286 7404
rect 256329 7395 256387 7401
rect 256329 7361 256341 7395
rect 256375 7392 256387 7395
rect 256970 7392 256976 7404
rect 256375 7364 256976 7392
rect 256375 7361 256387 7364
rect 256329 7355 256387 7361
rect 256970 7352 256976 7364
rect 257028 7352 257034 7404
rect 260834 7352 260840 7404
rect 260892 7352 260898 7404
rect 261389 7395 261447 7401
rect 261389 7361 261401 7395
rect 261435 7392 261447 7395
rect 262030 7392 262036 7404
rect 261435 7364 262036 7392
rect 261435 7361 261447 7364
rect 261389 7355 261447 7361
rect 262030 7352 262036 7364
rect 262088 7352 262094 7404
rect 266449 7395 266507 7401
rect 266449 7361 266461 7395
rect 266495 7392 266507 7395
rect 267090 7392 267096 7404
rect 266495 7364 267096 7392
rect 266495 7361 266507 7364
rect 266449 7355 266507 7361
rect 267090 7352 267096 7364
rect 267148 7352 267154 7404
rect 270954 7352 270960 7404
rect 271012 7352 271018 7404
rect 271509 7395 271567 7401
rect 271509 7361 271521 7395
rect 271555 7392 271567 7395
rect 272150 7392 272156 7404
rect 271555 7364 272156 7392
rect 271555 7361 271567 7364
rect 271509 7355 271567 7361
rect 272150 7352 272156 7364
rect 272208 7352 272214 7404
rect 364978 7352 364984 7404
rect 365036 7392 365042 7404
rect 370682 7392 370688 7404
rect 365036 7364 370688 7392
rect 365036 7352 365042 7364
rect 370682 7352 370688 7364
rect 370740 7352 370746 7404
rect 252002 7284 252008 7336
rect 252060 7284 252066 7336
rect 253201 7327 253259 7333
rect 253201 7293 253213 7327
rect 253247 7324 253259 7327
rect 253247 7296 253934 7324
rect 253247 7293 253259 7296
rect 253201 7287 253259 7293
rect 253906 7256 253934 7296
rect 255774 7284 255780 7336
rect 255832 7284 255838 7336
rect 264974 7284 264980 7336
rect 265032 7324 265038 7336
rect 265897 7327 265955 7333
rect 265897 7324 265909 7327
rect 265032 7296 265909 7324
rect 265032 7284 265038 7296
rect 265897 7293 265909 7296
rect 265943 7293 265955 7327
rect 265897 7287 265955 7293
rect 362034 7256 362040 7268
rect 253906 7228 362040 7256
rect 362034 7216 362040 7228
rect 362092 7216 362098 7268
rect 249613 7191 249671 7197
rect 249613 7188 249625 7191
rect 249576 7160 249625 7188
rect 249576 7148 249582 7160
rect 249613 7157 249625 7160
rect 249659 7157 249671 7191
rect 249613 7151 249671 7157
rect 1104 7098 528816 7120
rect 1104 7046 66914 7098
rect 66966 7046 66978 7098
rect 67030 7046 67042 7098
rect 67094 7046 67106 7098
rect 67158 7046 67170 7098
rect 67222 7046 198842 7098
rect 198894 7046 198906 7098
rect 198958 7046 198970 7098
rect 199022 7046 199034 7098
rect 199086 7046 199098 7098
rect 199150 7046 330770 7098
rect 330822 7046 330834 7098
rect 330886 7046 330898 7098
rect 330950 7046 330962 7098
rect 331014 7046 331026 7098
rect 331078 7046 462698 7098
rect 462750 7046 462762 7098
rect 462814 7046 462826 7098
rect 462878 7046 462890 7098
rect 462942 7046 462954 7098
rect 463006 7046 528816 7098
rect 1104 7024 528816 7046
rect 46934 6944 46940 6996
rect 46992 6984 46998 6996
rect 90542 6984 90548 6996
rect 46992 6956 90548 6984
rect 46992 6944 46998 6956
rect 90542 6944 90548 6956
rect 90600 6944 90606 6996
rect 94866 6944 94872 6996
rect 94924 6984 94930 6996
rect 186682 6984 186688 6996
rect 94924 6956 186688 6984
rect 94924 6944 94930 6956
rect 186682 6944 186688 6956
rect 186740 6944 186746 6996
rect 262214 6944 262220 6996
rect 262272 6984 262278 6996
rect 365254 6984 365260 6996
rect 262272 6956 365260 6984
rect 262272 6944 262278 6956
rect 365254 6944 365260 6956
rect 365312 6944 365318 6996
rect 78674 6876 78680 6928
rect 78732 6916 78738 6928
rect 92290 6916 92296 6928
rect 78732 6888 92296 6916
rect 78732 6876 78738 6888
rect 92290 6876 92296 6888
rect 92348 6876 92354 6928
rect 94498 6876 94504 6928
rect 94556 6916 94562 6928
rect 102226 6916 102232 6928
rect 94556 6888 102232 6916
rect 94556 6876 94562 6888
rect 102226 6876 102232 6888
rect 102284 6876 102290 6928
rect 124953 6919 125011 6925
rect 124953 6885 124965 6919
rect 124999 6916 125011 6919
rect 125134 6916 125140 6928
rect 124999 6888 125140 6916
rect 124999 6885 125011 6888
rect 124953 6879 125011 6885
rect 125134 6876 125140 6888
rect 125192 6876 125198 6928
rect 196710 6876 196716 6928
rect 196768 6916 196774 6928
rect 202690 6916 202696 6928
rect 196768 6888 202696 6916
rect 196768 6876 196774 6888
rect 202690 6876 202696 6888
rect 202748 6876 202754 6928
rect 252002 6876 252008 6928
rect 252060 6916 252066 6928
rect 360930 6916 360936 6928
rect 252060 6888 360936 6916
rect 252060 6876 252066 6888
rect 360930 6876 360936 6888
rect 360988 6876 360994 6928
rect 33134 6808 33140 6860
rect 33192 6848 33198 6860
rect 33192 6820 102456 6848
rect 33192 6808 33198 6820
rect 91649 6783 91707 6789
rect 91649 6780 91661 6783
rect 90928 6752 91661 6780
rect 90928 6656 90956 6752
rect 91649 6749 91661 6752
rect 91695 6749 91707 6783
rect 91649 6743 91707 6749
rect 92106 6740 92112 6792
rect 92164 6740 92170 6792
rect 93397 6783 93455 6789
rect 93397 6780 93409 6783
rect 92768 6752 93409 6780
rect 92768 6656 92796 6752
rect 93397 6749 93409 6752
rect 93443 6749 93455 6783
rect 93397 6743 93455 6749
rect 93762 6740 93768 6792
rect 93820 6740 93826 6792
rect 94314 6740 94320 6792
rect 94372 6780 94378 6792
rect 94593 6783 94651 6789
rect 94593 6780 94605 6783
rect 94372 6752 94605 6780
rect 94372 6740 94378 6752
rect 94593 6749 94605 6752
rect 94639 6749 94651 6783
rect 94593 6743 94651 6749
rect 95142 6740 95148 6792
rect 95200 6740 95206 6792
rect 96798 6740 96804 6792
rect 96856 6780 96862 6792
rect 96893 6783 96951 6789
rect 96893 6780 96905 6783
rect 96856 6752 96905 6780
rect 96856 6740 96862 6752
rect 96893 6749 96905 6752
rect 96939 6749 96951 6783
rect 96893 6743 96951 6749
rect 97442 6740 97448 6792
rect 97500 6740 97506 6792
rect 99009 6783 99067 6789
rect 99009 6780 99021 6783
rect 98380 6752 99021 6780
rect 98380 6656 98408 6752
rect 99009 6749 99021 6752
rect 99055 6749 99067 6783
rect 102321 6783 102379 6789
rect 102321 6780 102333 6783
rect 99009 6743 99067 6749
rect 101232 6752 102333 6780
rect 99561 6715 99619 6721
rect 99561 6681 99573 6715
rect 99607 6712 99619 6715
rect 100662 6712 100668 6724
rect 99607 6684 100668 6712
rect 99607 6681 99619 6684
rect 99561 6675 99619 6681
rect 100662 6672 100668 6684
rect 100720 6672 100726 6724
rect 101232 6656 101260 6752
rect 102321 6749 102333 6752
rect 102367 6749 102379 6783
rect 102428 6780 102456 6820
rect 102870 6808 102876 6860
rect 102928 6808 102934 6860
rect 104066 6808 104072 6860
rect 104124 6808 104130 6860
rect 105265 6851 105323 6857
rect 105265 6817 105277 6851
rect 105311 6848 105323 6851
rect 108577 6851 108635 6857
rect 105311 6820 108528 6848
rect 105311 6817 105323 6820
rect 105265 6811 105323 6817
rect 103238 6780 103244 6792
rect 102428 6752 103244 6780
rect 102321 6743 102379 6749
rect 103238 6740 103244 6752
rect 103296 6780 103302 6792
rect 103517 6783 103575 6789
rect 103517 6780 103529 6783
rect 103296 6752 103529 6780
rect 103296 6740 103302 6752
rect 103517 6749 103529 6752
rect 103563 6749 103575 6783
rect 103517 6743 103575 6749
rect 104434 6740 104440 6792
rect 104492 6780 104498 6792
rect 104713 6783 104771 6789
rect 104713 6780 104725 6783
rect 104492 6752 104725 6780
rect 104492 6740 104498 6752
rect 104713 6749 104725 6752
rect 104759 6749 104771 6783
rect 104713 6743 104771 6749
rect 108025 6783 108083 6789
rect 108025 6749 108037 6783
rect 108071 6749 108083 6783
rect 108025 6743 108083 6749
rect 107286 6672 107292 6724
rect 107344 6712 107350 6724
rect 107473 6715 107531 6721
rect 107473 6712 107485 6715
rect 107344 6684 107485 6712
rect 107344 6672 107350 6684
rect 107473 6681 107485 6684
rect 107519 6712 107531 6715
rect 108040 6712 108068 6743
rect 107519 6684 108068 6712
rect 108500 6712 108528 6820
rect 108577 6817 108589 6851
rect 108623 6848 108635 6851
rect 109494 6848 109500 6860
rect 108623 6820 109500 6848
rect 108623 6817 108635 6820
rect 108577 6811 108635 6817
rect 109494 6808 109500 6820
rect 109552 6808 109558 6860
rect 109604 6820 112576 6848
rect 109604 6712 109632 6820
rect 110325 6783 110383 6789
rect 110325 6780 110337 6783
rect 108500 6684 109632 6712
rect 109696 6752 110337 6780
rect 107519 6681 107531 6684
rect 107473 6675 107531 6681
rect 90910 6604 90916 6656
rect 90968 6604 90974 6656
rect 92750 6604 92756 6656
rect 92808 6604 92814 6656
rect 98362 6604 98368 6656
rect 98420 6604 98426 6656
rect 101214 6604 101220 6656
rect 101272 6604 101278 6656
rect 103698 6604 103704 6656
rect 103756 6644 103762 6656
rect 109696 6653 109724 6752
rect 110325 6749 110337 6752
rect 110371 6749 110383 6783
rect 112257 6783 112315 6789
rect 112257 6780 112269 6783
rect 110325 6743 110383 6749
rect 111536 6752 112269 6780
rect 110874 6672 110880 6724
rect 110932 6672 110938 6724
rect 111536 6656 111564 6752
rect 112257 6749 112269 6752
rect 112303 6749 112315 6783
rect 112257 6743 112315 6749
rect 109681 6647 109739 6653
rect 109681 6644 109693 6647
rect 103756 6616 109693 6644
rect 103756 6604 103762 6616
rect 109681 6613 109693 6616
rect 109727 6613 109739 6647
rect 109681 6607 109739 6613
rect 111518 6604 111524 6656
rect 111576 6604 111582 6656
rect 112548 6644 112576 6820
rect 112806 6808 112812 6860
rect 112864 6808 112870 6860
rect 115385 6851 115443 6857
rect 115385 6817 115397 6851
rect 115431 6848 115443 6851
rect 115431 6820 118694 6848
rect 115431 6817 115443 6820
rect 115385 6811 115443 6817
rect 112714 6740 112720 6792
rect 112772 6780 112778 6792
rect 113358 6780 113364 6792
rect 112772 6752 113364 6780
rect 112772 6740 112778 6752
rect 113358 6740 113364 6752
rect 113416 6780 113422 6792
rect 113637 6783 113695 6789
rect 113637 6780 113649 6783
rect 113416 6752 113649 6780
rect 113416 6740 113422 6752
rect 113637 6749 113649 6752
rect 113683 6749 113695 6783
rect 113637 6743 113695 6749
rect 114646 6740 114652 6792
rect 114704 6780 114710 6792
rect 114833 6783 114891 6789
rect 114833 6780 114845 6783
rect 114704 6752 114845 6780
rect 114704 6740 114710 6752
rect 114833 6749 114845 6752
rect 114879 6749 114891 6783
rect 117409 6783 117467 6789
rect 117409 6780 117421 6783
rect 114833 6743 114891 6749
rect 116688 6752 117421 6780
rect 114186 6672 114192 6724
rect 114244 6672 114250 6724
rect 116688 6656 116716 6752
rect 117409 6749 117421 6752
rect 117455 6749 117467 6783
rect 118666 6780 118694 6820
rect 118786 6808 118792 6860
rect 118844 6848 118850 6860
rect 224954 6848 224960 6860
rect 118844 6820 224960 6848
rect 118844 6808 118850 6820
rect 224954 6808 224960 6820
rect 225012 6808 225018 6860
rect 258350 6808 258356 6860
rect 258408 6808 258414 6860
rect 259549 6851 259607 6857
rect 259549 6817 259561 6851
rect 259595 6848 259607 6851
rect 268378 6848 268384 6860
rect 259595 6820 268384 6848
rect 259595 6817 259607 6820
rect 259549 6811 259607 6817
rect 268378 6808 268384 6820
rect 268436 6808 268442 6860
rect 327534 6808 327540 6860
rect 327592 6848 327598 6860
rect 377030 6848 377036 6860
rect 327592 6820 377036 6848
rect 327592 6808 327598 6820
rect 377030 6808 377036 6820
rect 377088 6808 377094 6860
rect 440970 6808 440976 6860
rect 441028 6848 441034 6860
rect 444742 6848 444748 6860
rect 441028 6820 444748 6848
rect 441028 6808 441034 6820
rect 444742 6808 444748 6820
rect 444800 6808 444806 6860
rect 223206 6780 223212 6792
rect 118666 6752 223212 6780
rect 117409 6743 117467 6749
rect 223206 6740 223212 6752
rect 223264 6740 223270 6792
rect 251913 6783 251971 6789
rect 251913 6749 251925 6783
rect 251959 6780 251971 6783
rect 255225 6783 255283 6789
rect 255225 6780 255237 6783
rect 251959 6752 252600 6780
rect 251959 6749 251971 6752
rect 251913 6743 251971 6749
rect 117961 6715 118019 6721
rect 117961 6681 117973 6715
rect 118007 6712 118019 6715
rect 225414 6712 225420 6724
rect 118007 6684 225420 6712
rect 118007 6681 118019 6684
rect 117961 6675 118019 6681
rect 225414 6672 225420 6684
rect 225472 6672 225478 6724
rect 251358 6672 251364 6724
rect 251416 6672 251422 6724
rect 252572 6656 252600 6752
rect 254596 6752 255237 6780
rect 254596 6656 254624 6752
rect 255225 6749 255237 6752
rect 255271 6749 255283 6783
rect 255225 6743 255283 6749
rect 256326 6740 256332 6792
rect 256384 6780 256390 6792
rect 256605 6783 256663 6789
rect 256605 6780 256617 6783
rect 256384 6752 256617 6780
rect 256384 6740 256390 6752
rect 256605 6749 256617 6752
rect 256651 6749 256663 6783
rect 256605 6743 256663 6749
rect 257522 6740 257528 6792
rect 257580 6780 257586 6792
rect 257801 6783 257859 6789
rect 257801 6780 257813 6783
rect 257580 6752 257813 6780
rect 257580 6740 257586 6752
rect 257801 6749 257813 6752
rect 257847 6749 257859 6783
rect 257801 6743 257859 6749
rect 258994 6740 259000 6792
rect 259052 6740 259058 6792
rect 259914 6740 259920 6792
rect 259972 6780 259978 6792
rect 260193 6783 260251 6789
rect 260193 6780 260205 6783
rect 259972 6752 260205 6780
rect 259972 6740 259978 6752
rect 260193 6749 260205 6752
rect 260239 6749 260251 6783
rect 267642 6780 267648 6792
rect 260193 6743 260251 6749
rect 260668 6752 267648 6780
rect 255777 6715 255835 6721
rect 255777 6681 255789 6715
rect 255823 6681 255835 6715
rect 255777 6675 255835 6681
rect 116026 6644 116032 6656
rect 112548 6616 116032 6644
rect 116026 6604 116032 6616
rect 116084 6604 116090 6656
rect 116670 6604 116676 6656
rect 116728 6604 116734 6656
rect 120261 6647 120319 6653
rect 120261 6613 120273 6647
rect 120307 6644 120319 6647
rect 120442 6644 120448 6656
rect 120307 6616 120448 6644
rect 120307 6613 120319 6616
rect 120261 6607 120319 6613
rect 120442 6604 120448 6616
rect 120500 6604 120506 6656
rect 121457 6647 121515 6653
rect 121457 6613 121469 6647
rect 121503 6644 121515 6647
rect 121638 6644 121644 6656
rect 121503 6616 121644 6644
rect 121503 6613 121515 6616
rect 121457 6607 121515 6613
rect 121638 6604 121644 6616
rect 121696 6604 121702 6656
rect 122098 6604 122104 6656
rect 122156 6644 122162 6656
rect 123386 6644 123392 6656
rect 122156 6616 123392 6644
rect 122156 6604 122162 6616
rect 123386 6604 123392 6616
rect 123444 6604 123450 6656
rect 124030 6604 124036 6656
rect 124088 6644 124094 6656
rect 230474 6644 230480 6656
rect 124088 6616 230480 6644
rect 124088 6604 124094 6616
rect 230474 6604 230480 6616
rect 230532 6604 230538 6656
rect 252554 6604 252560 6656
rect 252612 6604 252618 6656
rect 253934 6604 253940 6656
rect 253992 6604 253998 6656
rect 254578 6604 254584 6656
rect 254636 6604 254642 6656
rect 255792 6644 255820 6675
rect 257154 6672 257160 6724
rect 257212 6672 257218 6724
rect 260668 6644 260696 6752
rect 267642 6740 267648 6752
rect 267700 6740 267706 6792
rect 372798 6740 372804 6792
rect 372856 6780 372862 6792
rect 401962 6780 401968 6792
rect 372856 6752 401968 6780
rect 372856 6740 372862 6752
rect 401962 6740 401968 6752
rect 402020 6740 402026 6792
rect 260745 6715 260803 6721
rect 260745 6681 260757 6715
rect 260791 6712 260803 6715
rect 358814 6712 358820 6724
rect 260791 6684 358820 6712
rect 260791 6681 260803 6684
rect 260745 6675 260803 6681
rect 358814 6672 358820 6684
rect 358872 6672 358878 6724
rect 361574 6672 361580 6724
rect 361632 6712 361638 6724
rect 396074 6712 396080 6724
rect 361632 6684 396080 6712
rect 361632 6672 361638 6684
rect 396074 6672 396080 6684
rect 396132 6672 396138 6724
rect 432046 6672 432052 6724
rect 432104 6712 432110 6724
rect 444006 6712 444012 6724
rect 432104 6684 444012 6712
rect 432104 6672 432110 6684
rect 444006 6672 444012 6684
rect 444064 6672 444070 6724
rect 255792 6616 260696 6644
rect 365622 6604 365628 6656
rect 365680 6644 365686 6656
rect 400306 6644 400312 6656
rect 365680 6616 400312 6644
rect 365680 6604 365686 6616
rect 400306 6604 400312 6616
rect 400364 6604 400370 6656
rect 408494 6604 408500 6656
rect 408552 6644 408558 6656
rect 445018 6644 445024 6656
rect 408552 6616 445024 6644
rect 408552 6604 408558 6616
rect 445018 6604 445024 6616
rect 445076 6604 445082 6656
rect 1104 6554 528816 6576
rect 1104 6502 67574 6554
rect 67626 6502 67638 6554
rect 67690 6502 67702 6554
rect 67754 6502 67766 6554
rect 67818 6502 67830 6554
rect 67882 6502 199502 6554
rect 199554 6502 199566 6554
rect 199618 6502 199630 6554
rect 199682 6502 199694 6554
rect 199746 6502 199758 6554
rect 199810 6502 331430 6554
rect 331482 6502 331494 6554
rect 331546 6502 331558 6554
rect 331610 6502 331622 6554
rect 331674 6502 331686 6554
rect 331738 6502 463358 6554
rect 463410 6502 463422 6554
rect 463474 6502 463486 6554
rect 463538 6502 463550 6554
rect 463602 6502 463614 6554
rect 463666 6502 528816 6554
rect 1104 6480 528816 6502
rect 40402 6400 40408 6452
rect 40460 6440 40466 6452
rect 90910 6440 90916 6452
rect 40460 6412 90916 6440
rect 40460 6400 40466 6412
rect 90910 6400 90916 6412
rect 90968 6400 90974 6452
rect 107286 6440 107292 6452
rect 94516 6412 107292 6440
rect 62114 6332 62120 6384
rect 62172 6372 62178 6384
rect 94516 6372 94544 6412
rect 107286 6400 107292 6412
rect 107344 6400 107350 6452
rect 110984 6412 113312 6440
rect 62172 6344 94544 6372
rect 94608 6344 99512 6372
rect 62172 6332 62178 6344
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 29914 6304 29920 6316
rect 17368 6276 29920 6304
rect 17368 6264 17374 6276
rect 29914 6264 29920 6276
rect 29972 6264 29978 6316
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 42978 6236 42984 6248
rect 12952 6208 42984 6236
rect 12952 6196 12958 6208
rect 42978 6196 42984 6208
rect 43036 6196 43042 6248
rect 94608 6236 94636 6344
rect 99377 6307 99435 6313
rect 99377 6304 99389 6307
rect 84166 6208 94636 6236
rect 98656 6276 99389 6304
rect 1854 6128 1860 6180
rect 1912 6168 1918 6180
rect 46934 6168 46940 6180
rect 1912 6140 46940 6168
rect 1912 6128 1918 6140
rect 46934 6128 46940 6140
rect 46992 6128 46998 6180
rect 68922 6128 68928 6180
rect 68980 6168 68986 6180
rect 84166 6168 84194 6208
rect 98656 6177 98684 6276
rect 99377 6273 99389 6276
rect 99423 6273 99435 6307
rect 99377 6267 99435 6273
rect 99484 6236 99512 6344
rect 99926 6332 99932 6384
rect 99984 6332 99990 6384
rect 101950 6332 101956 6384
rect 102008 6332 102014 6384
rect 106182 6332 106188 6384
rect 106240 6332 106246 6384
rect 110984 6381 111012 6412
rect 107473 6375 107531 6381
rect 107473 6341 107485 6375
rect 107519 6372 107531 6375
rect 110969 6375 111027 6381
rect 107519 6344 109034 6372
rect 107519 6341 107531 6344
rect 107473 6335 107531 6341
rect 100570 6264 100576 6316
rect 100628 6304 100634 6316
rect 101401 6307 101459 6313
rect 101401 6304 101413 6307
rect 100628 6276 101413 6304
rect 100628 6264 100634 6276
rect 101401 6273 101413 6276
rect 101447 6273 101459 6307
rect 101401 6267 101459 6273
rect 102594 6264 102600 6316
rect 102652 6304 102658 6316
rect 103241 6307 103299 6313
rect 103241 6304 103253 6307
rect 102652 6276 103253 6304
rect 102652 6264 102658 6276
rect 103241 6273 103253 6276
rect 103287 6273 103299 6307
rect 105725 6307 105783 6313
rect 105725 6304 105737 6307
rect 103241 6267 103299 6273
rect 105096 6276 105737 6304
rect 103698 6236 103704 6248
rect 99484 6208 103704 6236
rect 103698 6196 103704 6208
rect 103756 6196 103762 6248
rect 103790 6196 103796 6248
rect 103848 6196 103854 6248
rect 98641 6171 98699 6177
rect 98641 6168 98653 6171
rect 68980 6140 84194 6168
rect 89686 6140 98653 6168
rect 68980 6128 68986 6140
rect 42886 6060 42892 6112
rect 42944 6100 42950 6112
rect 89686 6100 89714 6140
rect 98641 6137 98653 6140
rect 98687 6137 98699 6171
rect 98641 6131 98699 6137
rect 105096 6112 105124 6276
rect 105725 6273 105737 6276
rect 105771 6273 105783 6307
rect 105725 6267 105783 6273
rect 106918 6264 106924 6316
rect 106976 6304 106982 6316
rect 108025 6307 108083 6313
rect 108025 6304 108037 6307
rect 106976 6276 108037 6304
rect 106976 6264 106982 6276
rect 108025 6273 108037 6276
rect 108071 6273 108083 6307
rect 108025 6267 108083 6273
rect 109006 6168 109034 6344
rect 110969 6341 110981 6375
rect 111015 6341 111027 6375
rect 113284 6372 113312 6412
rect 113358 6400 113364 6452
rect 113416 6440 113422 6452
rect 122098 6440 122104 6452
rect 113416 6412 122104 6440
rect 113416 6400 113422 6412
rect 122098 6400 122104 6412
rect 122156 6400 122162 6452
rect 131390 6440 131396 6452
rect 122208 6412 131396 6440
rect 122208 6381 122236 6412
rect 131390 6400 131396 6412
rect 131448 6400 131454 6452
rect 257154 6400 257160 6452
rect 257212 6440 257218 6452
rect 262214 6440 262220 6452
rect 257212 6412 262220 6440
rect 257212 6400 257218 6412
rect 262214 6400 262220 6412
rect 262272 6400 262278 6452
rect 362310 6440 362316 6452
rect 263566 6412 362316 6440
rect 122193 6375 122251 6381
rect 113284 6344 122144 6372
rect 110969 6335 111027 6341
rect 109770 6264 109776 6316
rect 109828 6304 109834 6316
rect 110417 6307 110475 6313
rect 110417 6304 110429 6307
rect 109828 6276 110429 6304
rect 109828 6264 109834 6276
rect 110417 6273 110429 6276
rect 110463 6273 110475 6307
rect 110417 6267 110475 6273
rect 111978 6264 111984 6316
rect 112036 6304 112042 6316
rect 112349 6307 112407 6313
rect 112349 6304 112361 6307
rect 112036 6276 112361 6304
rect 112036 6264 112042 6276
rect 112349 6273 112361 6276
rect 112395 6273 112407 6307
rect 112349 6267 112407 6273
rect 112901 6307 112959 6313
rect 112901 6273 112913 6307
rect 112947 6304 112959 6307
rect 113174 6304 113180 6316
rect 112947 6276 113180 6304
rect 112947 6273 112959 6276
rect 112901 6267 112959 6273
rect 113174 6264 113180 6276
rect 113232 6264 113238 6316
rect 113542 6264 113548 6316
rect 113600 6264 113606 6316
rect 113652 6276 114232 6304
rect 109494 6196 109500 6248
rect 109552 6236 109558 6248
rect 113652 6236 113680 6276
rect 109552 6208 113680 6236
rect 109552 6196 109558 6208
rect 114094 6196 114100 6248
rect 114152 6196 114158 6248
rect 114204 6236 114232 6276
rect 117498 6264 117504 6316
rect 117556 6304 117562 6316
rect 118237 6307 118295 6313
rect 118237 6304 118249 6307
rect 117556 6276 118249 6304
rect 117556 6264 117562 6276
rect 118237 6273 118249 6276
rect 118283 6273 118295 6307
rect 118237 6267 118295 6273
rect 120442 6264 120448 6316
rect 120500 6264 120506 6316
rect 120994 6264 121000 6316
rect 121052 6264 121058 6316
rect 121638 6264 121644 6316
rect 121696 6264 121702 6316
rect 122116 6304 122144 6344
rect 122193 6341 122205 6375
rect 122239 6341 122251 6375
rect 122193 6335 122251 6341
rect 124401 6375 124459 6381
rect 124401 6341 124413 6375
rect 124447 6372 124459 6375
rect 231854 6372 231860 6384
rect 124447 6344 231860 6372
rect 124447 6341 124459 6344
rect 124401 6335 124459 6341
rect 231854 6332 231860 6344
rect 231912 6332 231918 6384
rect 261941 6375 261999 6381
rect 261941 6341 261953 6375
rect 261987 6372 261999 6375
rect 263566 6372 263594 6412
rect 362310 6400 362316 6412
rect 362368 6400 362374 6452
rect 367922 6400 367928 6452
rect 367980 6440 367986 6452
rect 397914 6440 397920 6452
rect 367980 6412 397920 6440
rect 367980 6400 367986 6412
rect 397914 6400 397920 6412
rect 397972 6400 397978 6452
rect 398834 6400 398840 6452
rect 398892 6440 398898 6452
rect 440234 6440 440240 6452
rect 398892 6412 440240 6440
rect 398892 6400 398898 6412
rect 440234 6400 440240 6412
rect 440292 6400 440298 6452
rect 261987 6344 263594 6372
rect 266817 6375 266875 6381
rect 261987 6341 261999 6344
rect 261941 6335 261999 6341
rect 266817 6341 266829 6375
rect 266863 6372 266875 6375
rect 368474 6372 368480 6384
rect 266863 6344 368480 6372
rect 266863 6341 266875 6344
rect 266817 6335 266875 6341
rect 368474 6332 368480 6344
rect 368532 6332 368538 6384
rect 369946 6332 369952 6384
rect 370004 6372 370010 6384
rect 399846 6372 399852 6384
rect 370004 6344 399852 6372
rect 370004 6332 370010 6344
rect 399846 6332 399852 6344
rect 399904 6332 399910 6384
rect 400306 6332 400312 6384
rect 400364 6372 400370 6384
rect 441706 6372 441712 6384
rect 400364 6344 441712 6372
rect 400364 6332 400370 6344
rect 441706 6332 441712 6344
rect 441764 6332 441770 6384
rect 442902 6332 442908 6384
rect 442960 6372 442966 6384
rect 445846 6372 445852 6384
rect 442960 6344 445852 6372
rect 442960 6332 442966 6344
rect 445846 6332 445852 6344
rect 445904 6332 445910 6384
rect 123478 6304 123484 6316
rect 122116 6276 123484 6304
rect 123478 6264 123484 6276
rect 123536 6264 123542 6316
rect 123849 6307 123907 6313
rect 123849 6273 123861 6307
rect 123895 6273 123907 6307
rect 123849 6267 123907 6273
rect 117958 6236 117964 6248
rect 114204 6208 117964 6236
rect 117958 6196 117964 6208
rect 118016 6196 118022 6248
rect 118510 6196 118516 6248
rect 118568 6196 118574 6248
rect 123864 6236 123892 6267
rect 125134 6264 125140 6316
rect 125192 6264 125198 6316
rect 125502 6264 125508 6316
rect 125560 6264 125566 6316
rect 126606 6264 126612 6316
rect 126664 6304 126670 6316
rect 127253 6307 127311 6313
rect 127253 6304 127265 6307
rect 126664 6276 127265 6304
rect 126664 6264 126670 6276
rect 127253 6273 127265 6276
rect 127299 6273 127311 6307
rect 127253 6267 127311 6273
rect 127802 6264 127808 6316
rect 127860 6264 127866 6316
rect 128354 6264 128360 6316
rect 128412 6304 128418 6316
rect 128449 6307 128507 6313
rect 128449 6304 128461 6307
rect 128412 6276 128461 6304
rect 128412 6264 128418 6276
rect 128449 6273 128461 6276
rect 128495 6273 128507 6307
rect 128449 6267 128507 6273
rect 131390 6264 131396 6316
rect 131448 6304 131454 6316
rect 229830 6304 229836 6316
rect 131448 6276 229836 6304
rect 131448 6264 131454 6276
rect 229830 6264 229836 6276
rect 229888 6264 229894 6316
rect 260834 6264 260840 6316
rect 260892 6304 260898 6316
rect 261389 6307 261447 6313
rect 261389 6304 261401 6307
rect 260892 6276 261401 6304
rect 260892 6264 260898 6276
rect 261389 6273 261401 6276
rect 261435 6273 261447 6307
rect 261389 6267 261447 6273
rect 262306 6264 262312 6316
rect 262364 6304 262370 6316
rect 262585 6307 262643 6313
rect 262585 6304 262597 6307
rect 262364 6276 262597 6304
rect 262364 6264 262370 6276
rect 262585 6273 262597 6276
rect 262631 6273 262643 6307
rect 262585 6267 262643 6273
rect 264330 6264 264336 6316
rect 264388 6304 264394 6316
rect 264977 6307 265035 6313
rect 264977 6304 264989 6307
rect 264388 6276 264989 6304
rect 264388 6264 264394 6276
rect 264977 6273 264989 6276
rect 265023 6273 265035 6307
rect 264977 6267 265035 6273
rect 265986 6264 265992 6316
rect 266044 6304 266050 6316
rect 266265 6307 266323 6313
rect 266265 6304 266277 6307
rect 266044 6276 266277 6304
rect 266044 6264 266050 6276
rect 266265 6273 266277 6276
rect 266311 6273 266323 6307
rect 367094 6304 367100 6316
rect 266265 6267 266323 6273
rect 269408 6276 367100 6304
rect 123220 6208 123892 6236
rect 129001 6239 129059 6245
rect 123110 6168 123116 6180
rect 109006 6140 123116 6168
rect 123110 6128 123116 6140
rect 123168 6128 123174 6180
rect 123220 6112 123248 6208
rect 129001 6205 129013 6239
rect 129047 6236 129059 6239
rect 236270 6236 236276 6248
rect 129047 6208 236276 6236
rect 129047 6205 129059 6208
rect 129001 6199 129059 6205
rect 236270 6196 236276 6208
rect 236328 6196 236334 6248
rect 262214 6196 262220 6248
rect 262272 6236 262278 6248
rect 262398 6236 262404 6248
rect 262272 6208 262404 6236
rect 262272 6196 262278 6208
rect 262398 6196 262404 6208
rect 262456 6196 262462 6248
rect 263137 6239 263195 6245
rect 263137 6205 263149 6239
rect 263183 6236 263195 6239
rect 265529 6239 265587 6245
rect 263183 6208 263594 6236
rect 263183 6205 263195 6208
rect 263137 6199 263195 6205
rect 124674 6128 124680 6180
rect 124732 6168 124738 6180
rect 231394 6168 231400 6180
rect 124732 6140 231400 6168
rect 124732 6128 124738 6140
rect 231394 6128 231400 6140
rect 231452 6128 231458 6180
rect 263566 6168 263594 6208
rect 265529 6205 265541 6239
rect 265575 6236 265587 6239
rect 269408 6236 269436 6276
rect 367094 6264 367100 6276
rect 367152 6264 367158 6316
rect 378134 6264 378140 6316
rect 378192 6304 378198 6316
rect 442626 6304 442632 6316
rect 378192 6276 442632 6304
rect 378192 6264 378198 6276
rect 442626 6264 442632 6276
rect 442684 6264 442690 6316
rect 464522 6264 464528 6316
rect 464580 6304 464586 6316
rect 482094 6304 482100 6316
rect 464580 6276 482100 6304
rect 464580 6264 464586 6276
rect 482094 6264 482100 6276
rect 482152 6264 482158 6316
rect 364978 6236 364984 6248
rect 265575 6208 269436 6236
rect 273226 6208 364984 6236
rect 265575 6205 265587 6208
rect 265529 6199 265587 6205
rect 273226 6168 273254 6208
rect 364978 6196 364984 6208
rect 365036 6196 365042 6248
rect 381538 6196 381544 6248
rect 381596 6236 381602 6248
rect 440694 6236 440700 6248
rect 381596 6208 440700 6236
rect 381596 6196 381602 6208
rect 440694 6196 440700 6208
rect 440752 6196 440758 6248
rect 459554 6196 459560 6248
rect 459612 6236 459618 6248
rect 480254 6236 480260 6248
rect 459612 6208 480260 6236
rect 459612 6196 459618 6208
rect 480254 6196 480260 6208
rect 480312 6196 480318 6248
rect 263566 6140 273254 6168
rect 369854 6128 369860 6180
rect 369912 6168 369918 6180
rect 441614 6168 441620 6180
rect 369912 6140 441620 6168
rect 369912 6128 369918 6140
rect 441614 6128 441620 6140
rect 441672 6128 441678 6180
rect 445662 6128 445668 6180
rect 445720 6168 445726 6180
rect 481266 6168 481272 6180
rect 445720 6140 481272 6168
rect 445720 6128 445726 6140
rect 481266 6128 481272 6140
rect 481324 6128 481330 6180
rect 42944 6072 89714 6100
rect 42944 6060 42950 6072
rect 94314 6060 94320 6112
rect 94372 6060 94378 6112
rect 96709 6103 96767 6109
rect 96709 6069 96721 6103
rect 96755 6100 96767 6103
rect 96798 6100 96804 6112
rect 96755 6072 96804 6100
rect 96755 6069 96767 6072
rect 96709 6063 96767 6069
rect 96798 6060 96804 6072
rect 96856 6060 96862 6112
rect 99558 6060 99564 6112
rect 99616 6100 99622 6112
rect 100570 6100 100576 6112
rect 99616 6072 100576 6100
rect 99616 6060 99622 6072
rect 100570 6060 100576 6072
rect 100628 6100 100634 6112
rect 100757 6103 100815 6109
rect 100757 6100 100769 6103
rect 100628 6072 100769 6100
rect 100628 6060 100634 6072
rect 100757 6069 100769 6072
rect 100803 6069 100815 6103
rect 100757 6063 100815 6069
rect 102594 6060 102600 6112
rect 102652 6060 102658 6112
rect 104434 6060 104440 6112
rect 104492 6060 104498 6112
rect 105078 6060 105084 6112
rect 105136 6060 105142 6112
rect 109770 6060 109776 6112
rect 109828 6060 109834 6112
rect 111797 6103 111855 6109
rect 111797 6069 111809 6103
rect 111843 6100 111855 6103
rect 111978 6100 111984 6112
rect 111843 6072 111984 6100
rect 111843 6069 111855 6072
rect 111797 6063 111855 6069
rect 111978 6060 111984 6072
rect 112036 6060 112042 6112
rect 114646 6060 114652 6112
rect 114704 6100 114710 6112
rect 114741 6103 114799 6109
rect 114741 6100 114753 6103
rect 114704 6072 114753 6100
rect 114704 6060 114710 6072
rect 114741 6069 114753 6072
rect 114787 6069 114799 6103
rect 114741 6063 114799 6069
rect 117498 6060 117504 6112
rect 117556 6100 117562 6112
rect 117593 6103 117651 6109
rect 117593 6100 117605 6103
rect 117556 6072 117605 6100
rect 117556 6060 117562 6072
rect 117593 6069 117605 6072
rect 117639 6069 117651 6103
rect 117593 6063 117651 6069
rect 123202 6060 123208 6112
rect 123260 6060 123266 6112
rect 126606 6060 126612 6112
rect 126664 6060 126670 6112
rect 131669 6103 131727 6109
rect 131669 6069 131681 6103
rect 131715 6100 131727 6103
rect 131758 6100 131764 6112
rect 131715 6072 131764 6100
rect 131715 6069 131727 6072
rect 131669 6063 131727 6069
rect 131758 6060 131764 6072
rect 131816 6060 131822 6112
rect 134426 6060 134432 6112
rect 134484 6100 134490 6112
rect 241606 6100 241612 6112
rect 134484 6072 241612 6100
rect 134484 6060 134490 6072
rect 241606 6060 241612 6072
rect 241664 6060 241670 6112
rect 256326 6060 256332 6112
rect 256384 6060 256390 6112
rect 257522 6060 257528 6112
rect 257580 6060 257586 6112
rect 258994 6060 259000 6112
rect 259052 6060 259058 6112
rect 259914 6060 259920 6112
rect 259972 6060 259978 6112
rect 260834 6060 260840 6112
rect 260892 6060 260898 6112
rect 264330 6060 264336 6112
rect 264388 6060 264394 6112
rect 1104 6010 528816 6032
rect 1104 5958 66914 6010
rect 66966 5958 66978 6010
rect 67030 5958 67042 6010
rect 67094 5958 67106 6010
rect 67158 5958 67170 6010
rect 67222 5958 198842 6010
rect 198894 5958 198906 6010
rect 198958 5958 198970 6010
rect 199022 5958 199034 6010
rect 199086 5958 199098 6010
rect 199150 5958 330770 6010
rect 330822 5958 330834 6010
rect 330886 5958 330898 6010
rect 330950 5958 330962 6010
rect 331014 5958 331026 6010
rect 331078 5958 462698 6010
rect 462750 5958 462762 6010
rect 462814 5958 462826 6010
rect 462878 5958 462890 6010
rect 462942 5958 462954 6010
rect 463006 5958 528816 6010
rect 1104 5936 528816 5958
rect 48774 5856 48780 5908
rect 48832 5896 48838 5908
rect 102594 5896 102600 5908
rect 48832 5868 102600 5896
rect 48832 5856 48838 5868
rect 102594 5856 102600 5868
rect 102652 5856 102658 5908
rect 111518 5896 111524 5908
rect 103486 5868 111524 5896
rect 75914 5788 75920 5840
rect 75972 5828 75978 5840
rect 103486 5828 103514 5868
rect 111518 5856 111524 5868
rect 111576 5856 111582 5908
rect 114094 5856 114100 5908
rect 114152 5896 114158 5908
rect 123294 5896 123300 5908
rect 114152 5868 123300 5896
rect 114152 5856 114158 5868
rect 123294 5856 123300 5868
rect 123352 5856 123358 5908
rect 127342 5856 127348 5908
rect 127400 5896 127406 5908
rect 149698 5896 149704 5908
rect 127400 5868 135760 5896
rect 127400 5856 127406 5868
rect 75972 5800 103514 5828
rect 75972 5788 75978 5800
rect 103790 5788 103796 5840
rect 103848 5828 103854 5840
rect 103848 5800 109034 5828
rect 103848 5788 103854 5800
rect 19886 5720 19892 5772
rect 19944 5760 19950 5772
rect 98362 5760 98368 5772
rect 19944 5732 98368 5760
rect 19944 5720 19950 5732
rect 98362 5720 98368 5732
rect 98420 5720 98426 5772
rect 107562 5720 107568 5772
rect 107620 5720 107626 5772
rect 109006 5760 109034 5800
rect 110874 5788 110880 5840
rect 110932 5828 110938 5840
rect 120166 5828 120172 5840
rect 110932 5800 120172 5828
rect 110932 5788 110938 5800
rect 120166 5788 120172 5800
rect 120224 5788 120230 5840
rect 121288 5800 125594 5828
rect 115382 5760 115388 5772
rect 109006 5732 115388 5760
rect 115382 5720 115388 5732
rect 115440 5720 115446 5772
rect 121288 5769 121316 5800
rect 116673 5763 116731 5769
rect 116673 5729 116685 5763
rect 116719 5760 116731 5763
rect 121273 5763 121331 5769
rect 116719 5732 120028 5760
rect 116719 5729 116731 5732
rect 116673 5723 116731 5729
rect 98638 5652 98644 5704
rect 98696 5692 98702 5704
rect 106369 5695 106427 5701
rect 106369 5692 106381 5695
rect 98696 5664 106381 5692
rect 98696 5652 98702 5664
rect 106369 5661 106381 5664
rect 106415 5692 106427 5695
rect 107105 5695 107163 5701
rect 107105 5692 107117 5695
rect 106415 5664 107117 5692
rect 106415 5661 106427 5664
rect 106369 5655 106427 5661
rect 107105 5661 107117 5664
rect 107151 5661 107163 5695
rect 109313 5695 109371 5701
rect 109313 5692 109325 5695
rect 107105 5655 107163 5661
rect 108684 5664 109325 5692
rect 47394 5584 47400 5636
rect 47452 5624 47458 5636
rect 106918 5624 106924 5636
rect 47452 5596 106924 5624
rect 47452 5584 47458 5596
rect 106918 5584 106924 5596
rect 106976 5584 106982 5636
rect 56502 5516 56508 5568
rect 56560 5556 56566 5568
rect 105078 5556 105084 5568
rect 56560 5528 105084 5556
rect 56560 5516 56566 5528
rect 105078 5516 105084 5528
rect 105136 5516 105142 5568
rect 107654 5516 107660 5568
rect 107712 5556 107718 5568
rect 108684 5565 108712 5664
rect 109313 5661 109325 5664
rect 109359 5661 109371 5695
rect 109313 5655 109371 5661
rect 109862 5652 109868 5704
rect 109920 5652 109926 5704
rect 116121 5695 116179 5701
rect 116121 5692 116133 5695
rect 115492 5664 116133 5692
rect 115492 5568 115520 5664
rect 116121 5661 116133 5664
rect 116167 5661 116179 5695
rect 116121 5655 116179 5661
rect 117130 5652 117136 5704
rect 117188 5692 117194 5704
rect 117409 5695 117467 5701
rect 117409 5692 117421 5695
rect 117188 5664 117421 5692
rect 117188 5652 117194 5664
rect 117409 5661 117421 5664
rect 117455 5661 117467 5695
rect 117409 5655 117467 5661
rect 117961 5695 118019 5701
rect 117961 5661 117973 5695
rect 118007 5692 118019 5695
rect 118786 5692 118792 5704
rect 118007 5664 118792 5692
rect 118007 5661 118019 5664
rect 117961 5655 118019 5661
rect 118786 5652 118792 5664
rect 118844 5652 118850 5704
rect 119525 5695 119583 5701
rect 119525 5692 119537 5695
rect 118896 5664 119537 5692
rect 118896 5568 118924 5664
rect 119525 5661 119537 5664
rect 119571 5661 119583 5695
rect 119525 5655 119583 5661
rect 108669 5559 108727 5565
rect 108669 5556 108681 5559
rect 107712 5528 108681 5556
rect 107712 5516 107718 5528
rect 108669 5525 108681 5528
rect 108715 5525 108727 5559
rect 108669 5519 108727 5525
rect 108758 5516 108764 5568
rect 108816 5556 108822 5568
rect 113269 5559 113327 5565
rect 113269 5556 113281 5559
rect 108816 5528 113281 5556
rect 108816 5516 108822 5528
rect 113269 5525 113281 5528
rect 113315 5556 113327 5559
rect 113542 5556 113548 5568
rect 113315 5528 113548 5556
rect 113315 5525 113327 5528
rect 113269 5519 113327 5525
rect 113542 5516 113548 5528
rect 113600 5516 113606 5568
rect 115474 5516 115480 5568
rect 115532 5516 115538 5568
rect 118878 5516 118884 5568
rect 118936 5516 118942 5568
rect 120000 5556 120028 5732
rect 121273 5729 121285 5763
rect 121319 5729 121331 5763
rect 121273 5723 121331 5729
rect 124232 5732 124444 5760
rect 120718 5652 120724 5704
rect 120776 5652 120782 5704
rect 122834 5652 122840 5704
rect 122892 5692 122898 5704
rect 122929 5695 122987 5701
rect 122929 5692 122941 5695
rect 122892 5664 122941 5692
rect 122892 5652 122898 5664
rect 122929 5661 122941 5664
rect 122975 5661 122987 5695
rect 122929 5655 122987 5661
rect 123481 5695 123539 5701
rect 123481 5661 123493 5695
rect 123527 5692 123539 5695
rect 124030 5692 124036 5704
rect 123527 5664 124036 5692
rect 123527 5661 123539 5664
rect 123481 5655 123539 5661
rect 124030 5652 124036 5664
rect 124088 5652 124094 5704
rect 124122 5652 124128 5704
rect 124180 5652 124186 5704
rect 120077 5627 120135 5633
rect 120077 5593 120089 5627
rect 120123 5624 120135 5627
rect 124232 5624 124260 5732
rect 124416 5692 124444 5732
rect 124674 5720 124680 5772
rect 124732 5720 124738 5772
rect 125566 5760 125594 5800
rect 130396 5800 135484 5828
rect 130396 5760 130424 5800
rect 125566 5732 130424 5760
rect 130856 5732 134564 5760
rect 127342 5692 127348 5704
rect 124416 5664 127348 5692
rect 127342 5652 127348 5664
rect 127400 5652 127406 5704
rect 130654 5652 130660 5704
rect 130712 5652 130718 5704
rect 130856 5624 130884 5732
rect 130930 5652 130936 5704
rect 130988 5652 130994 5704
rect 131758 5652 131764 5704
rect 131816 5652 131822 5704
rect 132034 5652 132040 5704
rect 132092 5652 132098 5704
rect 134153 5695 134211 5701
rect 134153 5692 134165 5695
rect 133616 5664 134165 5692
rect 120123 5596 124260 5624
rect 124324 5596 130884 5624
rect 120123 5593 120135 5596
rect 120077 5587 120135 5593
rect 124324 5556 124352 5596
rect 133616 5568 133644 5664
rect 134153 5661 134165 5664
rect 134199 5661 134211 5695
rect 134153 5655 134211 5661
rect 134426 5652 134432 5704
rect 134484 5652 134490 5704
rect 134536 5624 134564 5732
rect 135257 5695 135315 5701
rect 135257 5661 135269 5695
rect 135303 5692 135315 5695
rect 135346 5692 135352 5704
rect 135303 5664 135352 5692
rect 135303 5661 135315 5664
rect 135257 5655 135315 5661
rect 135346 5652 135352 5664
rect 135404 5652 135410 5704
rect 135456 5692 135484 5800
rect 135530 5720 135536 5772
rect 135588 5720 135594 5772
rect 135732 5760 135760 5868
rect 137986 5868 149704 5896
rect 137986 5760 138014 5868
rect 149698 5856 149704 5868
rect 149756 5856 149762 5908
rect 372522 5896 372528 5908
rect 269132 5868 372528 5896
rect 228082 5828 228088 5840
rect 135732 5732 138014 5760
rect 138216 5800 144914 5828
rect 138216 5692 138244 5800
rect 144886 5760 144914 5800
rect 147784 5800 228088 5828
rect 147784 5760 147812 5800
rect 228082 5788 228088 5800
rect 228140 5788 228146 5840
rect 144886 5732 147812 5760
rect 149698 5720 149704 5772
rect 149756 5760 149762 5772
rect 226978 5760 226984 5772
rect 149756 5732 226984 5760
rect 149756 5720 149762 5732
rect 226978 5720 226984 5732
rect 227036 5720 227042 5772
rect 269132 5769 269160 5868
rect 372522 5856 372528 5868
rect 372580 5856 372586 5908
rect 365714 5828 365720 5840
rect 269316 5800 365720 5828
rect 264333 5763 264391 5769
rect 264333 5729 264345 5763
rect 264379 5760 264391 5763
rect 269117 5763 269175 5769
rect 264379 5732 269068 5760
rect 264379 5729 264391 5732
rect 264333 5723 264391 5729
rect 135456 5664 138244 5692
rect 138290 5652 138296 5704
rect 138348 5692 138354 5704
rect 138753 5695 138811 5701
rect 138753 5692 138765 5695
rect 138348 5664 138765 5692
rect 138348 5652 138354 5664
rect 138753 5661 138765 5664
rect 138799 5661 138811 5695
rect 138753 5655 138811 5661
rect 138952 5664 147674 5692
rect 138952 5624 138980 5664
rect 134536 5596 138980 5624
rect 139026 5584 139032 5636
rect 139084 5584 139090 5636
rect 147646 5624 147674 5664
rect 263134 5652 263140 5704
rect 263192 5692 263198 5704
rect 263781 5695 263839 5701
rect 263781 5692 263793 5695
rect 263192 5664 263793 5692
rect 263192 5652 263198 5664
rect 263781 5661 263793 5664
rect 263827 5661 263839 5695
rect 266817 5695 266875 5701
rect 266817 5692 266829 5695
rect 263781 5655 263839 5661
rect 264256 5664 266829 5692
rect 223758 5624 223764 5636
rect 147646 5596 223764 5624
rect 223758 5584 223764 5596
rect 223816 5584 223822 5636
rect 252646 5584 252652 5636
rect 252704 5624 252710 5636
rect 264256 5624 264284 5664
rect 266817 5661 266829 5664
rect 266863 5692 266875 5695
rect 267461 5695 267519 5701
rect 267461 5692 267473 5695
rect 266863 5664 267473 5692
rect 266863 5661 266875 5664
rect 266817 5655 266875 5661
rect 267461 5661 267473 5664
rect 267507 5661 267519 5695
rect 267461 5655 267519 5661
rect 268378 5652 268384 5704
rect 268436 5692 268442 5704
rect 268657 5695 268715 5701
rect 268657 5692 268669 5695
rect 268436 5664 268669 5692
rect 268436 5652 268442 5664
rect 268657 5661 268669 5664
rect 268703 5661 268715 5695
rect 269040 5692 269068 5732
rect 269117 5729 269129 5763
rect 269163 5729 269175 5763
rect 269117 5723 269175 5729
rect 269316 5692 269344 5800
rect 365714 5788 365720 5800
rect 365772 5788 365778 5840
rect 370774 5760 370780 5772
rect 270420 5732 370780 5760
rect 269040 5664 269344 5692
rect 268657 5655 268715 5661
rect 269666 5652 269672 5704
rect 269724 5692 269730 5704
rect 269945 5695 270003 5701
rect 269945 5692 269957 5695
rect 269724 5664 269957 5692
rect 269724 5652 269730 5664
rect 269945 5661 269957 5664
rect 269991 5661 270003 5695
rect 269945 5655 270003 5661
rect 252704 5596 264284 5624
rect 268013 5627 268071 5633
rect 252704 5584 252710 5596
rect 268013 5593 268025 5627
rect 268059 5624 268071 5627
rect 270420 5624 270448 5732
rect 370774 5720 370780 5732
rect 370832 5720 370838 5772
rect 268059 5596 270448 5624
rect 270497 5627 270555 5633
rect 268059 5593 268071 5596
rect 268013 5587 268071 5593
rect 270497 5593 270509 5627
rect 270543 5624 270555 5627
rect 373442 5624 373448 5636
rect 270543 5596 373448 5624
rect 270543 5593 270555 5596
rect 270497 5587 270555 5593
rect 373442 5584 373448 5596
rect 373500 5584 373506 5636
rect 120000 5528 124352 5556
rect 128170 5516 128176 5568
rect 128228 5516 128234 5568
rect 130102 5516 130108 5568
rect 130160 5556 130166 5568
rect 130654 5556 130660 5568
rect 130160 5528 130660 5556
rect 130160 5516 130166 5528
rect 130654 5516 130660 5528
rect 130712 5516 130718 5568
rect 133598 5516 133604 5568
rect 133656 5516 133662 5568
rect 138198 5516 138204 5568
rect 138256 5516 138262 5568
rect 141694 5516 141700 5568
rect 141752 5556 141758 5568
rect 141973 5559 142031 5565
rect 141973 5556 141985 5559
rect 141752 5528 141985 5556
rect 141752 5516 141758 5528
rect 141973 5525 141985 5528
rect 142019 5525 142031 5559
rect 141973 5519 142031 5525
rect 262306 5516 262312 5568
rect 262364 5516 262370 5568
rect 263134 5516 263140 5568
rect 263192 5516 263198 5568
rect 265986 5516 265992 5568
rect 266044 5516 266050 5568
rect 1104 5466 528816 5488
rect 1104 5414 67574 5466
rect 67626 5414 67638 5466
rect 67690 5414 67702 5466
rect 67754 5414 67766 5466
rect 67818 5414 67830 5466
rect 67882 5414 199502 5466
rect 199554 5414 199566 5466
rect 199618 5414 199630 5466
rect 199682 5414 199694 5466
rect 199746 5414 199758 5466
rect 199810 5414 331430 5466
rect 331482 5414 331494 5466
rect 331546 5414 331558 5466
rect 331610 5414 331622 5466
rect 331674 5414 331686 5466
rect 331738 5414 463358 5466
rect 463410 5414 463422 5466
rect 463474 5414 463486 5466
rect 463538 5414 463550 5466
rect 463602 5414 463614 5466
rect 463666 5414 528816 5466
rect 1104 5392 528816 5414
rect 18046 5312 18052 5364
rect 18104 5352 18110 5364
rect 96614 5352 96620 5364
rect 18104 5324 96620 5352
rect 18104 5312 18110 5324
rect 96614 5312 96620 5324
rect 96672 5312 96678 5364
rect 241146 5352 241152 5364
rect 118666 5324 134472 5352
rect 9582 5244 9588 5296
rect 9640 5284 9646 5296
rect 92382 5284 92388 5296
rect 9640 5256 92388 5284
rect 9640 5244 9646 5256
rect 92382 5244 92388 5256
rect 92440 5244 92446 5296
rect 5166 5176 5172 5228
rect 5224 5216 5230 5228
rect 94498 5216 94504 5228
rect 5224 5188 94504 5216
rect 5224 5176 5230 5188
rect 94498 5176 94504 5188
rect 94556 5176 94562 5228
rect 115106 5176 115112 5228
rect 115164 5216 115170 5228
rect 118666 5216 118694 5324
rect 126885 5287 126943 5293
rect 126885 5253 126897 5287
rect 126931 5284 126943 5287
rect 126931 5256 133644 5284
rect 126931 5253 126943 5256
rect 126885 5247 126943 5253
rect 115164 5188 118694 5216
rect 115164 5176 115170 5188
rect 125686 5176 125692 5228
rect 125744 5216 125750 5228
rect 126333 5219 126391 5225
rect 126333 5216 126345 5219
rect 125744 5188 126345 5216
rect 125744 5176 125750 5188
rect 126333 5185 126345 5188
rect 126379 5185 126391 5219
rect 126333 5179 126391 5185
rect 127529 5219 127587 5225
rect 127529 5185 127541 5219
rect 127575 5216 127587 5219
rect 127618 5216 127624 5228
rect 127575 5188 127624 5216
rect 127575 5185 127587 5188
rect 127529 5179 127587 5185
rect 127618 5176 127624 5188
rect 127676 5176 127682 5228
rect 130289 5219 130347 5225
rect 130289 5216 130301 5219
rect 129568 5188 130301 5216
rect 6822 5108 6828 5160
rect 6880 5148 6886 5160
rect 78674 5148 78680 5160
rect 6880 5120 78680 5148
rect 6880 5108 6886 5120
rect 78674 5108 78680 5120
rect 78732 5108 78738 5160
rect 82814 5108 82820 5160
rect 82872 5148 82878 5160
rect 117130 5148 117136 5160
rect 82872 5120 117136 5148
rect 82872 5108 82878 5120
rect 117130 5108 117136 5120
rect 117188 5108 117194 5160
rect 128078 5108 128084 5160
rect 128136 5108 128142 5160
rect 68830 5040 68836 5092
rect 68888 5080 68894 5092
rect 68888 5052 70394 5080
rect 68888 5040 68894 5052
rect 45646 4972 45652 5024
rect 45704 5012 45710 5024
rect 68922 5012 68928 5024
rect 45704 4984 68928 5012
rect 45704 4972 45710 4984
rect 68922 4972 68928 4984
rect 68980 4972 68986 5024
rect 70366 5012 70394 5052
rect 76558 5040 76564 5092
rect 76616 5080 76622 5092
rect 123849 5083 123907 5089
rect 123849 5080 123861 5083
rect 76616 5052 123861 5080
rect 76616 5040 76622 5052
rect 123849 5049 123861 5052
rect 123895 5080 123907 5083
rect 124122 5080 124128 5092
rect 123895 5052 124128 5080
rect 123895 5049 123907 5052
rect 123849 5043 123907 5049
rect 124122 5040 124128 5052
rect 124180 5040 124186 5092
rect 129568 5024 129596 5188
rect 130289 5185 130301 5188
rect 130335 5185 130347 5219
rect 130289 5179 130347 5185
rect 131206 5176 131212 5228
rect 131264 5216 131270 5228
rect 131393 5219 131451 5225
rect 131393 5216 131405 5219
rect 131264 5188 131405 5216
rect 131264 5176 131270 5188
rect 131393 5185 131405 5188
rect 131439 5185 131451 5219
rect 131393 5179 131451 5185
rect 132678 5176 132684 5228
rect 132736 5216 132742 5228
rect 133233 5219 133291 5225
rect 133233 5216 133245 5219
rect 132736 5188 133245 5216
rect 132736 5176 132742 5188
rect 133233 5185 133245 5188
rect 133279 5185 133291 5219
rect 133233 5179 133291 5185
rect 130838 5108 130844 5160
rect 130896 5108 130902 5160
rect 131669 5151 131727 5157
rect 131669 5117 131681 5151
rect 131715 5117 131727 5151
rect 131669 5111 131727 5117
rect 131684 5080 131712 5111
rect 133506 5108 133512 5160
rect 133564 5108 133570 5160
rect 133616 5148 133644 5256
rect 134334 5176 134340 5228
rect 134392 5176 134398 5228
rect 134444 5216 134472 5324
rect 134628 5324 241152 5352
rect 134628 5293 134656 5324
rect 241146 5312 241152 5324
rect 241204 5312 241210 5364
rect 252554 5312 252560 5364
rect 252612 5352 252618 5364
rect 360746 5352 360752 5364
rect 252612 5324 360752 5352
rect 252612 5312 252618 5324
rect 360746 5312 360752 5324
rect 360804 5312 360810 5364
rect 389174 5312 389180 5364
rect 389232 5352 389238 5364
rect 403618 5352 403624 5364
rect 389232 5324 403624 5352
rect 389232 5312 389238 5324
rect 403618 5312 403624 5324
rect 403676 5312 403682 5364
rect 426986 5312 426992 5364
rect 427044 5352 427050 5364
rect 443086 5352 443092 5364
rect 427044 5324 443092 5352
rect 427044 5312 427050 5324
rect 443086 5312 443092 5324
rect 443144 5312 443150 5364
rect 443730 5312 443736 5364
rect 443788 5352 443794 5364
rect 446122 5352 446128 5364
rect 443788 5324 446128 5352
rect 443788 5312 443794 5324
rect 446122 5312 446128 5324
rect 446180 5312 446186 5364
rect 477494 5312 477500 5364
rect 477552 5352 477558 5364
rect 481634 5352 481640 5364
rect 477552 5324 481640 5352
rect 477552 5312 477558 5324
rect 481634 5312 481640 5324
rect 481692 5312 481698 5364
rect 134613 5287 134671 5293
rect 134613 5253 134625 5287
rect 134659 5253 134671 5287
rect 134613 5247 134671 5253
rect 137002 5244 137008 5296
rect 137060 5284 137066 5296
rect 137060 5256 137600 5284
rect 137060 5244 137066 5256
rect 137094 5216 137100 5228
rect 134444 5188 137100 5216
rect 137094 5176 137100 5188
rect 137152 5176 137158 5228
rect 137572 5225 137600 5256
rect 137986 5256 144960 5284
rect 137557 5219 137615 5225
rect 137557 5185 137569 5219
rect 137603 5185 137615 5219
rect 137986 5216 138014 5256
rect 137557 5179 137615 5185
rect 137664 5188 138014 5216
rect 137664 5148 137692 5188
rect 140498 5176 140504 5228
rect 140556 5216 140562 5228
rect 141053 5219 141111 5225
rect 141053 5216 141065 5219
rect 140556 5188 141065 5216
rect 140556 5176 140562 5188
rect 141053 5185 141065 5188
rect 141099 5185 141111 5219
rect 141053 5179 141111 5185
rect 141326 5176 141332 5228
rect 141384 5176 141390 5228
rect 141694 5176 141700 5228
rect 141752 5216 141758 5228
rect 142157 5219 142215 5225
rect 142157 5216 142169 5219
rect 141752 5188 142169 5216
rect 141752 5176 141758 5188
rect 142157 5185 142169 5188
rect 142203 5185 142215 5219
rect 142157 5179 142215 5185
rect 144546 5176 144552 5228
rect 144604 5176 144610 5228
rect 133616 5120 137692 5148
rect 137830 5108 137836 5160
rect 137888 5108 137894 5160
rect 142430 5108 142436 5160
rect 142488 5108 142494 5160
rect 144822 5108 144828 5160
rect 144880 5108 144886 5160
rect 144932 5148 144960 5256
rect 145834 5244 145840 5296
rect 145892 5284 145898 5296
rect 236914 5284 236920 5296
rect 145892 5256 236920 5284
rect 145892 5244 145898 5256
rect 236914 5244 236920 5256
rect 236972 5244 236978 5296
rect 291102 5244 291108 5296
rect 291160 5284 291166 5296
rect 391934 5284 391940 5296
rect 291160 5256 391940 5284
rect 291160 5244 291166 5256
rect 391934 5244 391940 5256
rect 391992 5244 391998 5296
rect 417050 5244 417056 5296
rect 417108 5284 417114 5296
rect 443178 5284 443184 5296
rect 417108 5256 443184 5284
rect 417108 5244 417114 5256
rect 443178 5244 443184 5256
rect 443236 5244 443242 5296
rect 145466 5176 145472 5228
rect 145524 5216 145530 5228
rect 145653 5219 145711 5225
rect 145653 5216 145665 5219
rect 145524 5188 145665 5216
rect 145524 5176 145530 5188
rect 145653 5185 145665 5188
rect 145699 5185 145711 5219
rect 145653 5179 145711 5185
rect 145926 5176 145932 5228
rect 145984 5176 145990 5228
rect 148042 5176 148048 5228
rect 148100 5176 148106 5228
rect 148152 5188 151814 5216
rect 148152 5148 148180 5188
rect 144932 5120 148180 5148
rect 148321 5151 148379 5157
rect 148321 5117 148333 5151
rect 148367 5148 148379 5151
rect 148962 5148 148968 5160
rect 148367 5120 148968 5148
rect 148367 5117 148379 5120
rect 148321 5111 148379 5117
rect 148962 5108 148968 5120
rect 149020 5108 149026 5160
rect 151786 5148 151814 5188
rect 270586 5176 270592 5228
rect 270644 5216 270650 5228
rect 271141 5219 271199 5225
rect 271141 5216 271153 5219
rect 270644 5188 271153 5216
rect 270644 5176 270650 5188
rect 271141 5185 271153 5188
rect 271187 5185 271199 5219
rect 271141 5179 271199 5185
rect 285950 5176 285956 5228
rect 286008 5216 286014 5228
rect 390554 5216 390560 5228
rect 286008 5188 390560 5216
rect 286008 5176 286014 5188
rect 390554 5176 390560 5188
rect 390612 5176 390618 5228
rect 403986 5176 403992 5228
rect 404044 5216 404050 5228
rect 442994 5216 443000 5228
rect 404044 5188 443000 5216
rect 404044 5176 404050 5188
rect 442994 5176 443000 5188
rect 443052 5176 443058 5228
rect 233602 5148 233608 5160
rect 151786 5120 233608 5148
rect 233602 5108 233608 5120
rect 233660 5108 233666 5160
rect 271690 5108 271696 5160
rect 271748 5108 271754 5160
rect 288526 5108 288532 5160
rect 288584 5148 288590 5160
rect 391382 5148 391388 5160
rect 288584 5120 391388 5148
rect 288584 5108 288590 5120
rect 391382 5108 391388 5120
rect 391440 5108 391446 5160
rect 400398 5108 400404 5160
rect 400456 5148 400462 5160
rect 441798 5148 441804 5160
rect 400456 5120 441804 5148
rect 400456 5108 400462 5120
rect 441798 5108 441804 5120
rect 441856 5108 441862 5160
rect 475286 5108 475292 5160
rect 475344 5148 475350 5160
rect 480714 5148 480720 5160
rect 475344 5120 480720 5148
rect 475344 5108 475350 5120
rect 480714 5108 480720 5120
rect 480772 5108 480778 5160
rect 481726 5108 481732 5160
rect 481784 5148 481790 5160
rect 482002 5148 482008 5160
rect 481784 5120 482008 5148
rect 481784 5108 481790 5120
rect 482002 5108 482008 5120
rect 482060 5108 482066 5160
rect 237926 5080 237932 5092
rect 131684 5052 237932 5080
rect 237926 5040 237932 5052
rect 237984 5040 237990 5092
rect 283374 5040 283380 5092
rect 283432 5080 283438 5092
rect 390646 5080 390652 5092
rect 283432 5052 390652 5080
rect 283432 5040 283438 5052
rect 390646 5040 390652 5052
rect 390704 5040 390710 5092
rect 404354 5040 404360 5092
rect 404412 5080 404418 5092
rect 439130 5080 439136 5092
rect 404412 5052 439136 5080
rect 404412 5040 404418 5052
rect 439130 5040 439136 5052
rect 439188 5040 439194 5092
rect 440326 5080 440332 5092
rect 439240 5052 440332 5080
rect 120445 5015 120503 5021
rect 120445 5012 120457 5015
rect 70366 4984 120457 5012
rect 120445 4981 120457 4984
rect 120491 5012 120503 5015
rect 120718 5012 120724 5024
rect 120491 4984 120724 5012
rect 120491 4981 120503 4984
rect 120445 4975 120503 4981
rect 120718 4972 120724 4984
rect 120776 4972 120782 5024
rect 122745 5015 122803 5021
rect 122745 4981 122757 5015
rect 122791 5012 122803 5015
rect 122834 5012 122840 5024
rect 122791 4984 122840 5012
rect 122791 4981 122803 4984
rect 122745 4975 122803 4981
rect 122834 4972 122840 4984
rect 122892 4972 122898 5024
rect 125686 4972 125692 5024
rect 125744 4972 125750 5024
rect 129550 4972 129556 5024
rect 129608 4972 129614 5024
rect 132678 4972 132684 5024
rect 132736 4972 132742 5024
rect 135346 4972 135352 5024
rect 135404 4972 135410 5024
rect 137002 4972 137008 5024
rect 137060 4972 137066 5024
rect 137094 4972 137100 5024
rect 137152 5012 137158 5024
rect 140498 5012 140504 5024
rect 137152 4984 140504 5012
rect 137152 4972 137158 4984
rect 140498 4972 140504 4984
rect 140556 4972 140562 5024
rect 140682 4972 140688 5024
rect 140740 5012 140746 5024
rect 143997 5015 144055 5021
rect 143997 5012 144009 5015
rect 140740 4984 144009 5012
rect 140740 4972 140746 4984
rect 143997 4981 144009 4984
rect 144043 5012 144055 5015
rect 144546 5012 144552 5024
rect 144043 4984 144552 5012
rect 144043 4981 144055 4984
rect 143997 4975 144055 4981
rect 144546 4972 144552 4984
rect 144604 4972 144610 5024
rect 144638 4972 144644 5024
rect 144696 5012 144702 5024
rect 147493 5015 147551 5021
rect 147493 5012 147505 5015
rect 144696 4984 147505 5012
rect 144696 4972 144702 4984
rect 147493 4981 147505 4984
rect 147539 5012 147551 5015
rect 148042 5012 148048 5024
rect 147539 4984 148048 5012
rect 147539 4981 147551 4984
rect 147493 4975 147551 4981
rect 148042 4972 148048 4984
rect 148100 4972 148106 5024
rect 268378 4972 268384 5024
rect 268436 4972 268442 5024
rect 269666 4972 269672 5024
rect 269724 4972 269730 5024
rect 270586 4972 270592 5024
rect 270644 4972 270650 5024
rect 360654 4972 360660 5024
rect 360712 5012 360718 5024
rect 439240 5012 439268 5052
rect 440326 5040 440332 5052
rect 440384 5040 440390 5092
rect 360712 4984 439268 5012
rect 360712 4972 360718 4984
rect 440142 4972 440148 5024
rect 440200 5012 440206 5024
rect 444558 5012 444564 5024
rect 440200 4984 444564 5012
rect 440200 4972 440206 4984
rect 444558 4972 444564 4984
rect 444616 4972 444622 5024
rect 456794 4972 456800 5024
rect 456852 5012 456858 5024
rect 478874 5012 478880 5024
rect 456852 4984 478880 5012
rect 456852 4972 456858 4984
rect 478874 4972 478880 4984
rect 478932 4972 478938 5024
rect 1104 4922 528816 4944
rect 1104 4870 66914 4922
rect 66966 4870 66978 4922
rect 67030 4870 67042 4922
rect 67094 4870 67106 4922
rect 67158 4870 67170 4922
rect 67222 4870 198842 4922
rect 198894 4870 198906 4922
rect 198958 4870 198970 4922
rect 199022 4870 199034 4922
rect 199086 4870 199098 4922
rect 199150 4870 330770 4922
rect 330822 4870 330834 4922
rect 330886 4870 330898 4922
rect 330950 4870 330962 4922
rect 331014 4870 331026 4922
rect 331078 4870 462698 4922
rect 462750 4870 462762 4922
rect 462814 4870 462826 4922
rect 462878 4870 462890 4922
rect 462942 4870 462954 4922
rect 463006 4870 528816 4922
rect 1104 4848 528816 4870
rect 12158 4768 12164 4820
rect 12216 4808 12222 4820
rect 63494 4808 63500 4820
rect 12216 4780 63500 4808
rect 12216 4768 12222 4780
rect 63494 4768 63500 4780
rect 63552 4768 63558 4820
rect 73982 4768 73988 4820
rect 74040 4808 74046 4820
rect 122834 4808 122840 4820
rect 74040 4780 122840 4808
rect 74040 4768 74046 4780
rect 122834 4768 122840 4780
rect 122892 4768 122898 4820
rect 123386 4768 123392 4820
rect 123444 4808 123450 4820
rect 128170 4808 128176 4820
rect 123444 4780 128176 4808
rect 123444 4768 123450 4780
rect 128170 4768 128176 4780
rect 128228 4768 128234 4820
rect 130838 4768 130844 4820
rect 130896 4808 130902 4820
rect 130896 4780 138014 4808
rect 130896 4768 130902 4780
rect 59170 4700 59176 4752
rect 59228 4740 59234 4752
rect 94314 4740 94320 4752
rect 59228 4712 94320 4740
rect 59228 4700 59234 4712
rect 94314 4700 94320 4712
rect 94372 4700 94378 4752
rect 97166 4700 97172 4752
rect 97224 4740 97230 4752
rect 132678 4740 132684 4752
rect 97224 4712 132684 4740
rect 97224 4700 97230 4712
rect 132678 4700 132684 4712
rect 132736 4700 132742 4752
rect 135346 4740 135352 4752
rect 132788 4712 135352 4740
rect 79226 4632 79232 4684
rect 79284 4672 79290 4684
rect 92750 4672 92756 4684
rect 79284 4644 92756 4672
rect 79284 4632 79290 4644
rect 92750 4632 92756 4644
rect 92808 4632 92814 4684
rect 94130 4632 94136 4684
rect 94188 4672 94194 4684
rect 129550 4672 129556 4684
rect 94188 4644 129556 4672
rect 94188 4632 94194 4644
rect 129550 4632 129556 4644
rect 129608 4632 129614 4684
rect 130378 4632 130384 4684
rect 130436 4672 130442 4684
rect 132788 4672 132816 4712
rect 135346 4700 135352 4712
rect 135404 4700 135410 4752
rect 137986 4740 138014 4780
rect 138106 4768 138112 4820
rect 138164 4808 138170 4820
rect 243354 4808 243360 4820
rect 138164 4780 243360 4808
rect 138164 4768 138170 4780
rect 243354 4768 243360 4780
rect 243412 4768 243418 4820
rect 280798 4768 280804 4820
rect 280856 4808 280862 4820
rect 389818 4808 389824 4820
rect 280856 4780 389824 4808
rect 280856 4768 280862 4780
rect 389818 4768 389824 4780
rect 389876 4768 389882 4820
rect 390554 4768 390560 4820
rect 390612 4808 390618 4820
rect 438854 4808 438860 4820
rect 390612 4780 438860 4808
rect 390612 4768 390618 4780
rect 438854 4768 438860 4780
rect 438912 4768 438918 4820
rect 439130 4768 439136 4820
rect 439188 4808 439194 4820
rect 445754 4808 445760 4820
rect 439188 4780 445760 4808
rect 439188 4768 439194 4780
rect 445754 4768 445760 4780
rect 445812 4768 445818 4820
rect 450814 4768 450820 4820
rect 450872 4808 450878 4820
rect 481910 4808 481916 4820
rect 450872 4780 481916 4808
rect 450872 4768 450878 4780
rect 481910 4768 481916 4780
rect 481968 4768 481974 4820
rect 488442 4768 488448 4820
rect 488500 4808 488506 4820
rect 511626 4808 511632 4820
rect 488500 4780 511632 4808
rect 488500 4768 488506 4780
rect 511626 4768 511632 4780
rect 511684 4768 511690 4820
rect 137986 4712 140544 4740
rect 137005 4675 137063 4681
rect 130436 4644 132816 4672
rect 135226 4644 136864 4672
rect 130436 4632 130442 4644
rect 23198 4564 23204 4616
rect 23256 4604 23262 4616
rect 96706 4604 96712 4616
rect 23256 4576 96712 4604
rect 23256 4564 23262 4576
rect 96706 4564 96712 4576
rect 96764 4564 96770 4616
rect 112622 4564 112628 4616
rect 112680 4604 112686 4616
rect 130838 4604 130844 4616
rect 112680 4576 130844 4604
rect 112680 4564 112686 4576
rect 130838 4564 130844 4576
rect 130896 4564 130902 4616
rect 131022 4564 131028 4616
rect 131080 4604 131086 4616
rect 135226 4604 135254 4644
rect 136729 4607 136787 4613
rect 136729 4604 136741 4607
rect 131080 4576 135254 4604
rect 136192 4576 136741 4604
rect 131080 4564 131086 4576
rect 91554 4496 91560 4548
rect 91612 4536 91618 4548
rect 123386 4536 123392 4548
rect 91612 4508 123392 4536
rect 91612 4496 91618 4508
rect 123386 4496 123392 4508
rect 123444 4496 123450 4548
rect 130378 4536 130384 4548
rect 123496 4508 130384 4536
rect 102318 4428 102324 4480
rect 102376 4468 102382 4480
rect 123496 4468 123524 4508
rect 130378 4496 130384 4508
rect 130436 4496 130442 4548
rect 131206 4496 131212 4548
rect 131264 4496 131270 4548
rect 136192 4480 136220 4576
rect 136729 4573 136741 4576
rect 136775 4573 136787 4607
rect 136729 4567 136787 4573
rect 136836 4536 136864 4644
rect 137005 4641 137017 4675
rect 137051 4672 137063 4675
rect 138106 4672 138112 4684
rect 137051 4644 138112 4672
rect 137051 4641 137063 4644
rect 137005 4635 137063 4641
rect 138106 4632 138112 4644
rect 138164 4632 138170 4684
rect 138201 4675 138259 4681
rect 138201 4641 138213 4675
rect 138247 4672 138259 4675
rect 140516 4672 140544 4712
rect 141602 4700 141608 4752
rect 141660 4740 141666 4752
rect 247678 4740 247684 4752
rect 141660 4712 247684 4740
rect 141660 4700 141666 4712
rect 247678 4700 247684 4712
rect 247736 4700 247742 4752
rect 293678 4700 293684 4752
rect 293736 4740 293742 4752
rect 392486 4740 392492 4752
rect 293736 4712 392492 4740
rect 293736 4700 293742 4712
rect 392486 4700 392492 4712
rect 392544 4700 392550 4752
rect 145834 4672 145840 4684
rect 138247 4644 140452 4672
rect 140516 4644 145840 4672
rect 138247 4641 138259 4644
rect 138201 4635 138259 4641
rect 137922 4564 137928 4616
rect 137980 4564 137986 4616
rect 140225 4607 140283 4613
rect 140225 4573 140237 4607
rect 140271 4573 140283 4607
rect 140225 4567 140283 4573
rect 139673 4539 139731 4545
rect 139673 4536 139685 4539
rect 136836 4508 139685 4536
rect 139673 4505 139685 4508
rect 139719 4536 139731 4539
rect 140240 4536 140268 4567
rect 139719 4508 140268 4536
rect 139719 4505 139731 4508
rect 139673 4499 139731 4505
rect 102376 4440 123524 4468
rect 102376 4428 102382 4440
rect 127618 4428 127624 4480
rect 127676 4428 127682 4480
rect 127710 4428 127716 4480
rect 127768 4468 127774 4480
rect 134153 4471 134211 4477
rect 134153 4468 134165 4471
rect 127768 4440 134165 4468
rect 127768 4428 127774 4440
rect 134153 4437 134165 4440
rect 134199 4468 134211 4471
rect 134334 4468 134340 4480
rect 134199 4440 134340 4468
rect 134199 4437 134211 4440
rect 134153 4431 134211 4437
rect 134334 4428 134340 4440
rect 134392 4428 134398 4480
rect 136174 4428 136180 4480
rect 136232 4428 136238 4480
rect 140424 4468 140452 4644
rect 145834 4632 145840 4644
rect 145892 4632 145898 4684
rect 246666 4672 246672 4684
rect 147646 4644 246672 4672
rect 141050 4564 141056 4616
rect 141108 4604 141114 4616
rect 141329 4607 141387 4613
rect 141329 4604 141341 4607
rect 141108 4576 141341 4604
rect 141108 4564 141114 4576
rect 141329 4573 141341 4576
rect 141375 4573 141387 4607
rect 147646 4604 147674 4644
rect 246666 4632 246672 4644
rect 246724 4632 246730 4684
rect 271690 4632 271696 4684
rect 271748 4672 271754 4684
rect 293862 4672 293868 4684
rect 271748 4644 293868 4672
rect 271748 4632 271754 4644
rect 293862 4632 293868 4644
rect 293920 4632 293926 4684
rect 309134 4632 309140 4684
rect 309192 4672 309198 4684
rect 395522 4672 395528 4684
rect 309192 4644 395528 4672
rect 309192 4632 309198 4644
rect 395522 4632 395528 4644
rect 395580 4632 395586 4684
rect 141329 4567 141387 4573
rect 141528 4576 147674 4604
rect 140501 4539 140559 4545
rect 140501 4505 140513 4539
rect 140547 4536 140559 4539
rect 141528 4536 141556 4576
rect 149146 4564 149152 4616
rect 149204 4564 149210 4616
rect 149425 4607 149483 4613
rect 149425 4573 149437 4607
rect 149471 4604 149483 4607
rect 255866 4604 255872 4616
rect 149471 4576 255872 4604
rect 149471 4573 149483 4576
rect 149425 4567 149483 4573
rect 255866 4564 255872 4576
rect 255924 4564 255930 4616
rect 322014 4564 322020 4616
rect 322072 4604 322078 4616
rect 398466 4604 398472 4616
rect 322072 4576 398472 4604
rect 322072 4564 322078 4576
rect 398466 4564 398472 4576
rect 398524 4564 398530 4616
rect 140547 4508 141556 4536
rect 140547 4505 140559 4508
rect 140501 4499 140559 4505
rect 141602 4496 141608 4548
rect 141660 4496 141666 4548
rect 244458 4536 244464 4548
rect 142908 4508 244464 4536
rect 142908 4468 142936 4508
rect 244458 4496 244464 4508
rect 244516 4496 244522 4548
rect 244826 4496 244832 4548
rect 244884 4536 244890 4548
rect 312906 4536 312912 4548
rect 244884 4508 312912 4536
rect 244884 4496 244890 4508
rect 312906 4496 312912 4508
rect 312964 4496 312970 4548
rect 334894 4496 334900 4548
rect 334952 4536 334958 4548
rect 361482 4536 361488 4548
rect 334952 4508 361488 4536
rect 334952 4496 334958 4508
rect 361482 4496 361488 4508
rect 361540 4496 361546 4548
rect 140424 4440 142936 4468
rect 145466 4428 145472 4480
rect 145524 4428 145530 4480
rect 249886 4428 249892 4480
rect 249944 4468 249950 4480
rect 357066 4468 357072 4480
rect 249944 4440 357072 4468
rect 249944 4428 249950 4440
rect 357066 4428 357072 4440
rect 357124 4428 357130 4480
rect 1104 4378 528816 4400
rect 1104 4326 67574 4378
rect 67626 4326 67638 4378
rect 67690 4326 67702 4378
rect 67754 4326 67766 4378
rect 67818 4326 67830 4378
rect 67882 4326 199502 4378
rect 199554 4326 199566 4378
rect 199618 4326 199630 4378
rect 199682 4326 199694 4378
rect 199746 4326 199758 4378
rect 199810 4326 331430 4378
rect 331482 4326 331494 4378
rect 331546 4326 331558 4378
rect 331610 4326 331622 4378
rect 331674 4326 331686 4378
rect 331738 4326 463358 4378
rect 463410 4326 463422 4378
rect 463474 4326 463486 4378
rect 463538 4326 463550 4378
rect 463602 4326 463614 4378
rect 463666 4326 528816 4378
rect 1104 4304 528816 4326
rect 109954 4224 109960 4276
rect 110012 4264 110018 4276
rect 138198 4264 138204 4276
rect 110012 4236 138204 4264
rect 110012 4224 110018 4236
rect 138198 4224 138204 4236
rect 138256 4224 138262 4276
rect 142430 4224 142436 4276
rect 142488 4264 142494 4276
rect 249334 4264 249340 4276
rect 142488 4236 249340 4264
rect 142488 4224 142494 4236
rect 249334 4224 249340 4236
rect 249392 4224 249398 4276
rect 128078 4156 128084 4208
rect 128136 4196 128142 4208
rect 234706 4196 234712 4208
rect 128136 4168 234712 4196
rect 128136 4156 128142 4168
rect 234706 4156 234712 4168
rect 234764 4156 234770 4208
rect 84286 4088 84292 4140
rect 84344 4128 84350 4140
rect 126606 4128 126612 4140
rect 84344 4100 126612 4128
rect 84344 4088 84350 4100
rect 126606 4088 126612 4100
rect 126664 4088 126670 4140
rect 126882 4088 126888 4140
rect 126940 4128 126946 4140
rect 137741 4131 137799 4137
rect 137741 4128 137753 4131
rect 126940 4100 137753 4128
rect 126940 4088 126946 4100
rect 137741 4097 137753 4100
rect 137787 4128 137799 4131
rect 137922 4128 137928 4140
rect 137787 4100 137928 4128
rect 137787 4097 137799 4100
rect 137741 4091 137799 4097
rect 137922 4088 137928 4100
rect 137980 4088 137986 4140
rect 141694 4128 141700 4140
rect 139320 4100 141700 4128
rect 48222 4020 48228 4072
rect 48280 4060 48286 4072
rect 75914 4060 75920 4072
rect 48280 4032 75920 4060
rect 48280 4020 48286 4032
rect 75914 4020 75920 4032
rect 75972 4020 75978 4072
rect 79042 4020 79048 4072
rect 79100 4060 79106 4072
rect 125134 4060 125140 4072
rect 79100 4032 125140 4060
rect 79100 4020 79106 4032
rect 125134 4020 125140 4032
rect 125192 4020 125198 4072
rect 133046 4020 133052 4072
rect 133104 4060 133110 4072
rect 139320 4060 139348 4100
rect 141694 4088 141700 4100
rect 141752 4088 141758 4140
rect 143721 4131 143779 4137
rect 143721 4128 143733 4131
rect 143184 4100 143733 4128
rect 133104 4032 139348 4060
rect 133104 4020 133110 4032
rect 143184 4004 143212 4100
rect 143721 4097 143733 4100
rect 143767 4097 143779 4131
rect 145653 4131 145711 4137
rect 145653 4128 145665 4131
rect 143721 4091 143779 4097
rect 144656 4100 145665 4128
rect 143994 4020 144000 4072
rect 144052 4020 144058 4072
rect 4430 3952 4436 4004
rect 4488 3992 4494 4004
rect 71038 3992 71044 4004
rect 4488 3964 71044 3992
rect 4488 3952 4494 3964
rect 71038 3952 71044 3964
rect 71096 3952 71102 4004
rect 76466 3952 76472 4004
rect 76524 3992 76530 4004
rect 123202 3992 123208 4004
rect 76524 3964 123208 3992
rect 76524 3952 76530 3964
rect 123202 3952 123208 3964
rect 123260 3952 123266 4004
rect 130838 3952 130844 4004
rect 130896 3992 130902 4004
rect 130896 3964 138014 3992
rect 130896 3952 130902 3964
rect 71406 3884 71412 3936
rect 71464 3924 71470 3936
rect 121638 3924 121644 3936
rect 71464 3896 121644 3924
rect 71464 3884 71470 3896
rect 121638 3884 121644 3896
rect 121696 3884 121702 3936
rect 122926 3884 122932 3936
rect 122984 3924 122990 3936
rect 133138 3924 133144 3936
rect 122984 3896 133144 3924
rect 122984 3884 122990 3896
rect 133138 3884 133144 3896
rect 133196 3884 133202 3936
rect 137986 3924 138014 3964
rect 143166 3952 143172 4004
rect 143224 3952 143230 4004
rect 140958 3924 140964 3936
rect 137986 3896 140964 3924
rect 140958 3884 140964 3896
rect 141016 3884 141022 3936
rect 141050 3884 141056 3936
rect 141108 3924 141114 3936
rect 141145 3927 141203 3933
rect 141145 3924 141157 3927
rect 141108 3896 141157 3924
rect 141108 3884 141114 3896
rect 141145 3893 141157 3896
rect 141191 3893 141203 3927
rect 141145 3887 141203 3893
rect 141694 3884 141700 3936
rect 141752 3924 141758 3936
rect 144656 3924 144684 4100
rect 145653 4097 145665 4100
rect 145699 4097 145711 4131
rect 147217 4131 147275 4137
rect 147217 4128 147229 4131
rect 145653 4091 145711 4097
rect 145852 4100 147229 4128
rect 144730 3952 144736 4004
rect 144788 3992 144794 4004
rect 145852 3992 145880 4100
rect 147217 4097 147229 4100
rect 147263 4097 147275 4131
rect 147217 4091 147275 4097
rect 148134 4088 148140 4140
rect 148192 4128 148198 4140
rect 148413 4131 148471 4137
rect 148413 4128 148425 4131
rect 148192 4100 148425 4128
rect 148192 4088 148198 4100
rect 148413 4097 148425 4100
rect 148459 4097 148471 4131
rect 148413 4091 148471 4097
rect 148612 4100 150756 4128
rect 145929 4063 145987 4069
rect 145929 4029 145941 4063
rect 145975 4029 145987 4063
rect 145929 4023 145987 4029
rect 147493 4063 147551 4069
rect 147493 4029 147505 4063
rect 147539 4060 147551 4063
rect 148612 4060 148640 4100
rect 147539 4032 148640 4060
rect 147539 4029 147551 4032
rect 147493 4023 147551 4029
rect 144788 3964 145880 3992
rect 145944 3992 145972 4023
rect 148686 4020 148692 4072
rect 148744 4020 148750 4072
rect 150728 4060 150756 4100
rect 150802 4088 150808 4140
rect 150860 4088 150866 4140
rect 151004 4100 151814 4128
rect 150894 4060 150900 4072
rect 150728 4032 150900 4060
rect 150894 4020 150900 4032
rect 150952 4020 150958 4072
rect 151004 3992 151032 4100
rect 151081 4063 151139 4069
rect 151081 4029 151093 4063
rect 151127 4029 151139 4063
rect 151786 4060 151814 4100
rect 205358 4088 205364 4140
rect 205416 4128 205422 4140
rect 210418 4128 210424 4140
rect 205416 4100 210424 4128
rect 205416 4088 205422 4100
rect 210418 4088 210424 4100
rect 210476 4088 210482 4140
rect 301406 4088 301412 4140
rect 301464 4128 301470 4140
rect 375374 4128 375380 4140
rect 301464 4100 375380 4128
rect 301464 4088 301470 4100
rect 375374 4088 375380 4100
rect 375432 4088 375438 4140
rect 440234 4088 440240 4140
rect 440292 4128 440298 4140
rect 445294 4128 445300 4140
rect 440292 4100 445300 4128
rect 440292 4088 440298 4100
rect 445294 4088 445300 4100
rect 445352 4088 445358 4140
rect 251266 4060 251272 4072
rect 151786 4032 251272 4060
rect 151081 4023 151139 4029
rect 145944 3964 151032 3992
rect 144788 3952 144794 3964
rect 145009 3927 145067 3933
rect 145009 3924 145021 3927
rect 141752 3896 145021 3924
rect 141752 3884 141758 3896
rect 145009 3893 145021 3896
rect 145055 3893 145067 3927
rect 145852 3924 145880 3964
rect 146665 3927 146723 3933
rect 146665 3924 146677 3927
rect 145852 3896 146677 3924
rect 145009 3887 145067 3893
rect 146665 3893 146677 3896
rect 146711 3893 146723 3927
rect 151096 3924 151124 4023
rect 251266 4020 251272 4032
rect 251324 4020 251330 4072
rect 298830 4020 298836 4072
rect 298888 4060 298894 4072
rect 374270 4060 374276 4072
rect 298888 4032 374276 4060
rect 298888 4020 298894 4032
rect 374270 4020 374276 4032
rect 374328 4020 374334 4072
rect 378686 4020 378692 4072
rect 378744 4060 378750 4072
rect 403066 4060 403072 4072
rect 378744 4032 403072 4060
rect 378744 4020 378750 4032
rect 403066 4020 403072 4032
rect 403124 4020 403130 4072
rect 151170 3952 151176 4004
rect 151228 3992 151234 4004
rect 253106 3992 253112 4004
rect 151228 3964 253112 3992
rect 151228 3952 151234 3964
rect 253106 3952 253112 3964
rect 253164 3952 253170 4004
rect 319254 3952 319260 4004
rect 319312 3992 319318 4004
rect 397454 3992 397460 4004
rect 319312 3964 397460 3992
rect 319312 3952 319318 3964
rect 397454 3952 397460 3964
rect 397512 3952 397518 4004
rect 256418 3924 256424 3936
rect 151096 3896 256424 3924
rect 146665 3887 146723 3893
rect 256418 3884 256424 3896
rect 256476 3884 256482 3936
rect 355502 3884 355508 3936
rect 355560 3924 355566 3936
rect 440418 3924 440424 3936
rect 355560 3896 440424 3924
rect 355560 3884 355566 3896
rect 440418 3884 440424 3896
rect 440476 3884 440482 3936
rect 1104 3834 528816 3856
rect 1104 3782 66914 3834
rect 66966 3782 66978 3834
rect 67030 3782 67042 3834
rect 67094 3782 67106 3834
rect 67158 3782 67170 3834
rect 67222 3782 198842 3834
rect 198894 3782 198906 3834
rect 198958 3782 198970 3834
rect 199022 3782 199034 3834
rect 199086 3782 199098 3834
rect 199150 3782 330770 3834
rect 330822 3782 330834 3834
rect 330886 3782 330898 3834
rect 330950 3782 330962 3834
rect 331014 3782 331026 3834
rect 331078 3782 462698 3834
rect 462750 3782 462762 3834
rect 462814 3782 462826 3834
rect 462878 3782 462890 3834
rect 462942 3782 462954 3834
rect 463006 3782 528816 3834
rect 1104 3760 528816 3782
rect 1854 3680 1860 3732
rect 1912 3680 1918 3732
rect 4430 3680 4436 3732
rect 4488 3680 4494 3732
rect 6822 3680 6828 3732
rect 6880 3680 6886 3732
rect 9582 3680 9588 3732
rect 9640 3680 9646 3732
rect 12158 3680 12164 3732
rect 12216 3680 12222 3732
rect 14734 3680 14740 3732
rect 14792 3680 14798 3732
rect 17310 3680 17316 3732
rect 17368 3680 17374 3732
rect 19886 3680 19892 3732
rect 19944 3680 19950 3732
rect 22462 3680 22468 3732
rect 22520 3680 22526 3732
rect 30193 3723 30251 3729
rect 30193 3689 30205 3723
rect 30239 3720 30251 3723
rect 33134 3720 33140 3732
rect 30239 3692 33140 3720
rect 30239 3689 30251 3692
rect 30193 3683 30251 3689
rect 33134 3680 33140 3692
rect 33192 3680 33198 3732
rect 36078 3680 36084 3732
rect 36136 3680 36142 3732
rect 43806 3680 43812 3732
rect 43864 3680 43870 3732
rect 45646 3680 45652 3732
rect 45704 3680 45710 3732
rect 48222 3680 48228 3732
rect 48280 3680 48286 3732
rect 59262 3680 59268 3732
rect 59320 3680 59326 3732
rect 62114 3720 62120 3732
rect 60016 3692 62120 3720
rect 31846 3612 31852 3664
rect 31904 3652 31910 3664
rect 35345 3655 35403 3661
rect 35345 3652 35357 3655
rect 31904 3624 35357 3652
rect 31904 3612 31910 3624
rect 35345 3621 35357 3624
rect 35391 3621 35403 3655
rect 35345 3615 35403 3621
rect 40497 3655 40555 3661
rect 40497 3621 40509 3655
rect 40543 3652 40555 3655
rect 60016 3652 60044 3692
rect 62114 3680 62120 3692
rect 62172 3680 62178 3732
rect 63494 3680 63500 3732
rect 63552 3720 63558 3732
rect 66257 3723 66315 3729
rect 66257 3720 66269 3723
rect 63552 3692 66269 3720
rect 63552 3680 63558 3692
rect 66257 3689 66269 3692
rect 66303 3689 66315 3723
rect 66257 3683 66315 3689
rect 66993 3723 67051 3729
rect 66993 3689 67005 3723
rect 67039 3720 67051 3723
rect 67266 3720 67272 3732
rect 67039 3692 67272 3720
rect 67039 3689 67051 3692
rect 66993 3683 67051 3689
rect 67266 3680 67272 3692
rect 67324 3680 67330 3732
rect 68833 3723 68891 3729
rect 68833 3689 68845 3723
rect 68879 3720 68891 3723
rect 120442 3720 120448 3732
rect 68879 3692 120448 3720
rect 68879 3689 68891 3692
rect 68833 3683 68891 3689
rect 120442 3680 120448 3692
rect 120500 3680 120506 3732
rect 122926 3680 122932 3732
rect 122984 3680 122990 3732
rect 130838 3680 130844 3732
rect 130896 3680 130902 3732
rect 133138 3680 133144 3732
rect 133196 3720 133202 3732
rect 140682 3720 140688 3732
rect 133196 3692 140688 3720
rect 133196 3680 133202 3692
rect 140682 3680 140688 3692
rect 140740 3680 140746 3732
rect 140958 3680 140964 3732
rect 141016 3720 141022 3732
rect 144638 3720 144644 3732
rect 141016 3692 144644 3720
rect 141016 3680 141022 3692
rect 144638 3680 144644 3692
rect 144696 3680 144702 3732
rect 148686 3680 148692 3732
rect 148744 3720 148750 3732
rect 194686 3720 194692 3732
rect 148744 3692 194692 3720
rect 148744 3680 148750 3692
rect 194686 3680 194692 3692
rect 194744 3680 194750 3732
rect 194778 3680 194784 3732
rect 194836 3720 194842 3732
rect 194836 3692 205634 3720
rect 194836 3680 194842 3692
rect 40543 3624 60044 3652
rect 61105 3655 61163 3661
rect 40543 3621 40555 3624
rect 40497 3615 40555 3621
rect 61105 3621 61117 3655
rect 61151 3621 61163 3655
rect 61105 3615 61163 3621
rect 63681 3655 63739 3661
rect 63681 3621 63693 3655
rect 63727 3652 63739 3655
rect 63727 3624 109908 3652
rect 63727 3621 63739 3624
rect 63681 3615 63739 3621
rect 24857 3587 24915 3593
rect 24857 3553 24869 3587
rect 24903 3584 24915 3587
rect 35894 3584 35900 3596
rect 24903 3556 35900 3584
rect 24903 3553 24915 3556
rect 24857 3547 24915 3553
rect 35894 3544 35900 3556
rect 35952 3544 35958 3596
rect 37737 3587 37795 3593
rect 37737 3553 37749 3587
rect 37783 3584 37795 3587
rect 47394 3584 47400 3596
rect 37783 3556 47400 3584
rect 37783 3553 37795 3556
rect 37737 3547 37795 3553
rect 47394 3544 47400 3556
rect 47452 3544 47458 3596
rect 61120 3584 61148 3615
rect 109678 3584 109684 3596
rect 61120 3556 109684 3584
rect 109678 3544 109684 3556
rect 109736 3544 109742 3596
rect 109880 3584 109908 3624
rect 109954 3612 109960 3664
rect 110012 3612 110018 3664
rect 115106 3612 115112 3664
rect 115164 3612 115170 3664
rect 117685 3655 117743 3661
rect 117685 3621 117697 3655
rect 117731 3652 117743 3655
rect 125413 3655 125471 3661
rect 117731 3624 123524 3652
rect 117731 3621 117743 3624
rect 117685 3615 117743 3621
rect 111058 3584 111064 3596
rect 109880 3556 111064 3584
rect 111058 3544 111064 3556
rect 111116 3544 111122 3596
rect 113361 3587 113419 3593
rect 113361 3584 113373 3587
rect 112824 3556 113373 3584
rect 29362 3476 29368 3528
rect 29420 3516 29426 3528
rect 31941 3519 31999 3525
rect 31941 3516 31953 3519
rect 29420 3488 31953 3516
rect 29420 3476 29426 3488
rect 31941 3485 31953 3488
rect 31987 3516 31999 3519
rect 32861 3519 32919 3525
rect 32861 3516 32873 3519
rect 31987 3488 32873 3516
rect 31987 3485 31999 3488
rect 31941 3479 31999 3485
rect 32861 3485 32873 3488
rect 32907 3485 32919 3519
rect 32861 3479 32919 3485
rect 35529 3519 35587 3525
rect 35529 3485 35541 3519
rect 35575 3516 35587 3519
rect 36078 3516 36084 3528
rect 35575 3488 36084 3516
rect 35575 3485 35587 3488
rect 35529 3479 35587 3485
rect 36078 3476 36084 3488
rect 36136 3476 36142 3528
rect 40678 3476 40684 3528
rect 40736 3476 40742 3528
rect 43257 3519 43315 3525
rect 43257 3485 43269 3519
rect 43303 3516 43315 3519
rect 43806 3516 43812 3528
rect 43303 3488 43812 3516
rect 43303 3485 43315 3488
rect 43257 3479 43315 3485
rect 43806 3476 43812 3488
rect 43864 3476 43870 3528
rect 45830 3476 45836 3528
rect 45888 3476 45894 3528
rect 48409 3519 48467 3525
rect 48409 3516 48421 3519
rect 47596 3488 48421 3516
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1949 3451 2007 3457
rect 1949 3448 1961 3451
rect 1360 3420 1961 3448
rect 1360 3408 1366 3420
rect 1949 3417 1961 3420
rect 1995 3417 2007 3451
rect 1949 3411 2007 3417
rect 3970 3408 3976 3460
rect 4028 3448 4034 3460
rect 4525 3451 4583 3457
rect 4525 3448 4537 3451
rect 4028 3420 4537 3448
rect 4028 3408 4034 3420
rect 4525 3417 4537 3420
rect 4571 3417 4583 3451
rect 7101 3451 7159 3457
rect 7101 3448 7113 3451
rect 4525 3411 4583 3417
rect 6886 3420 7113 3448
rect 6178 3340 6184 3392
rect 6236 3380 6242 3392
rect 6886 3380 6914 3420
rect 7101 3417 7113 3420
rect 7147 3417 7159 3451
rect 7101 3411 7159 3417
rect 9122 3408 9128 3460
rect 9180 3448 9186 3460
rect 9677 3451 9735 3457
rect 9677 3448 9689 3451
rect 9180 3420 9689 3448
rect 9180 3408 9186 3420
rect 9677 3417 9689 3420
rect 9723 3417 9735 3451
rect 9677 3411 9735 3417
rect 12253 3451 12311 3457
rect 12253 3417 12265 3451
rect 12299 3417 12311 3451
rect 12253 3411 12311 3417
rect 6236 3352 6914 3380
rect 6236 3340 6242 3352
rect 11330 3340 11336 3392
rect 11388 3380 11394 3392
rect 12268 3380 12296 3411
rect 14274 3408 14280 3460
rect 14332 3448 14338 3460
rect 14829 3451 14887 3457
rect 14829 3448 14841 3451
rect 14332 3420 14841 3448
rect 14332 3408 14338 3420
rect 14829 3417 14841 3420
rect 14875 3417 14887 3451
rect 17405 3451 17463 3457
rect 17405 3448 17417 3451
rect 14829 3411 14887 3417
rect 16592 3420 17417 3448
rect 16592 3392 16620 3420
rect 17405 3417 17417 3420
rect 17451 3417 17463 3451
rect 17405 3411 17463 3417
rect 19242 3408 19248 3460
rect 19300 3448 19306 3460
rect 19981 3451 20039 3457
rect 19981 3448 19993 3451
rect 19300 3420 19993 3448
rect 19300 3408 19306 3420
rect 19981 3417 19993 3420
rect 20027 3417 20039 3451
rect 19981 3411 20039 3417
rect 22557 3451 22615 3457
rect 22557 3417 22569 3451
rect 22603 3417 22615 3451
rect 22557 3411 22615 3417
rect 11388 3352 12296 3380
rect 11388 3340 11394 3352
rect 16574 3340 16580 3392
rect 16632 3340 16638 3392
rect 21634 3340 21640 3392
rect 21692 3380 21698 3392
rect 22572 3380 22600 3411
rect 24578 3408 24584 3460
rect 24636 3448 24642 3460
rect 25133 3451 25191 3457
rect 25133 3448 25145 3451
rect 24636 3420 25145 3448
rect 24636 3408 24642 3420
rect 25133 3417 25145 3420
rect 25179 3417 25191 3451
rect 26881 3451 26939 3457
rect 26881 3448 26893 3451
rect 25133 3411 25191 3417
rect 26206 3420 26893 3448
rect 21692 3352 22600 3380
rect 21692 3340 21698 3352
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 26206 3380 26234 3420
rect 26881 3417 26893 3420
rect 26927 3448 26939 3451
rect 27709 3451 27767 3457
rect 27709 3448 27721 3451
rect 26927 3420 27721 3448
rect 26927 3417 26939 3420
rect 26881 3411 26939 3417
rect 27709 3417 27721 3420
rect 27755 3417 27767 3451
rect 27709 3411 27767 3417
rect 28902 3408 28908 3460
rect 28960 3448 28966 3460
rect 30285 3451 30343 3457
rect 30285 3448 30297 3451
rect 28960 3420 30297 3448
rect 28960 3408 28966 3420
rect 30285 3417 30297 3420
rect 30331 3417 30343 3451
rect 30285 3411 30343 3417
rect 33134 3408 33140 3460
rect 33192 3448 33198 3460
rect 47596 3457 47624 3488
rect 48409 3485 48421 3488
rect 48455 3485 48467 3519
rect 48409 3479 48467 3485
rect 50985 3519 51043 3525
rect 50985 3485 50997 3519
rect 51031 3516 51043 3519
rect 53561 3519 53619 3525
rect 53561 3516 53573 3519
rect 51031 3488 51580 3516
rect 51031 3485 51043 3488
rect 50985 3479 51043 3485
rect 37093 3451 37151 3457
rect 37093 3448 37105 3451
rect 33192 3420 37105 3448
rect 33192 3408 33198 3420
rect 37093 3417 37105 3420
rect 37139 3448 37151 3451
rect 38013 3451 38071 3457
rect 38013 3448 38025 3451
rect 37139 3420 38025 3448
rect 37139 3417 37151 3420
rect 37093 3411 37151 3417
rect 38013 3417 38025 3420
rect 38059 3417 38071 3451
rect 47581 3451 47639 3457
rect 47581 3448 47593 3451
rect 38013 3411 38071 3417
rect 45526 3420 47593 3448
rect 24912 3352 26234 3380
rect 24912 3340 24918 3352
rect 27614 3340 27620 3392
rect 27672 3340 27678 3392
rect 32766 3340 32772 3392
rect 32824 3340 32830 3392
rect 39114 3340 39120 3392
rect 39172 3380 39178 3392
rect 43073 3383 43131 3389
rect 43073 3380 43085 3383
rect 39172 3352 43085 3380
rect 39172 3340 39178 3352
rect 43073 3349 43085 3352
rect 43119 3349 43131 3383
rect 43073 3343 43131 3349
rect 43162 3340 43168 3392
rect 43220 3380 43226 3392
rect 45526 3380 45554 3420
rect 47581 3417 47593 3420
rect 47627 3417 47639 3451
rect 47581 3411 47639 3417
rect 51552 3392 51580 3488
rect 52748 3488 53573 3516
rect 52748 3392 52776 3488
rect 53561 3485 53573 3488
rect 53607 3485 53619 3519
rect 53561 3479 53619 3485
rect 55122 3476 55128 3528
rect 55180 3516 55186 3528
rect 56137 3519 56195 3525
rect 56137 3516 56149 3519
rect 55180 3488 56149 3516
rect 55180 3476 55186 3488
rect 56137 3485 56149 3488
rect 56183 3485 56195 3519
rect 56137 3479 56195 3485
rect 58713 3519 58771 3525
rect 58713 3485 58725 3519
rect 58759 3516 58771 3519
rect 59262 3516 59268 3528
rect 58759 3488 59268 3516
rect 58759 3485 58771 3488
rect 58713 3479 58771 3485
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 60642 3476 60648 3528
rect 60700 3516 60706 3528
rect 61289 3519 61347 3525
rect 61289 3516 61301 3519
rect 60700 3488 61301 3516
rect 60700 3476 60706 3488
rect 61289 3485 61301 3488
rect 61335 3485 61347 3519
rect 63865 3519 63923 3525
rect 63865 3516 63877 3519
rect 61289 3479 61347 3485
rect 63052 3488 63877 3516
rect 62942 3448 62948 3460
rect 55186 3420 62948 3448
rect 43220 3352 45554 3380
rect 43220 3340 43226 3352
rect 49694 3340 49700 3392
rect 49752 3380 49758 3392
rect 50801 3383 50859 3389
rect 50801 3380 50813 3383
rect 49752 3352 50813 3380
rect 49752 3340 49758 3352
rect 50801 3349 50813 3352
rect 50847 3349 50859 3383
rect 50801 3343 50859 3349
rect 51534 3340 51540 3392
rect 51592 3340 51598 3392
rect 52730 3340 52736 3392
rect 52788 3340 52794 3392
rect 53377 3383 53435 3389
rect 53377 3349 53389 3383
rect 53423 3380 53435 3383
rect 55186 3380 55214 3420
rect 62942 3408 62948 3420
rect 63000 3408 63006 3460
rect 53423 3352 55214 3380
rect 53423 3349 53435 3352
rect 53377 3343 53435 3349
rect 55950 3340 55956 3392
rect 56008 3340 56014 3392
rect 56686 3340 56692 3392
rect 56744 3380 56750 3392
rect 58529 3383 58587 3389
rect 58529 3380 58541 3383
rect 56744 3352 58541 3380
rect 56744 3340 56750 3352
rect 58529 3349 58541 3352
rect 58575 3349 58587 3383
rect 58529 3343 58587 3349
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 63052 3389 63080 3488
rect 63865 3485 63877 3488
rect 63911 3485 63923 3519
rect 63865 3479 63923 3485
rect 66441 3519 66499 3525
rect 66441 3485 66453 3519
rect 66487 3516 66499 3519
rect 67266 3516 67272 3528
rect 66487 3488 67272 3516
rect 66487 3485 66499 3488
rect 66441 3479 66499 3485
rect 67266 3476 67272 3488
rect 67324 3476 67330 3528
rect 69014 3476 69020 3528
rect 69072 3476 69078 3528
rect 71222 3476 71228 3528
rect 71280 3516 71286 3528
rect 71593 3519 71651 3525
rect 71593 3516 71605 3519
rect 71280 3488 71605 3516
rect 71280 3476 71286 3488
rect 71593 3485 71605 3488
rect 71639 3485 71651 3519
rect 71593 3479 71651 3485
rect 74169 3519 74227 3525
rect 74169 3485 74181 3519
rect 74215 3516 74227 3519
rect 74718 3516 74724 3528
rect 74215 3488 74724 3516
rect 74215 3485 74227 3488
rect 74169 3479 74227 3485
rect 74718 3476 74724 3488
rect 74776 3476 74782 3528
rect 74920 3488 80054 3516
rect 63126 3408 63132 3460
rect 63184 3448 63190 3460
rect 74920 3448 74948 3488
rect 63184 3420 74948 3448
rect 63184 3408 63190 3420
rect 76466 3408 76472 3460
rect 76524 3408 76530 3460
rect 76650 3408 76656 3460
rect 76708 3408 76714 3460
rect 79042 3408 79048 3460
rect 79100 3408 79106 3460
rect 79229 3451 79287 3457
rect 79229 3417 79241 3451
rect 79275 3417 79287 3451
rect 80026 3448 80054 3488
rect 81894 3476 81900 3528
rect 81952 3476 81958 3528
rect 82004 3488 88748 3516
rect 82004 3448 82032 3488
rect 80026 3420 82032 3448
rect 79229 3411 79287 3417
rect 63037 3383 63095 3389
rect 63037 3380 63049 3383
rect 60792 3352 63049 3380
rect 60792 3340 60798 3352
rect 63037 3349 63049 3352
rect 63083 3349 63095 3383
rect 63037 3343 63095 3349
rect 64874 3340 64880 3392
rect 64932 3380 64938 3392
rect 68189 3383 68247 3389
rect 68189 3380 68201 3383
rect 64932 3352 68201 3380
rect 64932 3340 64938 3352
rect 68189 3349 68201 3352
rect 68235 3380 68247 3383
rect 69014 3380 69020 3392
rect 68235 3352 69020 3380
rect 68235 3349 68247 3352
rect 68189 3343 68247 3349
rect 69014 3340 69020 3352
rect 69072 3340 69078 3392
rect 71406 3340 71412 3392
rect 71464 3340 71470 3392
rect 71498 3340 71504 3392
rect 71556 3380 71562 3392
rect 73985 3383 74043 3389
rect 73985 3380 73997 3383
rect 71556 3352 73997 3380
rect 71556 3340 71562 3352
rect 73985 3349 73997 3352
rect 74031 3349 74043 3383
rect 73985 3343 74043 3349
rect 78490 3340 78496 3392
rect 78548 3380 78554 3392
rect 79244 3380 79272 3411
rect 82446 3408 82452 3460
rect 82504 3408 82510 3460
rect 84381 3451 84439 3457
rect 84381 3448 84393 3451
rect 84166 3420 84393 3448
rect 78548 3352 79272 3380
rect 78548 3340 78554 3352
rect 81526 3340 81532 3392
rect 81584 3380 81590 3392
rect 81713 3383 81771 3389
rect 81713 3380 81725 3383
rect 81584 3352 81725 3380
rect 81584 3340 81590 3352
rect 81713 3349 81725 3352
rect 81759 3349 81771 3383
rect 81713 3343 81771 3349
rect 81894 3340 81900 3392
rect 81952 3380 81958 3392
rect 82464 3380 82492 3408
rect 81952 3352 82492 3380
rect 81952 3340 81958 3352
rect 83642 3340 83648 3392
rect 83700 3380 83706 3392
rect 84166 3380 84194 3420
rect 84381 3417 84393 3420
rect 84427 3417 84439 3451
rect 84381 3411 84439 3417
rect 86954 3408 86960 3460
rect 87012 3408 87018 3460
rect 88720 3448 88748 3488
rect 89622 3476 89628 3528
rect 89680 3476 89686 3528
rect 89714 3476 89720 3528
rect 89772 3516 89778 3528
rect 90174 3516 90180 3528
rect 89772 3488 90180 3516
rect 89772 3476 89778 3488
rect 90174 3476 90180 3488
rect 90232 3476 90238 3528
rect 97353 3519 97411 3525
rect 90928 3488 94820 3516
rect 90928 3448 90956 3488
rect 88720 3420 90956 3448
rect 92106 3408 92112 3460
rect 92164 3408 92170 3460
rect 94685 3451 94743 3457
rect 94685 3448 94697 3451
rect 93964 3420 94697 3448
rect 83700 3352 84194 3380
rect 83700 3340 83706 3352
rect 84286 3340 84292 3392
rect 84344 3340 84350 3392
rect 86862 3340 86868 3392
rect 86920 3340 86926 3392
rect 87414 3340 87420 3392
rect 87472 3380 87478 3392
rect 89441 3383 89499 3389
rect 89441 3380 89453 3383
rect 87472 3352 89453 3380
rect 87472 3340 87478 3352
rect 89441 3349 89453 3352
rect 89487 3349 89499 3383
rect 89441 3343 89499 3349
rect 92014 3340 92020 3392
rect 92072 3340 92078 3392
rect 92566 3340 92572 3392
rect 92624 3380 92630 3392
rect 93964 3389 93992 3420
rect 94685 3417 94697 3420
rect 94731 3417 94743 3451
rect 94792 3448 94820 3488
rect 97353 3485 97365 3519
rect 97399 3516 97411 3519
rect 97902 3516 97908 3528
rect 97399 3488 97908 3516
rect 97399 3485 97411 3488
rect 97353 3479 97411 3485
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98012 3488 103514 3516
rect 98012 3448 98040 3488
rect 99837 3451 99895 3457
rect 99837 3448 99849 3451
rect 94792 3420 98040 3448
rect 99346 3420 99849 3448
rect 94685 3411 94743 3417
rect 93949 3383 94007 3389
rect 93949 3380 93961 3383
rect 92624 3352 93961 3380
rect 92624 3340 92630 3352
rect 93949 3349 93961 3352
rect 93995 3349 94007 3383
rect 93949 3343 94007 3349
rect 94590 3340 94596 3392
rect 94648 3340 94654 3392
rect 94774 3340 94780 3392
rect 94832 3380 94838 3392
rect 97169 3383 97227 3389
rect 97169 3380 97181 3383
rect 94832 3352 97181 3380
rect 94832 3340 94838 3352
rect 97169 3349 97181 3352
rect 97215 3349 97227 3383
rect 97169 3343 97227 3349
rect 97902 3340 97908 3392
rect 97960 3340 97966 3392
rect 99098 3340 99104 3392
rect 99156 3380 99162 3392
rect 99346 3380 99374 3420
rect 99837 3417 99849 3420
rect 99883 3417 99895 3451
rect 99837 3411 99895 3417
rect 102134 3408 102140 3460
rect 102192 3448 102198 3460
rect 102413 3451 102471 3457
rect 102413 3448 102425 3451
rect 102192 3420 102425 3448
rect 102192 3408 102198 3420
rect 102413 3417 102425 3420
rect 102459 3417 102471 3451
rect 103486 3448 103514 3488
rect 105078 3476 105084 3528
rect 105136 3476 105142 3528
rect 112714 3516 112720 3528
rect 105188 3488 112720 3516
rect 105188 3448 105216 3488
rect 112714 3476 112720 3488
rect 112772 3476 112778 3528
rect 112824 3525 112852 3556
rect 113361 3553 113373 3556
rect 113407 3584 113419 3587
rect 123496 3584 123524 3624
rect 125413 3621 125425 3655
rect 125459 3652 125471 3655
rect 133417 3655 133475 3661
rect 125459 3624 133184 3652
rect 125459 3621 125471 3624
rect 125413 3615 125471 3621
rect 133046 3584 133052 3596
rect 113407 3556 123432 3584
rect 123496 3556 133052 3584
rect 113407 3553 113419 3556
rect 113361 3547 113419 3553
rect 112809 3519 112867 3525
rect 112809 3485 112821 3519
rect 112855 3485 112867 3519
rect 117498 3516 117504 3528
rect 112809 3479 112867 3485
rect 112916 3488 117504 3516
rect 103486 3420 105216 3448
rect 102413 3411 102471 3417
rect 105630 3408 105636 3460
rect 105688 3408 105694 3460
rect 107562 3408 107568 3460
rect 107620 3408 107626 3460
rect 110141 3451 110199 3457
rect 110141 3448 110153 3451
rect 109420 3420 110153 3448
rect 99156 3352 99374 3380
rect 99156 3340 99162 3352
rect 99742 3340 99748 3392
rect 99800 3340 99806 3392
rect 102318 3340 102324 3392
rect 102376 3340 102382 3392
rect 102502 3340 102508 3392
rect 102560 3380 102566 3392
rect 104897 3383 104955 3389
rect 104897 3380 104909 3383
rect 102560 3352 104909 3380
rect 102560 3340 102566 3352
rect 104897 3349 104909 3352
rect 104943 3349 104955 3383
rect 104897 3343 104955 3349
rect 107470 3340 107476 3392
rect 107528 3340 107534 3392
rect 109126 3340 109132 3392
rect 109184 3380 109190 3392
rect 109420 3389 109448 3420
rect 110141 3417 110153 3420
rect 110187 3417 110199 3451
rect 110141 3411 110199 3417
rect 111058 3408 111064 3460
rect 111116 3448 111122 3460
rect 112916 3448 112944 3488
rect 117498 3476 117504 3488
rect 117556 3476 117562 3528
rect 120537 3519 120595 3525
rect 120537 3485 120549 3519
rect 120583 3516 120595 3519
rect 123404 3516 123432 3556
rect 133046 3544 133052 3556
rect 133104 3544 133110 3596
rect 133156 3584 133184 3624
rect 133417 3621 133429 3655
rect 133463 3652 133475 3655
rect 134334 3652 134340 3664
rect 133463 3624 134340 3652
rect 133463 3621 133475 3624
rect 133417 3615 133475 3621
rect 134334 3612 134340 3624
rect 134392 3612 134398 3664
rect 135254 3612 135260 3664
rect 135312 3652 135318 3664
rect 135809 3655 135867 3661
rect 135809 3652 135821 3655
rect 135312 3624 135821 3652
rect 135312 3612 135318 3624
rect 135809 3621 135821 3624
rect 135855 3621 135867 3655
rect 135809 3615 135867 3621
rect 188062 3612 188068 3664
rect 188120 3652 188126 3664
rect 195146 3652 195152 3664
rect 188120 3624 195152 3652
rect 188120 3612 188126 3624
rect 195146 3612 195152 3624
rect 195204 3612 195210 3664
rect 196158 3652 196164 3664
rect 195256 3624 196164 3652
rect 145466 3584 145472 3596
rect 133156 3556 145472 3584
rect 145466 3544 145472 3556
rect 145524 3544 145530 3596
rect 148134 3544 148140 3596
rect 148192 3584 148198 3596
rect 148229 3587 148287 3593
rect 148229 3584 148241 3587
rect 148192 3556 148241 3584
rect 148192 3544 148198 3556
rect 148229 3553 148241 3556
rect 148275 3553 148287 3587
rect 148229 3547 148287 3553
rect 158714 3544 158720 3596
rect 158772 3584 158778 3596
rect 179414 3584 179420 3596
rect 158772 3556 179420 3584
rect 158772 3544 158778 3556
rect 179414 3544 179420 3556
rect 179472 3544 179478 3596
rect 180794 3544 180800 3596
rect 180852 3584 180858 3596
rect 195256 3584 195284 3624
rect 196158 3612 196164 3624
rect 196216 3612 196222 3664
rect 205606 3652 205634 3692
rect 210418 3680 210424 3732
rect 210476 3720 210482 3732
rect 265986 3720 265992 3732
rect 210476 3692 265992 3720
rect 210476 3680 210482 3692
rect 265986 3680 265992 3692
rect 266044 3680 266050 3732
rect 270494 3680 270500 3732
rect 270552 3720 270558 3732
rect 357434 3720 357440 3732
rect 270552 3692 357440 3720
rect 270552 3680 270558 3692
rect 357434 3680 357440 3692
rect 357492 3680 357498 3732
rect 372614 3680 372620 3732
rect 372672 3720 372678 3732
rect 399294 3720 399300 3732
rect 372672 3692 399300 3720
rect 372672 3680 372678 3692
rect 399294 3680 399300 3692
rect 399352 3680 399358 3732
rect 301222 3652 301228 3664
rect 205606 3624 301228 3652
rect 301222 3612 301228 3624
rect 301280 3612 301286 3664
rect 306558 3612 306564 3664
rect 306616 3652 306622 3664
rect 395154 3652 395160 3664
rect 306616 3624 395160 3652
rect 306616 3612 306622 3624
rect 395154 3612 395160 3624
rect 395212 3612 395218 3664
rect 420914 3612 420920 3664
rect 420972 3652 420978 3664
rect 444374 3652 444380 3664
rect 420972 3624 444380 3652
rect 420972 3612 420978 3624
rect 444374 3612 444380 3624
rect 444432 3612 444438 3664
rect 180852 3556 195284 3584
rect 180852 3544 180858 3556
rect 195330 3544 195336 3596
rect 195388 3584 195394 3596
rect 296162 3584 296168 3596
rect 195388 3556 296168 3584
rect 195388 3544 195394 3556
rect 296162 3544 296168 3556
rect 296220 3544 296226 3596
rect 303982 3544 303988 3596
rect 304040 3584 304046 3596
rect 392118 3584 392124 3596
rect 304040 3556 392124 3584
rect 304040 3544 304046 3556
rect 392118 3544 392124 3556
rect 392176 3544 392182 3596
rect 435358 3544 435364 3596
rect 435416 3584 435422 3596
rect 480346 3584 480352 3596
rect 435416 3556 480352 3584
rect 435416 3544 435422 3556
rect 480346 3544 480352 3556
rect 480404 3544 480410 3596
rect 128265 3519 128323 3525
rect 120583 3488 121132 3516
rect 123404 3488 128216 3516
rect 120583 3485 120595 3488
rect 120537 3479 120595 3485
rect 115293 3451 115351 3457
rect 115293 3448 115305 3451
rect 111116 3420 112944 3448
rect 114572 3420 115305 3448
rect 111116 3408 111122 3420
rect 114572 3392 114600 3420
rect 115293 3417 115305 3420
rect 115339 3417 115351 3451
rect 115293 3411 115351 3417
rect 117590 3408 117596 3460
rect 117648 3448 117654 3460
rect 117869 3451 117927 3457
rect 117869 3448 117881 3451
rect 117648 3420 117881 3448
rect 117648 3408 117654 3420
rect 117869 3417 117881 3420
rect 117915 3417 117927 3451
rect 117869 3411 117927 3417
rect 121104 3392 121132 3488
rect 122650 3408 122656 3460
rect 122708 3448 122714 3460
rect 123021 3451 123079 3457
rect 123021 3448 123033 3451
rect 122708 3420 123033 3448
rect 122708 3408 122714 3420
rect 123021 3417 123033 3420
rect 123067 3417 123079 3451
rect 125597 3451 125655 3457
rect 125597 3448 125609 3451
rect 123021 3411 123079 3417
rect 124876 3420 125609 3448
rect 109405 3383 109463 3389
rect 109405 3380 109417 3383
rect 109184 3352 109417 3380
rect 109184 3340 109190 3352
rect 109405 3349 109417 3352
rect 109451 3349 109463 3383
rect 109405 3343 109463 3349
rect 111886 3340 111892 3392
rect 111944 3380 111950 3392
rect 112625 3383 112683 3389
rect 112625 3380 112637 3383
rect 111944 3352 112637 3380
rect 111944 3340 111950 3352
rect 112625 3349 112637 3352
rect 112671 3349 112683 3383
rect 112625 3343 112683 3349
rect 114554 3340 114560 3392
rect 114612 3340 114618 3392
rect 119338 3340 119344 3392
rect 119396 3380 119402 3392
rect 120353 3383 120411 3389
rect 120353 3380 120365 3383
rect 119396 3352 120365 3380
rect 119396 3340 119402 3352
rect 120353 3349 120365 3352
rect 120399 3349 120411 3383
rect 120353 3343 120411 3349
rect 121086 3340 121092 3392
rect 121144 3340 121150 3392
rect 124214 3340 124220 3392
rect 124272 3380 124278 3392
rect 124876 3389 124904 3420
rect 125597 3417 125609 3420
rect 125643 3417 125655 3451
rect 125597 3411 125655 3417
rect 124861 3383 124919 3389
rect 124861 3380 124873 3383
rect 124272 3352 124873 3380
rect 124272 3340 124278 3352
rect 124861 3349 124873 3352
rect 124907 3349 124919 3383
rect 124861 3343 124919 3349
rect 125686 3340 125692 3392
rect 125744 3380 125750 3392
rect 128081 3383 128139 3389
rect 128081 3380 128093 3383
rect 125744 3352 128093 3380
rect 125744 3340 125750 3352
rect 128081 3349 128093 3352
rect 128127 3349 128139 3383
rect 128188 3380 128216 3488
rect 128265 3485 128277 3519
rect 128311 3516 128323 3519
rect 128311 3488 128860 3516
rect 128311 3485 128323 3488
rect 128265 3479 128323 3485
rect 128832 3457 128860 3488
rect 130470 3476 130476 3528
rect 130528 3516 130534 3528
rect 130657 3519 130715 3525
rect 130657 3516 130669 3519
rect 130528 3488 130669 3516
rect 130528 3476 130534 3488
rect 130657 3485 130669 3488
rect 130703 3516 130715 3519
rect 131301 3519 131359 3525
rect 131301 3516 131313 3519
rect 130703 3488 131313 3516
rect 130703 3485 130715 3488
rect 130657 3479 130715 3485
rect 131301 3485 131313 3488
rect 131347 3485 131359 3519
rect 131301 3479 131359 3485
rect 132494 3476 132500 3528
rect 132552 3516 132558 3528
rect 133233 3519 133291 3525
rect 133233 3516 133245 3519
rect 132552 3488 133245 3516
rect 132552 3476 132558 3488
rect 133233 3485 133245 3488
rect 133279 3516 133291 3519
rect 133877 3519 133935 3525
rect 133877 3516 133889 3519
rect 133279 3488 133889 3516
rect 133279 3485 133291 3488
rect 133233 3479 133291 3485
rect 133877 3485 133889 3488
rect 133923 3485 133935 3519
rect 133877 3479 133935 3485
rect 135993 3519 136051 3525
rect 135993 3485 136005 3519
rect 136039 3516 136051 3519
rect 136545 3519 136603 3525
rect 136545 3516 136557 3519
rect 136039 3488 136557 3516
rect 136039 3485 136051 3488
rect 135993 3479 136051 3485
rect 136545 3485 136557 3488
rect 136591 3516 136603 3519
rect 243722 3516 243728 3528
rect 136591 3488 243728 3516
rect 136591 3485 136603 3488
rect 136545 3479 136603 3485
rect 243722 3476 243728 3488
rect 243780 3476 243786 3528
rect 273070 3476 273076 3528
rect 273128 3516 273134 3528
rect 365806 3516 365812 3528
rect 273128 3488 365812 3516
rect 273128 3476 273134 3488
rect 365806 3476 365812 3488
rect 365864 3476 365870 3528
rect 395430 3476 395436 3528
rect 395488 3516 395494 3528
rect 442074 3516 442080 3528
rect 395488 3488 442080 3516
rect 395488 3476 395494 3488
rect 442074 3476 442080 3488
rect 442132 3476 442138 3528
rect 128817 3451 128875 3457
rect 128817 3417 128829 3451
rect 128863 3448 128875 3451
rect 128863 3420 135852 3448
rect 128863 3417 128875 3420
rect 128817 3411 128875 3417
rect 128354 3380 128360 3392
rect 128188 3352 128360 3380
rect 128081 3343 128139 3349
rect 128354 3340 128360 3352
rect 128412 3340 128418 3392
rect 135824 3380 135852 3420
rect 136082 3408 136088 3460
rect 136140 3448 136146 3460
rect 220538 3448 220544 3460
rect 136140 3420 220544 3448
rect 136140 3408 136146 3420
rect 220538 3408 220544 3420
rect 220596 3408 220602 3460
rect 257614 3408 257620 3460
rect 257672 3448 257678 3460
rect 363690 3448 363696 3460
rect 257672 3420 363696 3448
rect 257672 3408 257678 3420
rect 363690 3408 363696 3420
rect 363748 3408 363754 3460
rect 397362 3408 397368 3460
rect 397420 3448 397426 3460
rect 443454 3448 443460 3460
rect 397420 3420 443460 3448
rect 397420 3408 397426 3420
rect 443454 3408 443460 3420
rect 443512 3408 443518 3460
rect 455966 3408 455972 3460
rect 456024 3448 456030 3460
rect 482278 3448 482284 3460
rect 456024 3420 482284 3448
rect 456024 3408 456030 3420
rect 482278 3408 482284 3420
rect 482336 3408 482342 3460
rect 235994 3380 236000 3392
rect 135824 3352 236000 3380
rect 235994 3340 236000 3352
rect 236052 3340 236058 3392
rect 296254 3340 296260 3392
rect 296312 3380 296318 3392
rect 364702 3380 364708 3392
rect 296312 3352 364708 3380
rect 296312 3340 296318 3352
rect 364702 3340 364708 3352
rect 364760 3340 364766 3392
rect 1104 3290 528816 3312
rect 1104 3238 67574 3290
rect 67626 3238 67638 3290
rect 67690 3238 67702 3290
rect 67754 3238 67766 3290
rect 67818 3238 67830 3290
rect 67882 3238 199502 3290
rect 199554 3238 199566 3290
rect 199618 3238 199630 3290
rect 199682 3238 199694 3290
rect 199746 3238 199758 3290
rect 199810 3238 331430 3290
rect 331482 3238 331494 3290
rect 331546 3238 331558 3290
rect 331610 3238 331622 3290
rect 331674 3238 331686 3290
rect 331738 3238 463358 3290
rect 463410 3238 463422 3290
rect 463474 3238 463486 3290
rect 463538 3238 463550 3290
rect 463602 3238 463614 3290
rect 463666 3238 528816 3290
rect 1104 3216 528816 3238
rect 61102 3136 61108 3188
rect 61160 3176 61166 3188
rect 82814 3176 82820 3188
rect 61160 3148 82820 3176
rect 61160 3136 61166 3148
rect 82814 3136 82820 3148
rect 82872 3136 82878 3188
rect 94590 3136 94596 3188
rect 94648 3176 94654 3188
rect 131758 3176 131764 3188
rect 94648 3148 131764 3176
rect 94648 3136 94654 3148
rect 131758 3136 131764 3148
rect 131816 3136 131822 3188
rect 132862 3136 132868 3188
rect 132920 3176 132926 3188
rect 189166 3176 189172 3188
rect 132920 3148 189172 3176
rect 132920 3136 132926 3148
rect 189166 3136 189172 3148
rect 189224 3136 189230 3188
rect 194686 3136 194692 3188
rect 194744 3176 194750 3188
rect 254210 3176 254216 3188
rect 194744 3148 254216 3176
rect 194744 3136 194750 3148
rect 254210 3136 254216 3148
rect 254268 3136 254274 3188
rect 351914 3136 351920 3188
rect 351972 3176 351978 3188
rect 396258 3176 396264 3188
rect 351972 3148 396264 3176
rect 351972 3136 351978 3148
rect 396258 3136 396264 3148
rect 396316 3136 396322 3188
rect 485774 3136 485780 3188
rect 485832 3176 485838 3188
rect 485869 3179 485927 3185
rect 485869 3176 485881 3179
rect 485832 3148 485881 3176
rect 485832 3136 485838 3148
rect 485869 3145 485881 3148
rect 485915 3145 485927 3179
rect 485869 3139 485927 3145
rect 488534 3136 488540 3188
rect 488592 3136 488598 3188
rect 491018 3136 491024 3188
rect 491076 3136 491082 3188
rect 493594 3136 493600 3188
rect 493652 3136 493658 3188
rect 496170 3136 496176 3188
rect 496228 3136 496234 3188
rect 498746 3136 498752 3188
rect 498804 3136 498810 3188
rect 501322 3136 501328 3188
rect 501380 3136 501386 3188
rect 503898 3136 503904 3188
rect 503956 3136 503962 3188
rect 506474 3136 506480 3188
rect 506532 3136 506538 3188
rect 509050 3136 509056 3188
rect 509108 3136 509114 3188
rect 511626 3136 511632 3188
rect 511684 3136 511690 3188
rect 71222 3068 71228 3120
rect 71280 3068 71286 3120
rect 74534 3068 74540 3120
rect 74592 3108 74598 3120
rect 78490 3108 78496 3120
rect 74592 3080 78496 3108
rect 74592 3068 74598 3080
rect 78490 3068 78496 3080
rect 78548 3068 78554 3120
rect 78674 3068 78680 3120
rect 78732 3108 78738 3120
rect 83642 3108 83648 3120
rect 78732 3080 83648 3108
rect 78732 3068 78738 3080
rect 83642 3068 83648 3080
rect 83700 3068 83706 3120
rect 86862 3068 86868 3120
rect 86920 3108 86926 3120
rect 91554 3108 91560 3120
rect 86920 3080 91560 3108
rect 86920 3068 86926 3080
rect 91554 3068 91560 3080
rect 91612 3068 91618 3120
rect 96706 3068 96712 3120
rect 96764 3108 96770 3120
rect 99098 3108 99104 3120
rect 96764 3080 99104 3108
rect 96764 3068 96770 3080
rect 99098 3068 99104 3080
rect 99156 3068 99162 3120
rect 99742 3068 99748 3120
rect 99800 3108 99806 3120
rect 133598 3108 133604 3120
rect 99800 3080 133604 3108
rect 99800 3068 99806 3080
rect 133598 3068 133604 3080
rect 133656 3068 133662 3120
rect 136082 3108 136088 3120
rect 133708 3080 136088 3108
rect 27614 3000 27620 3052
rect 27672 3040 27678 3052
rect 27672 3012 89714 3040
rect 27672 3000 27678 3012
rect 51534 2932 51540 2984
rect 51592 2972 51598 2984
rect 85574 2972 85580 2984
rect 51592 2944 85580 2972
rect 51592 2932 51598 2944
rect 85574 2932 85580 2944
rect 85632 2932 85638 2984
rect 89686 2972 89714 3012
rect 100846 3000 100852 3052
rect 100904 3040 100910 3052
rect 107197 3043 107255 3049
rect 107197 3040 107209 3043
rect 100904 3012 107209 3040
rect 100904 3000 100910 3012
rect 107197 3009 107209 3012
rect 107243 3040 107255 3043
rect 107562 3040 107568 3052
rect 107243 3012 107568 3040
rect 107243 3009 107255 3012
rect 107197 3003 107255 3009
rect 107562 3000 107568 3012
rect 107620 3000 107626 3052
rect 109678 3000 109684 3052
rect 109736 3040 109742 3052
rect 116670 3040 116676 3052
rect 109736 3012 116676 3040
rect 109736 3000 109742 3012
rect 116670 3000 116676 3012
rect 116728 3000 116734 3052
rect 117590 3000 117596 3052
rect 117648 3000 117654 3052
rect 128354 3000 128360 3052
rect 128412 3040 128418 3052
rect 133708 3040 133736 3080
rect 136082 3068 136088 3080
rect 136140 3068 136146 3120
rect 181070 3068 181076 3120
rect 181128 3108 181134 3120
rect 205450 3108 205456 3120
rect 181128 3080 205456 3108
rect 181128 3068 181134 3080
rect 205450 3068 205456 3080
rect 205508 3068 205514 3120
rect 210510 3068 210516 3120
rect 210568 3108 210574 3120
rect 252646 3108 252652 3120
rect 210568 3080 252652 3108
rect 210568 3068 210574 3080
rect 252646 3068 252652 3080
rect 252704 3068 252710 3120
rect 128412 3012 133736 3040
rect 128412 3000 128418 3012
rect 134334 3000 134340 3052
rect 134392 3040 134398 3052
rect 149146 3040 149152 3052
rect 134392 3012 149152 3040
rect 134392 3000 134398 3012
rect 149146 3000 149152 3012
rect 149204 3000 149210 3052
rect 184198 3000 184204 3052
rect 184256 3040 184262 3052
rect 192846 3040 192852 3052
rect 184256 3012 192852 3040
rect 184256 3000 184262 3012
rect 192846 3000 192852 3012
rect 192904 3000 192910 3052
rect 195974 3000 195980 3052
rect 196032 3040 196038 3052
rect 212534 3040 212540 3052
rect 196032 3012 212540 3040
rect 196032 3000 196038 3012
rect 212534 3000 212540 3012
rect 212592 3000 212598 3052
rect 101214 2972 101220 2984
rect 89686 2944 101220 2972
rect 101214 2932 101220 2944
rect 101272 2932 101278 2984
rect 107470 2932 107476 2984
rect 107528 2972 107534 2984
rect 137002 2972 137008 2984
rect 107528 2944 137008 2972
rect 107528 2932 107534 2944
rect 137002 2932 137008 2944
rect 137060 2932 137066 2984
rect 143994 2932 144000 2984
rect 144052 2972 144058 2984
rect 249978 2972 249984 2984
rect 144052 2944 249984 2972
rect 144052 2932 144058 2944
rect 249978 2932 249984 2944
rect 250036 2932 250042 2984
rect 36814 2864 36820 2916
rect 36872 2904 36878 2916
rect 40221 2907 40279 2913
rect 40221 2904 40233 2907
rect 36872 2876 40233 2904
rect 36872 2864 36878 2876
rect 40221 2873 40233 2876
rect 40267 2904 40279 2907
rect 40678 2904 40684 2916
rect 40267 2876 40684 2904
rect 40267 2873 40279 2876
rect 40221 2867 40279 2873
rect 40678 2864 40684 2876
rect 40736 2864 40742 2916
rect 41322 2864 41328 2916
rect 41380 2904 41386 2916
rect 45373 2907 45431 2913
rect 45373 2904 45385 2907
rect 41380 2876 45385 2904
rect 41380 2864 41386 2876
rect 45373 2873 45385 2876
rect 45419 2904 45431 2907
rect 45830 2904 45836 2916
rect 45419 2876 45836 2904
rect 45419 2873 45431 2876
rect 45373 2867 45431 2873
rect 45830 2864 45836 2876
rect 45888 2864 45894 2916
rect 67910 2864 67916 2916
rect 67968 2904 67974 2916
rect 71222 2904 71228 2916
rect 67968 2876 71228 2904
rect 67968 2864 67974 2876
rect 71222 2864 71228 2876
rect 71280 2864 71286 2916
rect 71774 2864 71780 2916
rect 71832 2904 71838 2916
rect 76285 2907 76343 2913
rect 76285 2904 76297 2907
rect 71832 2876 76297 2904
rect 71832 2864 71838 2876
rect 76285 2873 76297 2876
rect 76331 2904 76343 2907
rect 76650 2904 76656 2916
rect 76331 2876 76656 2904
rect 76331 2873 76343 2876
rect 76285 2867 76343 2873
rect 76650 2864 76656 2876
rect 76708 2864 76714 2916
rect 80054 2864 80060 2916
rect 80112 2904 80118 2916
rect 86589 2907 86647 2913
rect 86589 2904 86601 2907
rect 80112 2876 86601 2904
rect 80112 2864 80118 2876
rect 86589 2873 86601 2876
rect 86635 2904 86647 2907
rect 86954 2904 86960 2916
rect 86635 2876 86960 2904
rect 86635 2873 86647 2876
rect 86589 2867 86647 2873
rect 86954 2864 86960 2876
rect 87012 2864 87018 2916
rect 92014 2864 92020 2916
rect 92072 2904 92078 2916
rect 130102 2904 130108 2916
rect 92072 2876 130108 2904
rect 92072 2864 92078 2876
rect 130102 2864 130108 2876
rect 130160 2864 130166 2916
rect 166902 2864 166908 2916
rect 166960 2904 166966 2916
rect 194597 2907 194655 2913
rect 194597 2904 194609 2907
rect 166960 2876 194609 2904
rect 166960 2864 166966 2876
rect 194597 2873 194609 2876
rect 194643 2904 194655 2907
rect 195146 2904 195152 2916
rect 194643 2876 195152 2904
rect 194643 2873 194655 2876
rect 194597 2867 194655 2873
rect 195146 2864 195152 2876
rect 195204 2864 195210 2916
rect 202414 2904 202420 2916
rect 195256 2876 202420 2904
rect 1302 2796 1308 2848
rect 1360 2836 1366 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1360 2808 1593 2836
rect 1360 2796 1366 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 3970 2796 3976 2848
rect 4028 2796 4034 2848
rect 6546 2796 6552 2848
rect 6604 2796 6610 2848
rect 8478 2796 8484 2848
rect 8536 2836 8542 2848
rect 9122 2836 9128 2848
rect 8536 2808 9128 2836
rect 8536 2796 8542 2808
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 14274 2796 14280 2848
rect 14332 2796 14338 2848
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 19429 2839 19487 2845
rect 19429 2836 19441 2839
rect 19300 2808 19441 2836
rect 19300 2796 19306 2808
rect 19429 2805 19441 2808
rect 19475 2805 19487 2839
rect 19429 2799 19487 2805
rect 23842 2796 23848 2848
rect 23900 2836 23906 2848
rect 24578 2836 24584 2848
rect 23900 2808 24584 2836
rect 23900 2796 23906 2808
rect 24578 2796 24584 2808
rect 24636 2796 24642 2848
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 29733 2839 29791 2845
rect 29733 2836 29745 2839
rect 28960 2808 29745 2836
rect 28960 2796 28966 2808
rect 29733 2805 29745 2808
rect 29779 2805 29791 2839
rect 29733 2799 29791 2805
rect 34882 2796 34888 2848
rect 34940 2796 34946 2848
rect 37458 2796 37464 2848
rect 37516 2796 37522 2848
rect 42794 2796 42800 2848
rect 42852 2796 42858 2848
rect 50522 2796 50528 2848
rect 50580 2796 50586 2848
rect 53098 2796 53104 2848
rect 53156 2796 53162 2848
rect 53834 2796 53840 2848
rect 53892 2836 53898 2848
rect 55122 2836 55128 2848
rect 53892 2808 55128 2836
rect 53892 2796 53898 2808
rect 55122 2796 55128 2808
rect 55180 2836 55186 2848
rect 55677 2839 55735 2845
rect 55677 2836 55689 2839
rect 55180 2808 55689 2836
rect 55180 2796 55186 2808
rect 55677 2805 55689 2808
rect 55723 2805 55735 2839
rect 55677 2799 55735 2805
rect 58250 2796 58256 2848
rect 58308 2796 58314 2848
rect 59354 2796 59360 2848
rect 59412 2836 59418 2848
rect 60642 2836 60648 2848
rect 59412 2808 60648 2836
rect 59412 2796 59418 2808
rect 60642 2796 60648 2808
rect 60700 2836 60706 2848
rect 60829 2839 60887 2845
rect 60829 2836 60841 2839
rect 60700 2808 60841 2836
rect 60700 2796 60706 2808
rect 60829 2805 60841 2808
rect 60875 2805 60887 2839
rect 60829 2799 60887 2805
rect 65242 2796 65248 2848
rect 65300 2836 65306 2848
rect 65981 2839 66039 2845
rect 65981 2836 65993 2839
rect 65300 2808 65993 2836
rect 65300 2796 65306 2808
rect 65981 2805 65993 2808
rect 66027 2805 66039 2839
rect 65981 2799 66039 2805
rect 68554 2796 68560 2848
rect 68612 2796 68618 2848
rect 70394 2796 70400 2848
rect 70452 2836 70458 2848
rect 71498 2836 71504 2848
rect 70452 2808 71504 2836
rect 70452 2796 70458 2808
rect 71498 2796 71504 2808
rect 71556 2796 71562 2848
rect 73154 2796 73160 2848
rect 73212 2836 73218 2848
rect 73709 2839 73767 2845
rect 73709 2836 73721 2839
rect 73212 2808 73721 2836
rect 73212 2796 73218 2808
rect 73709 2805 73721 2808
rect 73755 2805 73767 2839
rect 73709 2799 73767 2805
rect 81434 2796 81440 2848
rect 81492 2796 81498 2848
rect 84010 2796 84016 2848
rect 84068 2796 84074 2848
rect 89257 2839 89315 2845
rect 89257 2805 89269 2839
rect 89303 2836 89315 2839
rect 89530 2836 89536 2848
rect 89303 2808 89536 2836
rect 89303 2805 89315 2808
rect 89257 2799 89315 2805
rect 89530 2796 89536 2808
rect 89588 2796 89594 2848
rect 89714 2796 89720 2848
rect 89772 2836 89778 2848
rect 91741 2839 91799 2845
rect 91741 2836 91753 2839
rect 89772 2808 91753 2836
rect 89772 2796 89778 2808
rect 91741 2805 91753 2808
rect 91787 2836 91799 2839
rect 92106 2836 92112 2848
rect 91787 2808 92112 2836
rect 91787 2805 91799 2808
rect 91741 2799 91799 2805
rect 92106 2796 92112 2808
rect 92164 2796 92170 2848
rect 96614 2796 96620 2848
rect 96672 2836 96678 2848
rect 96893 2839 96951 2845
rect 96893 2836 96905 2839
rect 96672 2808 96905 2836
rect 96672 2796 96678 2808
rect 96893 2805 96905 2808
rect 96939 2805 96951 2839
rect 96893 2799 96951 2805
rect 99466 2796 99472 2848
rect 99524 2796 99530 2848
rect 102134 2796 102140 2848
rect 102192 2796 102198 2848
rect 104618 2796 104624 2848
rect 104676 2796 104682 2848
rect 107378 2796 107384 2848
rect 107436 2836 107442 2848
rect 111702 2836 111708 2848
rect 107436 2808 111708 2836
rect 107436 2796 107442 2808
rect 111702 2796 111708 2808
rect 111760 2796 111766 2848
rect 112346 2796 112352 2848
rect 112404 2796 112410 2848
rect 112990 2796 112996 2848
rect 113048 2836 113054 2848
rect 114646 2836 114652 2848
rect 113048 2808 114652 2836
rect 113048 2796 113054 2808
rect 114646 2796 114652 2808
rect 114704 2796 114710 2848
rect 115017 2839 115075 2845
rect 115017 2805 115029 2839
rect 115063 2836 115075 2839
rect 115290 2836 115296 2848
rect 115063 2808 115296 2836
rect 115063 2805 115075 2808
rect 115017 2799 115075 2805
rect 115290 2796 115296 2808
rect 115348 2796 115354 2848
rect 120074 2796 120080 2848
rect 120132 2796 120138 2848
rect 121454 2796 121460 2848
rect 121512 2836 121518 2848
rect 122650 2836 122656 2848
rect 121512 2808 122656 2836
rect 121512 2796 121518 2808
rect 122650 2796 122656 2808
rect 122708 2796 122714 2848
rect 127897 2839 127955 2845
rect 127897 2805 127909 2839
rect 127943 2836 127955 2839
rect 128170 2836 128176 2848
rect 127943 2808 128176 2836
rect 127943 2805 127955 2808
rect 127897 2799 127955 2805
rect 128170 2796 128176 2808
rect 128228 2796 128234 2848
rect 138014 2796 138020 2848
rect 138072 2796 138078 2848
rect 143074 2796 143080 2848
rect 143132 2796 143138 2848
rect 148226 2796 148232 2848
rect 148284 2796 148290 2848
rect 153378 2796 153384 2848
rect 153436 2796 153442 2848
rect 158530 2796 158536 2848
rect 158588 2796 158594 2848
rect 163682 2796 163688 2848
rect 163740 2796 163746 2848
rect 168374 2796 168380 2848
rect 168432 2836 168438 2848
rect 168837 2839 168895 2845
rect 168837 2836 168849 2839
rect 168432 2808 168849 2836
rect 168432 2796 168438 2808
rect 168837 2805 168849 2808
rect 168883 2805 168895 2839
rect 168837 2799 168895 2805
rect 173986 2796 173992 2848
rect 174044 2796 174050 2848
rect 178034 2796 178040 2848
rect 178092 2836 178098 2848
rect 179138 2836 179144 2848
rect 178092 2808 179144 2836
rect 178092 2796 178098 2808
rect 179138 2796 179144 2808
rect 179196 2796 179202 2848
rect 183554 2796 183560 2848
rect 183612 2836 183618 2848
rect 184293 2839 184351 2845
rect 184293 2836 184305 2839
rect 183612 2808 184305 2836
rect 183612 2796 183618 2808
rect 184293 2805 184305 2808
rect 184339 2805 184351 2839
rect 184293 2799 184351 2805
rect 189074 2796 189080 2848
rect 189132 2836 189138 2848
rect 189445 2839 189503 2845
rect 189445 2836 189457 2839
rect 189132 2808 189457 2836
rect 189132 2796 189138 2808
rect 189445 2805 189457 2808
rect 189491 2805 189503 2839
rect 189445 2799 189503 2805
rect 190454 2796 190460 2848
rect 190512 2836 190518 2848
rect 195256 2836 195284 2876
rect 202414 2864 202420 2876
rect 202472 2864 202478 2916
rect 190512 2808 195284 2836
rect 190512 2796 190518 2808
rect 200022 2796 200028 2848
rect 200080 2796 200086 2848
rect 205082 2796 205088 2848
rect 205140 2796 205146 2848
rect 210234 2796 210240 2848
rect 210292 2796 210298 2848
rect 215386 2796 215392 2848
rect 215444 2796 215450 2848
rect 220538 2796 220544 2848
rect 220596 2796 220602 2848
rect 225785 2839 225843 2845
rect 225785 2805 225797 2839
rect 225831 2836 225843 2839
rect 226058 2836 226064 2848
rect 225831 2808 226064 2836
rect 225831 2805 225843 2808
rect 225785 2799 225843 2805
rect 226058 2796 226064 2808
rect 226116 2796 226122 2848
rect 514202 2796 514208 2848
rect 514260 2796 514266 2848
rect 1104 2746 528816 2768
rect 1104 2694 66914 2746
rect 66966 2694 66978 2746
rect 67030 2694 67042 2746
rect 67094 2694 67106 2746
rect 67158 2694 67170 2746
rect 67222 2694 198842 2746
rect 198894 2694 198906 2746
rect 198958 2694 198970 2746
rect 199022 2694 199034 2746
rect 199086 2694 199098 2746
rect 199150 2694 330770 2746
rect 330822 2694 330834 2746
rect 330886 2694 330898 2746
rect 330950 2694 330962 2746
rect 331014 2694 331026 2746
rect 331078 2694 462698 2746
rect 462750 2694 462762 2746
rect 462814 2694 462826 2746
rect 462878 2694 462890 2746
rect 462942 2694 462954 2746
rect 463006 2694 528816 2746
rect 1104 2672 528816 2694
rect 5166 2592 5172 2644
rect 5224 2592 5230 2644
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 59170 2632 59176 2644
rect 9631 2604 59176 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 59170 2592 59176 2604
rect 59228 2592 59234 2644
rect 61102 2592 61108 2644
rect 61160 2592 61166 2644
rect 68830 2592 68836 2644
rect 68888 2592 68894 2644
rect 73982 2592 73988 2644
rect 74040 2592 74046 2644
rect 76558 2592 76564 2644
rect 76616 2592 76622 2644
rect 81710 2592 81716 2644
rect 81768 2592 81774 2644
rect 87598 2592 87604 2644
rect 87656 2592 87662 2644
rect 92017 2635 92075 2641
rect 92017 2601 92029 2635
rect 92063 2632 92075 2635
rect 92382 2632 92388 2644
rect 92063 2604 92388 2632
rect 92063 2601 92075 2604
rect 92017 2595 92075 2601
rect 92382 2592 92388 2604
rect 92440 2592 92446 2644
rect 97166 2592 97172 2644
rect 97224 2592 97230 2644
rect 99098 2592 99104 2644
rect 99156 2632 99162 2644
rect 102321 2635 102379 2641
rect 102321 2632 102333 2635
rect 99156 2604 102333 2632
rect 99156 2592 99162 2604
rect 102321 2601 102333 2604
rect 102367 2601 102379 2635
rect 102321 2595 102379 2601
rect 103054 2592 103060 2644
rect 103112 2592 103118 2644
rect 103422 2592 103428 2644
rect 103480 2632 103486 2644
rect 107838 2632 107844 2644
rect 103480 2604 107844 2632
rect 103480 2592 103486 2604
rect 107838 2592 107844 2604
rect 107896 2592 107902 2644
rect 107930 2592 107936 2644
rect 107988 2632 107994 2644
rect 109034 2632 109040 2644
rect 107988 2604 109040 2632
rect 107988 2592 107994 2604
rect 109034 2592 109040 2604
rect 109092 2592 109098 2644
rect 110046 2592 110052 2644
rect 110104 2592 110110 2644
rect 110782 2592 110788 2644
rect 110840 2592 110846 2644
rect 112622 2592 112628 2644
rect 112680 2592 112686 2644
rect 126882 2632 126888 2644
rect 115906 2604 126888 2632
rect 12894 2524 12900 2576
rect 12952 2524 12958 2576
rect 18046 2524 18052 2576
rect 18104 2524 18110 2576
rect 19797 2567 19855 2573
rect 19797 2533 19809 2567
rect 19843 2564 19855 2567
rect 42886 2564 42892 2576
rect 19843 2536 42892 2564
rect 19843 2533 19855 2536
rect 19797 2527 19855 2533
rect 42886 2524 42892 2536
rect 42944 2524 42950 2576
rect 43073 2567 43131 2573
rect 43073 2533 43085 2567
rect 43119 2564 43131 2567
rect 45649 2567 45707 2573
rect 43119 2536 45554 2564
rect 43119 2533 43131 2536
rect 43073 2527 43131 2533
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 1719 2468 31754 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2428 4675 2431
rect 5166 2428 5172 2440
rect 4663 2400 5172 2428
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 6788 2400 8493 2428
rect 6788 2388 6794 2400
rect 8481 2397 8493 2400
rect 8527 2428 8539 2431
rect 9677 2431 9735 2437
rect 9677 2428 9689 2431
rect 8527 2400 9689 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 9677 2397 9689 2400
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12894 2428 12900 2440
rect 12391 2400 12900 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2428 17555 2431
rect 18046 2428 18052 2440
rect 17543 2400 18052 2428
rect 17543 2397 17555 2400
rect 17497 2391 17555 2397
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 27801 2431 27859 2437
rect 27801 2397 27813 2431
rect 27847 2428 27859 2431
rect 27847 2400 28396 2428
rect 27847 2397 27859 2400
rect 27801 2391 27859 2397
rect 842 2320 848 2372
rect 900 2360 906 2372
rect 1949 2363 2007 2369
rect 1949 2360 1961 2363
rect 900 2332 1961 2360
rect 900 2320 906 2332
rect 1949 2329 1961 2332
rect 1995 2360 2007 2363
rect 2501 2363 2559 2369
rect 2501 2360 2513 2363
rect 1995 2332 2513 2360
rect 1995 2329 2007 2332
rect 1949 2323 2007 2329
rect 2501 2329 2513 2332
rect 2547 2329 2559 2363
rect 2501 2323 2559 2329
rect 5994 2320 6000 2372
rect 6052 2360 6058 2372
rect 6546 2360 6552 2372
rect 6052 2332 6552 2360
rect 6052 2320 6058 2332
rect 6546 2320 6552 2332
rect 6604 2360 6610 2372
rect 7101 2363 7159 2369
rect 7101 2360 7113 2363
rect 6604 2332 7113 2360
rect 6604 2320 6610 2332
rect 7101 2329 7113 2332
rect 7147 2329 7159 2363
rect 7101 2323 7159 2329
rect 10778 2320 10784 2372
rect 10836 2360 10842 2372
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 10836 2332 13645 2360
rect 10836 2320 10842 2332
rect 13633 2329 13645 2332
rect 13679 2360 13691 2363
rect 14829 2363 14887 2369
rect 14829 2360 14841 2363
rect 13679 2332 14841 2360
rect 13679 2329 13691 2332
rect 13633 2323 13691 2329
rect 14829 2329 14841 2332
rect 14875 2329 14887 2363
rect 14829 2323 14887 2329
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 18785 2363 18843 2369
rect 18785 2360 18797 2363
rect 15988 2332 18797 2360
rect 15988 2320 15994 2332
rect 18785 2329 18797 2332
rect 18831 2360 18843 2363
rect 19981 2363 20039 2369
rect 19981 2360 19993 2363
rect 18831 2332 19993 2360
rect 18831 2329 18843 2332
rect 18785 2323 18843 2329
rect 19981 2329 19993 2332
rect 20027 2329 20039 2363
rect 22664 2360 22692 2391
rect 28368 2372 28396 2400
rect 23198 2360 23204 2372
rect 22664 2332 23204 2360
rect 19981 2323 20039 2329
rect 23198 2320 23204 2332
rect 23256 2320 23262 2372
rect 25133 2363 25191 2369
rect 25133 2360 25145 2363
rect 23952 2332 25145 2360
rect 23952 2304 23980 2332
rect 25133 2329 25145 2332
rect 25179 2329 25191 2363
rect 25133 2323 25191 2329
rect 28350 2320 28356 2372
rect 28408 2320 28414 2372
rect 30285 2363 30343 2369
rect 30285 2360 30297 2363
rect 29104 2332 30297 2360
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4433 2295 4491 2301
rect 4433 2292 4445 2295
rect 4212 2264 4445 2292
rect 4212 2252 4218 2264
rect 4433 2261 4445 2264
rect 4479 2261 4491 2295
rect 4433 2255 4491 2261
rect 7006 2252 7012 2304
rect 7064 2252 7070 2304
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 12161 2295 12219 2301
rect 12161 2292 12173 2295
rect 9640 2264 12173 2292
rect 9640 2252 9646 2264
rect 12161 2261 12173 2264
rect 12207 2261 12219 2295
rect 12161 2255 12219 2261
rect 14734 2252 14740 2304
rect 14792 2252 14798 2304
rect 17310 2252 17316 2304
rect 17368 2252 17374 2304
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 22465 2295 22523 2301
rect 22465 2292 22477 2295
rect 20772 2264 22477 2292
rect 20772 2252 20778 2264
rect 22465 2261 22477 2264
rect 22511 2261 22523 2295
rect 22465 2255 22523 2261
rect 23934 2252 23940 2304
rect 23992 2252 23998 2304
rect 25038 2252 25044 2304
rect 25096 2252 25102 2304
rect 27614 2252 27620 2304
rect 27672 2252 27678 2304
rect 28258 2252 28264 2304
rect 28316 2292 28322 2304
rect 29104 2301 29132 2332
rect 30285 2329 30297 2332
rect 30331 2329 30343 2363
rect 31726 2360 31754 2468
rect 33502 2456 33508 2508
rect 33560 2456 33566 2508
rect 41230 2496 41236 2508
rect 40696 2468 41236 2496
rect 32953 2431 33011 2437
rect 32953 2397 32965 2431
rect 32999 2428 33011 2431
rect 33520 2428 33548 2456
rect 40402 2428 40408 2440
rect 32999 2400 33548 2428
rect 33612 2400 40408 2428
rect 32999 2397 33011 2400
rect 32953 2391 33011 2397
rect 33612 2360 33640 2400
rect 40402 2388 40408 2400
rect 40460 2388 40466 2440
rect 40696 2437 40724 2468
rect 41230 2456 41236 2468
rect 41288 2456 41294 2508
rect 45526 2496 45554 2536
rect 45649 2533 45661 2567
rect 45695 2564 45707 2567
rect 45695 2536 104112 2564
rect 45695 2533 45707 2536
rect 45649 2527 45707 2533
rect 103974 2496 103980 2508
rect 45526 2468 103980 2496
rect 103974 2456 103980 2468
rect 104032 2456 104038 2508
rect 40681 2431 40739 2437
rect 40681 2397 40693 2431
rect 40727 2397 40739 2431
rect 40681 2391 40739 2397
rect 42794 2388 42800 2440
rect 42852 2428 42858 2440
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 42852 2400 43269 2428
rect 42852 2388 42858 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 43257 2391 43315 2397
rect 44560 2400 45845 2428
rect 31726 2332 33640 2360
rect 30285 2323 30343 2329
rect 34882 2320 34888 2372
rect 34940 2360 34946 2372
rect 35437 2363 35495 2369
rect 35437 2360 35449 2363
rect 34940 2332 35449 2360
rect 34940 2320 34946 2332
rect 35437 2329 35449 2332
rect 35483 2329 35495 2363
rect 35437 2323 35495 2329
rect 37458 2320 37464 2372
rect 37516 2360 37522 2372
rect 38013 2363 38071 2369
rect 38013 2360 38025 2363
rect 37516 2332 38025 2360
rect 37516 2320 37522 2332
rect 38013 2329 38025 2332
rect 38059 2329 38071 2363
rect 38013 2323 38071 2329
rect 29089 2295 29147 2301
rect 29089 2292 29101 2295
rect 28316 2264 29101 2292
rect 28316 2252 28322 2264
rect 29089 2261 29101 2264
rect 29135 2261 29147 2295
rect 29089 2255 29147 2261
rect 30190 2252 30196 2304
rect 30248 2252 30254 2304
rect 32766 2252 32772 2304
rect 32824 2252 32830 2304
rect 35342 2252 35348 2304
rect 35400 2252 35406 2304
rect 37918 2252 37924 2304
rect 37976 2252 37982 2304
rect 38654 2252 38660 2304
rect 38712 2292 38718 2304
rect 40497 2295 40555 2301
rect 40497 2292 40509 2295
rect 38712 2264 40509 2292
rect 38712 2252 38718 2264
rect 40497 2261 40509 2264
rect 40543 2261 40555 2295
rect 40497 2255 40555 2261
rect 44082 2252 44088 2304
rect 44140 2292 44146 2304
rect 44560 2301 44588 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 48409 2431 48467 2437
rect 48409 2397 48421 2431
rect 48455 2428 48467 2431
rect 48958 2428 48964 2440
rect 48455 2400 48964 2428
rect 48455 2397 48467 2400
rect 48409 2391 48467 2397
rect 48958 2388 48964 2400
rect 49016 2388 49022 2440
rect 50522 2388 50528 2440
rect 50580 2428 50586 2440
rect 50985 2431 51043 2437
rect 50985 2428 50997 2431
rect 50580 2400 50997 2428
rect 50580 2388 50586 2400
rect 50985 2397 50997 2400
rect 51031 2397 51043 2431
rect 50985 2391 51043 2397
rect 53098 2388 53104 2440
rect 53156 2428 53162 2440
rect 53558 2428 53564 2440
rect 53156 2400 53564 2428
rect 53156 2388 53162 2400
rect 53558 2388 53564 2400
rect 53616 2388 53622 2440
rect 56137 2431 56195 2437
rect 56137 2397 56149 2431
rect 56183 2428 56195 2431
rect 56594 2428 56600 2440
rect 56183 2400 56600 2428
rect 56183 2397 56195 2400
rect 56137 2391 56195 2397
rect 56594 2388 56600 2400
rect 56652 2388 56658 2440
rect 57974 2388 57980 2440
rect 58032 2428 58038 2440
rect 58250 2428 58256 2440
rect 58032 2400 58256 2428
rect 58032 2388 58038 2400
rect 58250 2388 58256 2400
rect 58308 2428 58314 2440
rect 58713 2431 58771 2437
rect 58713 2428 58725 2431
rect 58308 2400 58725 2428
rect 58308 2388 58314 2400
rect 58713 2397 58725 2400
rect 58759 2397 58771 2431
rect 61289 2431 61347 2437
rect 61289 2428 61301 2431
rect 58713 2391 58771 2397
rect 60706 2400 61301 2428
rect 52638 2320 52644 2372
rect 52696 2360 52702 2372
rect 52696 2332 55996 2360
rect 52696 2320 52702 2332
rect 44545 2295 44603 2301
rect 44545 2292 44557 2295
rect 44140 2264 44557 2292
rect 44140 2252 44146 2264
rect 44545 2261 44557 2264
rect 44591 2261 44603 2295
rect 44545 2255 44603 2261
rect 46014 2252 46020 2304
rect 46072 2292 46078 2304
rect 48225 2295 48283 2301
rect 48225 2292 48237 2295
rect 46072 2264 48237 2292
rect 46072 2252 46078 2264
rect 48225 2261 48237 2264
rect 48271 2261 48283 2295
rect 48225 2255 48283 2261
rect 50798 2252 50804 2304
rect 50856 2252 50862 2304
rect 53374 2252 53380 2304
rect 53432 2252 53438 2304
rect 55968 2301 55996 2332
rect 57882 2320 57888 2372
rect 57940 2360 57946 2372
rect 60001 2363 60059 2369
rect 60001 2360 60013 2363
rect 57940 2332 60013 2360
rect 57940 2320 57946 2332
rect 60001 2329 60013 2332
rect 60047 2360 60059 2363
rect 60706 2360 60734 2400
rect 61289 2397 61301 2400
rect 61335 2397 61347 2431
rect 61289 2391 61347 2397
rect 63865 2431 63923 2437
rect 63865 2397 63877 2431
rect 63911 2428 63923 2431
rect 63911 2400 64460 2428
rect 63911 2397 63923 2400
rect 63865 2391 63923 2397
rect 60047 2332 60734 2360
rect 60047 2329 60059 2332
rect 60001 2323 60059 2329
rect 64432 2304 64460 2400
rect 65242 2388 65248 2440
rect 65300 2428 65306 2440
rect 66441 2431 66499 2437
rect 66441 2428 66453 2431
rect 65300 2400 66453 2428
rect 65300 2388 65306 2400
rect 66441 2397 66453 2400
rect 66487 2397 66499 2431
rect 66441 2391 66499 2397
rect 68554 2388 68560 2440
rect 68612 2428 68618 2440
rect 69017 2431 69075 2437
rect 69017 2428 69029 2431
rect 68612 2400 69029 2428
rect 68612 2388 68618 2400
rect 69017 2397 69029 2400
rect 69063 2397 69075 2431
rect 69017 2391 69075 2397
rect 71593 2431 71651 2437
rect 71593 2397 71605 2431
rect 71639 2428 71651 2431
rect 71639 2400 72188 2428
rect 71639 2397 71651 2400
rect 71593 2391 71651 2397
rect 72160 2304 72188 2400
rect 73154 2388 73160 2440
rect 73212 2428 73218 2440
rect 74169 2431 74227 2437
rect 74169 2428 74181 2431
rect 73212 2400 74181 2428
rect 73212 2388 73218 2400
rect 74169 2397 74181 2400
rect 74215 2397 74227 2431
rect 74169 2391 74227 2397
rect 75546 2388 75552 2440
rect 75604 2428 75610 2440
rect 79226 2428 79232 2440
rect 75604 2400 79232 2428
rect 75604 2388 75610 2400
rect 79226 2388 79232 2400
rect 79284 2388 79290 2440
rect 79321 2431 79379 2437
rect 79321 2397 79333 2431
rect 79367 2428 79379 2431
rect 87049 2431 87107 2437
rect 79367 2400 79916 2428
rect 79367 2397 79379 2400
rect 79321 2391 79379 2397
rect 76653 2363 76711 2369
rect 76653 2360 76665 2363
rect 75472 2332 76665 2360
rect 75472 2304 75500 2332
rect 76653 2329 76665 2332
rect 76699 2329 76711 2363
rect 76653 2323 76711 2329
rect 79888 2304 79916 2400
rect 87049 2397 87061 2431
rect 87095 2428 87107 2431
rect 87598 2428 87604 2440
rect 87095 2400 87604 2428
rect 87095 2397 87107 2400
rect 87049 2391 87107 2397
rect 87598 2388 87604 2400
rect 87656 2388 87662 2440
rect 89349 2431 89407 2437
rect 89349 2397 89361 2431
rect 89395 2428 89407 2431
rect 94130 2428 94136 2440
rect 89395 2400 94136 2428
rect 89395 2397 89407 2400
rect 89349 2391 89407 2397
rect 94130 2388 94136 2400
rect 94188 2388 94194 2440
rect 94777 2431 94835 2437
rect 94777 2397 94789 2431
rect 94823 2428 94835 2431
rect 95326 2428 95332 2440
rect 94823 2400 95332 2428
rect 94823 2397 94835 2400
rect 94777 2391 94835 2397
rect 95326 2388 95332 2400
rect 95384 2388 95390 2440
rect 99190 2388 99196 2440
rect 99248 2428 99254 2440
rect 102505 2431 102563 2437
rect 99248 2400 102088 2428
rect 99248 2388 99254 2400
rect 81434 2320 81440 2372
rect 81492 2360 81498 2372
rect 81805 2363 81863 2369
rect 81805 2360 81817 2363
rect 81492 2332 81817 2360
rect 81492 2320 81498 2332
rect 81805 2329 81817 2332
rect 81851 2329 81863 2363
rect 81805 2323 81863 2329
rect 84102 2320 84108 2372
rect 84160 2360 84166 2372
rect 84381 2363 84439 2369
rect 84381 2360 84393 2363
rect 84160 2332 84393 2360
rect 84160 2320 84166 2332
rect 84381 2329 84393 2332
rect 84427 2329 84439 2363
rect 84381 2323 84439 2329
rect 86770 2320 86776 2372
rect 86828 2360 86834 2372
rect 89530 2360 89536 2372
rect 86828 2332 89536 2360
rect 86828 2320 86834 2332
rect 89530 2320 89536 2332
rect 89588 2320 89594 2372
rect 91005 2363 91063 2369
rect 91005 2360 91017 2363
rect 89686 2332 91017 2360
rect 55953 2295 56011 2301
rect 55953 2261 55965 2295
rect 55999 2261 56011 2295
rect 55953 2255 56011 2261
rect 58526 2252 58532 2304
rect 58584 2252 58590 2304
rect 63678 2252 63684 2304
rect 63736 2252 63742 2304
rect 64414 2252 64420 2304
rect 64472 2252 64478 2304
rect 66254 2252 66260 2304
rect 66312 2252 66318 2304
rect 71406 2252 71412 2304
rect 71464 2252 71470 2304
rect 72142 2252 72148 2304
rect 72200 2252 72206 2304
rect 75454 2252 75460 2304
rect 75512 2252 75518 2304
rect 77294 2252 77300 2304
rect 77352 2292 77358 2304
rect 79137 2295 79195 2301
rect 79137 2292 79149 2295
rect 77352 2264 79149 2292
rect 77352 2252 77358 2264
rect 79137 2261 79149 2264
rect 79183 2261 79195 2295
rect 79137 2255 79195 2261
rect 79870 2252 79876 2304
rect 79928 2252 79934 2304
rect 84286 2252 84292 2304
rect 84344 2252 84350 2304
rect 84470 2252 84476 2304
rect 84528 2292 84534 2304
rect 86865 2295 86923 2301
rect 86865 2292 86877 2295
rect 84528 2264 86877 2292
rect 84528 2252 84534 2264
rect 86865 2261 86877 2264
rect 86911 2261 86923 2295
rect 86865 2255 86923 2261
rect 86954 2252 86960 2304
rect 87012 2292 87018 2304
rect 89686 2292 89714 2332
rect 91005 2329 91017 2332
rect 91051 2360 91063 2363
rect 92109 2363 92167 2369
rect 92109 2360 92121 2363
rect 91051 2332 92121 2360
rect 91051 2329 91063 2332
rect 91005 2323 91063 2329
rect 92109 2329 92121 2332
rect 92155 2329 92167 2363
rect 92109 2323 92167 2329
rect 92216 2332 94728 2360
rect 87012 2264 89714 2292
rect 87012 2252 87018 2264
rect 91278 2252 91284 2304
rect 91336 2292 91342 2304
rect 92216 2292 92244 2332
rect 91336 2264 92244 2292
rect 91336 2252 91342 2264
rect 92290 2252 92296 2304
rect 92348 2292 92354 2304
rect 94593 2295 94651 2301
rect 94593 2292 94605 2295
rect 92348 2264 94605 2292
rect 92348 2252 92354 2264
rect 94593 2261 94605 2264
rect 94639 2261 94651 2295
rect 94700 2292 94728 2332
rect 96614 2320 96620 2372
rect 96672 2360 96678 2372
rect 97261 2363 97319 2369
rect 97261 2360 97273 2363
rect 96672 2332 97273 2360
rect 96672 2320 96678 2332
rect 97261 2329 97273 2332
rect 97307 2329 97319 2363
rect 99466 2360 99472 2372
rect 97261 2323 97319 2329
rect 99346 2332 99472 2360
rect 99346 2292 99374 2332
rect 99466 2320 99472 2332
rect 99524 2360 99530 2372
rect 99837 2363 99895 2369
rect 99837 2360 99849 2363
rect 99524 2332 99849 2360
rect 99524 2320 99530 2332
rect 99837 2329 99849 2332
rect 99883 2329 99895 2363
rect 102060 2360 102088 2400
rect 102505 2397 102517 2431
rect 102551 2428 102563 2431
rect 103054 2428 103060 2440
rect 102551 2400 103060 2428
rect 102551 2397 102563 2400
rect 102505 2391 102563 2397
rect 103054 2388 103060 2400
rect 103112 2388 103118 2440
rect 104084 2428 104112 2536
rect 104158 2524 104164 2576
rect 104216 2564 104222 2576
rect 104216 2536 104296 2564
rect 104216 2524 104222 2536
rect 104268 2496 104296 2536
rect 107378 2524 107384 2576
rect 107436 2524 107442 2576
rect 111702 2524 111708 2576
rect 111760 2564 111766 2576
rect 115906 2564 115934 2604
rect 126882 2592 126888 2604
rect 126940 2592 126946 2644
rect 141142 2592 141148 2644
rect 141200 2632 141206 2644
rect 141697 2635 141755 2641
rect 141697 2632 141709 2635
rect 141200 2604 141709 2632
rect 141200 2592 141206 2604
rect 141697 2601 141709 2604
rect 141743 2632 141755 2635
rect 187326 2632 187332 2644
rect 141743 2604 187332 2632
rect 141743 2601 141755 2604
rect 141697 2595 141755 2601
rect 187326 2592 187332 2604
rect 187384 2592 187390 2644
rect 187418 2592 187424 2644
rect 187476 2632 187482 2644
rect 192481 2635 192539 2641
rect 192481 2632 192493 2635
rect 187476 2604 192493 2632
rect 187476 2592 187482 2604
rect 192481 2601 192493 2604
rect 192527 2601 192539 2635
rect 192481 2595 192539 2601
rect 193214 2592 193220 2644
rect 193272 2632 193278 2644
rect 194502 2632 194508 2644
rect 193272 2604 194508 2632
rect 193272 2592 193278 2604
rect 194502 2592 194508 2604
rect 194560 2592 194566 2644
rect 205358 2592 205364 2644
rect 205416 2592 205422 2644
rect 208578 2592 208584 2644
rect 208636 2592 208642 2644
rect 210510 2592 210516 2644
rect 210568 2592 210574 2644
rect 224126 2592 224132 2644
rect 224184 2592 224190 2644
rect 229186 2592 229192 2644
rect 229244 2592 229250 2644
rect 231854 2592 231860 2644
rect 231912 2632 231918 2644
rect 232866 2632 232872 2644
rect 231912 2604 232872 2632
rect 231912 2592 231918 2604
rect 232866 2592 232872 2604
rect 232924 2592 232930 2644
rect 234430 2592 234436 2644
rect 234488 2592 234494 2644
rect 237006 2592 237012 2644
rect 237064 2592 237070 2644
rect 242158 2592 242164 2644
rect 242216 2592 242222 2644
rect 244737 2635 244795 2641
rect 244737 2601 244749 2635
rect 244783 2632 244795 2635
rect 244826 2632 244832 2644
rect 244783 2604 244832 2632
rect 244783 2601 244795 2604
rect 244737 2595 244795 2601
rect 244826 2592 244832 2604
rect 244884 2592 244890 2644
rect 247218 2592 247224 2644
rect 247276 2592 247282 2644
rect 249886 2592 249892 2644
rect 249944 2592 249950 2644
rect 257614 2592 257620 2644
rect 257672 2592 257678 2644
rect 260190 2592 260196 2644
rect 260248 2592 260254 2644
rect 265342 2592 265348 2644
rect 265400 2592 265406 2644
rect 270494 2592 270500 2644
rect 270552 2592 270558 2644
rect 273070 2592 273076 2644
rect 273128 2592 273134 2644
rect 275646 2592 275652 2644
rect 275704 2592 275710 2644
rect 280798 2592 280804 2644
rect 280856 2592 280862 2644
rect 283374 2592 283380 2644
rect 283432 2592 283438 2644
rect 285950 2592 285956 2644
rect 286008 2592 286014 2644
rect 288526 2592 288532 2644
rect 288584 2592 288590 2644
rect 291102 2592 291108 2644
rect 291160 2592 291166 2644
rect 293678 2592 293684 2644
rect 293736 2592 293742 2644
rect 296254 2592 296260 2644
rect 296312 2592 296318 2644
rect 298830 2592 298836 2644
rect 298888 2592 298894 2644
rect 301406 2592 301412 2644
rect 301464 2592 301470 2644
rect 303249 2635 303307 2641
rect 303249 2632 303261 2635
rect 302206 2604 303261 2632
rect 111760 2536 115934 2564
rect 117777 2567 117835 2573
rect 111760 2524 111766 2536
rect 117777 2533 117789 2567
rect 117823 2533 117835 2567
rect 117777 2527 117835 2533
rect 118513 2567 118571 2573
rect 118513 2533 118525 2567
rect 118559 2564 118571 2567
rect 172514 2564 172520 2576
rect 118559 2536 172520 2564
rect 118559 2533 118571 2536
rect 118513 2527 118571 2533
rect 107654 2496 107660 2508
rect 104268 2468 107660 2496
rect 107654 2456 107660 2468
rect 107712 2456 107718 2508
rect 107838 2456 107844 2508
rect 107896 2496 107902 2508
rect 110046 2496 110052 2508
rect 107896 2468 110052 2496
rect 107896 2456 107902 2468
rect 110046 2456 110052 2468
rect 110104 2456 110110 2508
rect 110322 2456 110328 2508
rect 110380 2496 110386 2508
rect 117792 2496 117820 2527
rect 110380 2468 117820 2496
rect 110380 2456 110386 2468
rect 109770 2428 109776 2440
rect 104084 2400 109776 2428
rect 109770 2388 109776 2400
rect 109828 2388 109834 2440
rect 110233 2431 110291 2437
rect 110233 2397 110245 2431
rect 110279 2428 110291 2431
rect 110782 2428 110788 2440
rect 110279 2400 110788 2428
rect 110279 2397 110291 2400
rect 110233 2391 110291 2397
rect 110782 2388 110788 2400
rect 110840 2388 110846 2440
rect 117961 2431 118019 2437
rect 117961 2397 117973 2431
rect 118007 2428 118019 2431
rect 118528 2428 118556 2527
rect 172514 2524 172520 2536
rect 172572 2524 172578 2576
rect 172606 2524 172612 2576
rect 172664 2564 172670 2576
rect 176746 2564 176752 2576
rect 172664 2536 176752 2564
rect 172664 2524 172670 2536
rect 176746 2524 176752 2536
rect 176804 2524 176810 2576
rect 177206 2524 177212 2576
rect 177264 2564 177270 2576
rect 177761 2567 177819 2573
rect 177761 2564 177773 2567
rect 177264 2536 177773 2564
rect 177264 2524 177270 2536
rect 177761 2533 177773 2536
rect 177807 2564 177819 2567
rect 180794 2564 180800 2576
rect 177807 2536 180800 2564
rect 177807 2533 177819 2536
rect 177761 2527 177819 2533
rect 180794 2524 180800 2536
rect 180852 2524 180858 2576
rect 182910 2524 182916 2576
rect 182968 2524 182974 2576
rect 184661 2567 184719 2573
rect 184661 2533 184673 2567
rect 184707 2564 184719 2567
rect 260834 2564 260840 2576
rect 184707 2536 260840 2564
rect 184707 2533 184719 2536
rect 184661 2527 184719 2533
rect 260834 2524 260840 2536
rect 260892 2524 260898 2576
rect 282454 2524 282460 2576
rect 282512 2564 282518 2576
rect 290369 2567 290427 2573
rect 290369 2564 290381 2567
rect 282512 2536 290381 2564
rect 282512 2524 282518 2536
rect 290369 2533 290381 2536
rect 290415 2533 290427 2567
rect 290369 2527 290427 2533
rect 291194 2524 291200 2576
rect 291252 2564 291258 2576
rect 295521 2567 295579 2573
rect 295521 2564 295533 2567
rect 291252 2536 295533 2564
rect 291252 2524 291258 2536
rect 295521 2533 295533 2536
rect 295567 2533 295579 2567
rect 300673 2567 300731 2573
rect 300673 2564 300685 2567
rect 295521 2527 295579 2533
rect 295628 2536 300685 2564
rect 126422 2456 126428 2508
rect 126480 2496 126486 2508
rect 130470 2496 130476 2508
rect 126480 2468 130476 2496
rect 126480 2456 126486 2468
rect 130470 2456 130476 2468
rect 130528 2456 130534 2508
rect 136453 2499 136511 2505
rect 136453 2496 136465 2499
rect 130580 2468 136465 2496
rect 118007 2400 118556 2428
rect 118007 2397 118019 2400
rect 117961 2391 118019 2397
rect 119430 2388 119436 2440
rect 119488 2428 119494 2440
rect 121825 2431 121883 2437
rect 121825 2428 121837 2431
rect 119488 2400 121837 2428
rect 119488 2388 119494 2400
rect 121825 2397 121837 2400
rect 121871 2428 121883 2431
rect 123021 2431 123079 2437
rect 123021 2428 123033 2431
rect 121871 2400 123033 2428
rect 121871 2397 121883 2400
rect 121825 2391 121883 2397
rect 123021 2397 123033 2400
rect 123067 2397 123079 2431
rect 123021 2391 123079 2397
rect 125689 2431 125747 2437
rect 125689 2397 125701 2431
rect 125735 2428 125747 2431
rect 125735 2400 126284 2428
rect 125735 2397 125747 2400
rect 125689 2391 125747 2397
rect 104618 2360 104624 2372
rect 102060 2332 104624 2360
rect 99837 2323 99895 2329
rect 104618 2320 104624 2332
rect 104676 2360 104682 2372
rect 104989 2363 105047 2369
rect 104989 2360 105001 2363
rect 104676 2332 105001 2360
rect 104676 2320 104682 2332
rect 104989 2329 105001 2332
rect 105035 2329 105047 2363
rect 104989 2323 105047 2329
rect 107565 2363 107623 2369
rect 107565 2329 107577 2363
rect 107611 2329 107623 2363
rect 107565 2323 107623 2329
rect 94700 2264 99374 2292
rect 94593 2255 94651 2261
rect 99742 2252 99748 2304
rect 99800 2252 99806 2304
rect 104894 2252 104900 2304
rect 104952 2252 104958 2304
rect 106366 2252 106372 2304
rect 106424 2292 106430 2304
rect 107580 2292 107608 2323
rect 112346 2320 112352 2372
rect 112404 2360 112410 2372
rect 112717 2363 112775 2369
rect 112717 2360 112729 2363
rect 112404 2332 112729 2360
rect 112404 2320 112410 2332
rect 112717 2329 112729 2332
rect 112763 2329 112775 2363
rect 112717 2323 112775 2329
rect 115290 2320 115296 2372
rect 115348 2320 115354 2372
rect 120074 2320 120080 2372
rect 120132 2360 120138 2372
rect 120445 2363 120503 2369
rect 120445 2360 120457 2363
rect 120132 2332 120457 2360
rect 120132 2320 120138 2332
rect 120445 2329 120457 2332
rect 120491 2329 120503 2363
rect 120445 2323 120503 2329
rect 126256 2304 126284 2400
rect 128262 2388 128268 2440
rect 128320 2428 128326 2440
rect 130580 2428 130608 2468
rect 128320 2400 130608 2428
rect 128320 2388 128326 2400
rect 130654 2388 130660 2440
rect 130712 2428 130718 2440
rect 135824 2437 135852 2468
rect 136453 2465 136465 2468
rect 136499 2465 136511 2499
rect 150802 2496 150808 2508
rect 136453 2459 136511 2465
rect 137986 2468 150808 2496
rect 131301 2431 131359 2437
rect 131301 2428 131313 2431
rect 130712 2400 131313 2428
rect 130712 2388 130718 2400
rect 131301 2397 131313 2400
rect 131347 2397 131359 2431
rect 131301 2391 131359 2397
rect 133417 2431 133475 2437
rect 133417 2397 133429 2431
rect 133463 2428 133475 2431
rect 135809 2431 135867 2437
rect 133463 2400 134012 2428
rect 133463 2397 133475 2400
rect 133417 2391 133475 2397
rect 127066 2320 127072 2372
rect 127124 2360 127130 2372
rect 128170 2360 128176 2372
rect 127124 2332 128176 2360
rect 127124 2320 127130 2332
rect 128170 2320 128176 2332
rect 128228 2320 128234 2372
rect 128354 2320 128360 2372
rect 128412 2360 128418 2372
rect 128412 2332 133276 2360
rect 128412 2320 128418 2332
rect 106424 2264 107608 2292
rect 106424 2252 106430 2264
rect 107746 2252 107752 2304
rect 107804 2292 107810 2304
rect 109218 2292 109224 2304
rect 107804 2264 109224 2292
rect 107804 2252 107810 2264
rect 109218 2252 109224 2264
rect 109276 2252 109282 2304
rect 115198 2252 115204 2304
rect 115256 2252 115262 2304
rect 120350 2252 120356 2304
rect 120408 2252 120414 2304
rect 122926 2252 122932 2304
rect 122984 2252 122990 2304
rect 125502 2252 125508 2304
rect 125560 2252 125566 2304
rect 126238 2252 126244 2304
rect 126296 2252 126302 2304
rect 128078 2252 128084 2304
rect 128136 2252 128142 2304
rect 130838 2252 130844 2304
rect 130896 2252 130902 2304
rect 133248 2301 133276 2332
rect 133984 2304 134012 2400
rect 135809 2397 135821 2431
rect 135855 2397 135867 2431
rect 137986 2428 138014 2468
rect 150802 2456 150808 2468
rect 150860 2456 150866 2508
rect 153841 2499 153899 2505
rect 153841 2465 153853 2499
rect 153887 2496 153899 2499
rect 253934 2496 253940 2508
rect 153887 2468 253940 2496
rect 153887 2465 153899 2468
rect 153841 2459 153899 2465
rect 253934 2456 253940 2468
rect 253992 2456 253998 2508
rect 263410 2456 263416 2508
rect 263468 2496 263474 2508
rect 263468 2468 268056 2496
rect 263468 2456 263474 2468
rect 135809 2391 135867 2397
rect 136008 2400 138014 2428
rect 133233 2295 133291 2301
rect 133233 2261 133245 2295
rect 133279 2261 133291 2295
rect 133233 2255 133291 2261
rect 133966 2252 133972 2304
rect 134024 2252 134030 2304
rect 136008 2301 136036 2400
rect 138106 2388 138112 2440
rect 138164 2428 138170 2440
rect 138569 2431 138627 2437
rect 138569 2428 138581 2431
rect 138164 2400 138581 2428
rect 138164 2388 138170 2400
rect 138569 2397 138581 2400
rect 138615 2397 138627 2431
rect 138569 2391 138627 2397
rect 141142 2388 141148 2440
rect 141200 2388 141206 2440
rect 143074 2388 143080 2440
rect 143132 2428 143138 2440
rect 143721 2431 143779 2437
rect 143721 2428 143733 2431
rect 143132 2400 143733 2428
rect 143132 2388 143138 2400
rect 143721 2397 143733 2400
rect 143767 2397 143779 2431
rect 143721 2391 143779 2397
rect 146297 2431 146355 2437
rect 146297 2397 146309 2431
rect 146343 2397 146355 2431
rect 146297 2391 146355 2397
rect 138293 2363 138351 2369
rect 138293 2329 138305 2363
rect 138339 2360 138351 2363
rect 138339 2332 143396 2360
rect 138339 2329 138351 2332
rect 138293 2323 138351 2329
rect 135993 2295 136051 2301
rect 135993 2261 136005 2295
rect 136039 2261 136051 2295
rect 135993 2255 136051 2261
rect 136450 2252 136456 2304
rect 136508 2292 136514 2304
rect 140961 2295 141019 2301
rect 140961 2292 140973 2295
rect 136508 2264 140973 2292
rect 136508 2252 136514 2264
rect 140961 2261 140973 2264
rect 141007 2261 141019 2295
rect 143368 2292 143396 2332
rect 143442 2320 143448 2372
rect 143500 2320 143506 2372
rect 146312 2360 146340 2391
rect 148226 2388 148232 2440
rect 148284 2428 148290 2440
rect 148873 2431 148931 2437
rect 148873 2428 148885 2431
rect 148284 2400 148885 2428
rect 148284 2388 148290 2400
rect 148873 2397 148885 2400
rect 148919 2397 148931 2431
rect 148873 2391 148931 2397
rect 151449 2431 151507 2437
rect 151449 2397 151461 2431
rect 151495 2428 151507 2431
rect 151495 2400 152044 2428
rect 151495 2397 151507 2400
rect 151449 2391 151507 2397
rect 146846 2360 146852 2372
rect 144748 2332 146248 2360
rect 146312 2332 146852 2360
rect 144748 2292 144776 2332
rect 143368 2264 144776 2292
rect 140961 2255 141019 2261
rect 144914 2252 144920 2304
rect 144972 2292 144978 2304
rect 146113 2295 146171 2301
rect 146113 2292 146125 2295
rect 144972 2264 146125 2292
rect 144972 2252 144978 2264
rect 146113 2261 146125 2264
rect 146159 2261 146171 2295
rect 146220 2292 146248 2332
rect 146846 2320 146852 2332
rect 146904 2320 146910 2372
rect 148594 2320 148600 2372
rect 148652 2320 148658 2372
rect 152016 2304 152044 2400
rect 153378 2388 153384 2440
rect 153436 2428 153442 2440
rect 154025 2431 154083 2437
rect 154025 2428 154037 2431
rect 153436 2400 154037 2428
rect 153436 2388 153442 2400
rect 154025 2397 154037 2400
rect 154071 2397 154083 2431
rect 154025 2391 154083 2397
rect 156601 2431 156659 2437
rect 156601 2397 156613 2431
rect 156647 2428 156659 2431
rect 156647 2400 157196 2428
rect 156647 2397 156659 2400
rect 156601 2391 156659 2397
rect 157168 2304 157196 2400
rect 158898 2388 158904 2440
rect 158956 2388 158962 2440
rect 159177 2431 159235 2437
rect 159177 2397 159189 2431
rect 159223 2397 159235 2431
rect 159177 2391 159235 2397
rect 161753 2431 161811 2437
rect 161753 2397 161765 2431
rect 161799 2397 161811 2431
rect 161753 2391 161811 2397
rect 158530 2320 158536 2372
rect 158588 2360 158594 2372
rect 159192 2360 159220 2391
rect 158588 2332 159220 2360
rect 161768 2360 161796 2391
rect 161934 2388 161940 2440
rect 161992 2428 161998 2440
rect 166905 2431 166963 2437
rect 161992 2400 166764 2428
rect 161992 2388 161998 2400
rect 161768 2332 162348 2360
rect 158588 2320 158594 2332
rect 162320 2304 162348 2332
rect 163682 2320 163688 2372
rect 163740 2360 163746 2372
rect 164237 2363 164295 2369
rect 164237 2360 164249 2363
rect 163740 2332 164249 2360
rect 163740 2320 163746 2332
rect 164237 2329 164249 2332
rect 164283 2329 164295 2363
rect 164237 2323 164295 2329
rect 146662 2292 146668 2304
rect 146220 2264 146668 2292
rect 146113 2255 146171 2261
rect 146662 2252 146668 2264
rect 146720 2252 146726 2304
rect 151262 2252 151268 2304
rect 151320 2252 151326 2304
rect 151998 2252 152004 2304
rect 152056 2252 152062 2304
rect 156414 2252 156420 2304
rect 156472 2252 156478 2304
rect 157150 2252 157156 2304
rect 157208 2252 157214 2304
rect 161566 2252 161572 2304
rect 161624 2252 161630 2304
rect 162302 2252 162308 2304
rect 162360 2252 162366 2304
rect 164142 2252 164148 2304
rect 164200 2252 164206 2304
rect 166736 2301 166764 2400
rect 166905 2397 166917 2431
rect 166951 2397 166963 2431
rect 166905 2391 166963 2397
rect 172057 2431 172115 2437
rect 172057 2397 172069 2431
rect 172103 2428 172115 2431
rect 172103 2400 172652 2428
rect 172103 2397 172115 2400
rect 172057 2391 172115 2397
rect 166721 2295 166779 2301
rect 166721 2261 166733 2295
rect 166767 2261 166779 2295
rect 166920 2292 166948 2391
rect 168374 2320 168380 2372
rect 168432 2360 168438 2372
rect 169389 2363 169447 2369
rect 169389 2360 169401 2363
rect 168432 2332 169401 2360
rect 168432 2320 168438 2332
rect 169389 2329 169401 2332
rect 169435 2329 169447 2363
rect 169389 2323 169447 2329
rect 172624 2304 172652 2400
rect 177206 2388 177212 2440
rect 177264 2388 177270 2440
rect 179138 2388 179144 2440
rect 179196 2428 179202 2440
rect 179693 2431 179751 2437
rect 179693 2428 179705 2431
rect 179196 2400 179705 2428
rect 179196 2388 179202 2400
rect 179693 2397 179705 2400
rect 179739 2397 179751 2431
rect 179693 2391 179751 2397
rect 182361 2431 182419 2437
rect 182361 2397 182373 2431
rect 182407 2428 182419 2431
rect 182910 2428 182916 2440
rect 182407 2400 182916 2428
rect 182407 2397 182419 2400
rect 182361 2391 182419 2397
rect 182910 2388 182916 2400
rect 182968 2388 182974 2440
rect 184290 2388 184296 2440
rect 184348 2428 184354 2440
rect 187418 2428 187424 2440
rect 184348 2400 187424 2428
rect 184348 2388 184354 2400
rect 187418 2388 187424 2400
rect 187476 2388 187482 2440
rect 187513 2431 187571 2437
rect 187513 2397 187525 2431
rect 187559 2428 187571 2431
rect 188062 2428 188068 2440
rect 187559 2400 188068 2428
rect 187559 2397 187571 2400
rect 187513 2391 187571 2397
rect 188062 2388 188068 2400
rect 188120 2388 188126 2440
rect 191742 2428 191748 2440
rect 188172 2400 191748 2428
rect 173986 2320 173992 2372
rect 174044 2360 174050 2372
rect 174541 2363 174599 2369
rect 174541 2360 174553 2363
rect 174044 2332 174553 2360
rect 174044 2320 174050 2332
rect 174541 2329 174553 2332
rect 174587 2329 174599 2363
rect 174541 2323 174599 2329
rect 174998 2320 175004 2372
rect 175056 2360 175062 2372
rect 183554 2360 183560 2372
rect 175056 2332 183560 2360
rect 175056 2320 175062 2332
rect 183554 2320 183560 2332
rect 183612 2360 183618 2372
rect 184845 2363 184903 2369
rect 184845 2360 184857 2363
rect 183612 2332 184857 2360
rect 183612 2320 183618 2332
rect 184845 2329 184857 2332
rect 184891 2329 184903 2363
rect 184845 2323 184903 2329
rect 185486 2320 185492 2372
rect 185544 2360 185550 2372
rect 186774 2360 186780 2372
rect 185544 2332 186780 2360
rect 185544 2320 185550 2332
rect 186774 2320 186780 2332
rect 186832 2320 186838 2372
rect 186866 2320 186872 2372
rect 186924 2360 186930 2372
rect 188172 2360 188200 2400
rect 191742 2388 191748 2400
rect 191800 2388 191806 2440
rect 192665 2431 192723 2437
rect 192665 2397 192677 2431
rect 192711 2428 192723 2431
rect 193214 2428 193220 2440
rect 192711 2400 193220 2428
rect 192711 2397 192723 2400
rect 192665 2391 192723 2397
rect 193214 2388 193220 2400
rect 193272 2388 193278 2440
rect 195146 2388 195152 2440
rect 195204 2388 195210 2440
rect 197814 2388 197820 2440
rect 197872 2428 197878 2440
rect 198277 2431 198335 2437
rect 198277 2428 198289 2431
rect 197872 2400 198289 2428
rect 197872 2388 197878 2400
rect 198277 2397 198289 2400
rect 198323 2397 198335 2431
rect 198277 2391 198335 2397
rect 200022 2388 200028 2440
rect 200080 2428 200086 2440
rect 200393 2431 200451 2437
rect 200393 2428 200405 2431
rect 200080 2400 200405 2428
rect 200080 2388 200114 2400
rect 200393 2397 200405 2400
rect 200439 2397 200451 2431
rect 200393 2391 200451 2397
rect 202969 2431 203027 2437
rect 202969 2397 202981 2431
rect 203015 2428 203027 2431
rect 203058 2428 203064 2440
rect 203015 2400 203064 2428
rect 203015 2397 203027 2400
rect 202969 2391 203027 2397
rect 203058 2388 203064 2400
rect 203116 2428 203122 2440
rect 203429 2431 203487 2437
rect 203429 2428 203441 2431
rect 203116 2400 203441 2428
rect 203116 2388 203122 2400
rect 203429 2397 203441 2400
rect 203475 2397 203487 2431
rect 203429 2391 203487 2397
rect 205082 2388 205088 2440
rect 205140 2428 205146 2440
rect 205545 2431 205603 2437
rect 205545 2428 205557 2431
rect 205140 2400 205557 2428
rect 205140 2388 205146 2400
rect 205545 2397 205557 2400
rect 205591 2397 205603 2431
rect 205545 2391 205603 2397
rect 208121 2431 208179 2437
rect 208121 2397 208133 2431
rect 208167 2428 208179 2431
rect 208578 2428 208584 2440
rect 208167 2400 208584 2428
rect 208167 2397 208179 2400
rect 208121 2391 208179 2397
rect 208578 2388 208584 2400
rect 208636 2388 208642 2440
rect 210234 2388 210240 2440
rect 210292 2428 210298 2440
rect 210697 2431 210755 2437
rect 210697 2428 210709 2431
rect 210292 2400 210709 2428
rect 210292 2388 210298 2400
rect 210697 2397 210709 2400
rect 210743 2397 210755 2431
rect 210697 2391 210755 2397
rect 213270 2388 213276 2440
rect 213328 2428 213334 2440
rect 213733 2431 213791 2437
rect 213733 2428 213745 2431
rect 213328 2400 213745 2428
rect 213328 2388 213334 2400
rect 213733 2397 213745 2400
rect 213779 2397 213791 2431
rect 213733 2391 213791 2397
rect 215386 2388 215392 2440
rect 215444 2428 215450 2440
rect 215849 2431 215907 2437
rect 215849 2428 215861 2431
rect 215444 2400 215861 2428
rect 215444 2388 215450 2400
rect 215849 2397 215861 2400
rect 215895 2397 215907 2431
rect 215849 2391 215907 2397
rect 218422 2388 218428 2440
rect 218480 2428 218486 2440
rect 218885 2431 218943 2437
rect 218885 2428 218897 2431
rect 218480 2400 218897 2428
rect 218480 2388 218486 2400
rect 218885 2397 218897 2400
rect 218931 2397 218943 2431
rect 218885 2391 218943 2397
rect 220538 2388 220544 2440
rect 220596 2428 220602 2440
rect 221001 2431 221059 2437
rect 221001 2428 221013 2431
rect 220596 2400 221013 2428
rect 220596 2388 220602 2400
rect 221001 2397 221013 2400
rect 221047 2397 221059 2431
rect 221001 2391 221059 2397
rect 223577 2431 223635 2437
rect 223577 2397 223589 2431
rect 223623 2428 223635 2431
rect 224126 2428 224132 2440
rect 223623 2400 224132 2428
rect 223623 2397 223635 2400
rect 223577 2391 223635 2397
rect 224126 2388 224132 2400
rect 224184 2388 224190 2440
rect 228729 2431 228787 2437
rect 228729 2397 228741 2431
rect 228775 2428 228787 2431
rect 229186 2428 229192 2440
rect 228775 2400 229192 2428
rect 228775 2397 228787 2400
rect 228729 2391 228787 2397
rect 229186 2388 229192 2400
rect 229244 2388 229250 2440
rect 231305 2431 231363 2437
rect 231305 2397 231317 2431
rect 231351 2428 231363 2431
rect 231854 2428 231860 2440
rect 231351 2400 231860 2428
rect 231351 2397 231363 2400
rect 231305 2391 231363 2397
rect 231854 2388 231860 2400
rect 231912 2388 231918 2440
rect 233881 2431 233939 2437
rect 233881 2397 233893 2431
rect 233927 2428 233939 2431
rect 234430 2428 234436 2440
rect 233927 2400 234436 2428
rect 233927 2397 233939 2400
rect 233881 2391 233939 2397
rect 234430 2388 234436 2400
rect 234488 2388 234494 2440
rect 236457 2431 236515 2437
rect 236457 2397 236469 2431
rect 236503 2428 236515 2431
rect 237006 2428 237012 2440
rect 236503 2400 237012 2428
rect 236503 2397 236515 2400
rect 236457 2391 236515 2397
rect 237006 2388 237012 2400
rect 237064 2388 237070 2440
rect 239030 2388 239036 2440
rect 239088 2428 239094 2440
rect 239493 2431 239551 2437
rect 239493 2428 239505 2431
rect 239088 2400 239505 2428
rect 239088 2388 239094 2400
rect 239493 2397 239505 2400
rect 239539 2397 239551 2431
rect 239493 2391 239551 2397
rect 241609 2431 241667 2437
rect 241609 2397 241621 2431
rect 241655 2428 241667 2431
rect 242158 2428 242164 2440
rect 241655 2400 242164 2428
rect 241655 2397 241667 2400
rect 241609 2391 241667 2397
rect 242158 2388 242164 2400
rect 242216 2388 242222 2440
rect 244185 2431 244243 2437
rect 244185 2397 244197 2431
rect 244231 2428 244243 2431
rect 244826 2428 244832 2440
rect 244231 2400 244832 2428
rect 244231 2397 244243 2400
rect 244185 2391 244243 2397
rect 244826 2388 244832 2400
rect 244884 2388 244890 2440
rect 246761 2431 246819 2437
rect 246761 2397 246773 2431
rect 246807 2428 246819 2431
rect 247218 2428 247224 2440
rect 246807 2400 247224 2428
rect 246807 2397 246819 2400
rect 246761 2391 246819 2397
rect 247218 2388 247224 2400
rect 247276 2388 247282 2440
rect 249337 2431 249395 2437
rect 249337 2397 249349 2431
rect 249383 2428 249395 2431
rect 249886 2428 249892 2440
rect 249383 2400 249892 2428
rect 249383 2397 249395 2400
rect 249337 2391 249395 2397
rect 249886 2388 249892 2400
rect 249944 2388 249950 2440
rect 251910 2388 251916 2440
rect 251968 2428 251974 2440
rect 252373 2431 252431 2437
rect 252373 2428 252385 2431
rect 251968 2400 252385 2428
rect 251968 2388 251974 2400
rect 252373 2397 252385 2400
rect 252419 2397 252431 2431
rect 252373 2391 252431 2397
rect 254489 2431 254547 2437
rect 254489 2397 254501 2431
rect 254535 2428 254547 2431
rect 257065 2431 257123 2437
rect 254535 2400 255084 2428
rect 254535 2397 254547 2400
rect 254489 2391 254547 2397
rect 186924 2332 188200 2360
rect 186924 2320 186930 2332
rect 189074 2320 189080 2372
rect 189132 2360 189138 2372
rect 189997 2363 190055 2369
rect 189997 2360 190009 2363
rect 189132 2332 190009 2360
rect 189132 2320 189138 2332
rect 189997 2329 190009 2332
rect 190043 2329 190055 2363
rect 195330 2360 195336 2372
rect 189997 2323 190055 2329
rect 192404 2332 195336 2360
rect 167454 2292 167460 2304
rect 166920 2264 167460 2292
rect 166721 2255 166779 2261
rect 167454 2252 167460 2264
rect 167512 2252 167518 2304
rect 169294 2252 169300 2304
rect 169352 2252 169358 2304
rect 171134 2252 171140 2304
rect 171192 2292 171198 2304
rect 171873 2295 171931 2301
rect 171873 2292 171885 2295
rect 171192 2264 171885 2292
rect 171192 2252 171198 2264
rect 171873 2261 171885 2264
rect 171919 2261 171931 2295
rect 171873 2255 171931 2261
rect 172606 2252 172612 2304
rect 172664 2252 172670 2304
rect 174446 2252 174452 2304
rect 174504 2252 174510 2304
rect 174630 2252 174636 2304
rect 174688 2292 174694 2304
rect 177025 2295 177083 2301
rect 177025 2292 177037 2295
rect 174688 2264 177037 2292
rect 174688 2252 174694 2264
rect 177025 2261 177037 2264
rect 177071 2261 177083 2295
rect 177025 2255 177083 2261
rect 179598 2252 179604 2304
rect 179656 2252 179662 2304
rect 182174 2252 182180 2304
rect 182232 2252 182238 2304
rect 183646 2252 183652 2304
rect 183704 2292 183710 2304
rect 187329 2295 187387 2301
rect 187329 2292 187341 2295
rect 183704 2264 187341 2292
rect 183704 2252 183710 2264
rect 187329 2261 187341 2264
rect 187375 2261 187387 2295
rect 187329 2255 187387 2261
rect 189905 2295 189963 2301
rect 189905 2261 189917 2295
rect 189951 2292 189963 2295
rect 192404 2292 192432 2332
rect 195330 2320 195336 2332
rect 195388 2320 195394 2372
rect 200086 2360 200114 2388
rect 195440 2332 200114 2360
rect 189951 2264 192432 2292
rect 189951 2261 189963 2264
rect 189905 2255 189963 2261
rect 195054 2252 195060 2304
rect 195112 2252 195118 2304
rect 195146 2252 195152 2304
rect 195204 2292 195210 2304
rect 195440 2292 195468 2332
rect 226058 2320 226064 2372
rect 226116 2320 226122 2372
rect 233234 2320 233240 2372
rect 233292 2360 233298 2372
rect 233292 2332 238892 2360
rect 233292 2320 233298 2332
rect 195204 2264 195468 2292
rect 195204 2252 195210 2264
rect 195974 2252 195980 2304
rect 196032 2292 196038 2304
rect 197633 2295 197691 2301
rect 197633 2292 197645 2295
rect 196032 2264 197645 2292
rect 196032 2252 196038 2264
rect 197633 2261 197645 2264
rect 197679 2261 197691 2295
rect 197633 2255 197691 2261
rect 200206 2252 200212 2304
rect 200264 2252 200270 2304
rect 202782 2252 202788 2304
rect 202840 2252 202846 2304
rect 207934 2252 207940 2304
rect 207992 2252 207998 2304
rect 213086 2252 213092 2304
rect 213144 2252 213150 2304
rect 215662 2252 215668 2304
rect 215720 2252 215726 2304
rect 218238 2252 218244 2304
rect 218296 2252 218302 2304
rect 220814 2252 220820 2304
rect 220872 2252 220878 2304
rect 223390 2252 223396 2304
rect 223448 2252 223454 2304
rect 225966 2252 225972 2304
rect 226024 2252 226030 2304
rect 228542 2252 228548 2304
rect 228600 2252 228606 2304
rect 229094 2252 229100 2304
rect 229152 2292 229158 2304
rect 231121 2295 231179 2301
rect 231121 2292 231133 2295
rect 229152 2264 231133 2292
rect 229152 2252 229158 2264
rect 231121 2261 231133 2264
rect 231167 2261 231179 2295
rect 231121 2255 231179 2261
rect 233694 2252 233700 2304
rect 233752 2252 233758 2304
rect 236270 2252 236276 2304
rect 236328 2252 236334 2304
rect 238864 2301 238892 2332
rect 243906 2320 243912 2372
rect 243964 2360 243970 2372
rect 243964 2332 251174 2360
rect 243964 2320 243970 2332
rect 238849 2295 238907 2301
rect 238849 2261 238861 2295
rect 238895 2261 238907 2295
rect 238849 2255 238907 2261
rect 241422 2252 241428 2304
rect 241480 2252 241486 2304
rect 242894 2252 242900 2304
rect 242952 2292 242958 2304
rect 244001 2295 244059 2301
rect 244001 2292 244013 2295
rect 242952 2264 244013 2292
rect 242952 2252 242958 2264
rect 244001 2261 244013 2264
rect 244047 2261 244059 2295
rect 244001 2255 244059 2261
rect 244090 2252 244096 2304
rect 244148 2292 244154 2304
rect 246577 2295 246635 2301
rect 246577 2292 246589 2295
rect 244148 2264 246589 2292
rect 244148 2252 244154 2264
rect 246577 2261 246589 2264
rect 246623 2261 246635 2295
rect 246577 2255 246635 2261
rect 247034 2252 247040 2304
rect 247092 2292 247098 2304
rect 249153 2295 249211 2301
rect 249153 2292 249165 2295
rect 247092 2264 249165 2292
rect 247092 2252 247098 2264
rect 249153 2261 249165 2264
rect 249199 2261 249211 2295
rect 251146 2292 251174 2332
rect 255056 2304 255084 2400
rect 257065 2397 257077 2431
rect 257111 2428 257123 2431
rect 257614 2428 257620 2440
rect 257111 2400 257620 2428
rect 257111 2397 257123 2400
rect 257065 2391 257123 2397
rect 257614 2388 257620 2400
rect 257672 2388 257678 2440
rect 259641 2431 259699 2437
rect 259641 2397 259653 2431
rect 259687 2428 259699 2431
rect 260190 2428 260196 2440
rect 259687 2400 260196 2428
rect 259687 2397 259699 2400
rect 259641 2391 259699 2397
rect 260190 2388 260196 2400
rect 260248 2388 260254 2440
rect 262214 2388 262220 2440
rect 262272 2428 262278 2440
rect 262677 2431 262735 2437
rect 262677 2428 262689 2431
rect 262272 2400 262689 2428
rect 262272 2388 262278 2400
rect 262677 2397 262689 2400
rect 262723 2397 262735 2431
rect 262677 2391 262735 2397
rect 264793 2431 264851 2437
rect 264793 2397 264805 2431
rect 264839 2428 264851 2431
rect 265342 2428 265348 2440
rect 264839 2400 265348 2428
rect 264839 2397 264851 2400
rect 264793 2391 264851 2397
rect 265342 2388 265348 2400
rect 265400 2388 265406 2440
rect 267369 2431 267427 2437
rect 267369 2397 267381 2431
rect 267415 2428 267427 2431
rect 267415 2400 267964 2428
rect 267415 2397 267427 2400
rect 267369 2391 267427 2397
rect 267936 2304 267964 2400
rect 268028 2360 268056 2468
rect 291746 2456 291752 2508
rect 291804 2496 291810 2508
rect 295628 2496 295656 2536
rect 300673 2533 300685 2536
rect 300719 2533 300731 2567
rect 300673 2527 300731 2533
rect 291804 2468 295656 2496
rect 291804 2456 291810 2468
rect 298186 2456 298192 2508
rect 298244 2496 298250 2508
rect 302206 2496 302234 2604
rect 303249 2601 303261 2604
rect 303295 2601 303307 2635
rect 303249 2595 303307 2601
rect 303982 2592 303988 2644
rect 304040 2592 304046 2644
rect 306558 2592 306564 2644
rect 306616 2592 306622 2644
rect 309134 2592 309140 2644
rect 309192 2592 309198 2644
rect 316865 2635 316923 2641
rect 316865 2601 316877 2635
rect 316911 2632 316923 2635
rect 319254 2632 319260 2644
rect 316911 2604 319260 2632
rect 316911 2601 316923 2604
rect 316865 2595 316923 2601
rect 303522 2524 303528 2576
rect 303580 2564 303586 2576
rect 308401 2567 308459 2573
rect 308401 2564 308413 2567
rect 303580 2536 308413 2564
rect 303580 2524 303586 2536
rect 308401 2533 308413 2536
rect 308447 2533 308459 2567
rect 313553 2567 313611 2573
rect 313553 2564 313565 2567
rect 308401 2527 308459 2533
rect 308508 2536 313565 2564
rect 298244 2468 302234 2496
rect 298244 2456 298250 2468
rect 306374 2456 306380 2508
rect 306432 2496 306438 2508
rect 308508 2496 308536 2536
rect 313553 2533 313565 2536
rect 313599 2533 313611 2567
rect 316880 2564 316908 2595
rect 319254 2592 319260 2604
rect 319312 2592 319318 2644
rect 322014 2592 322020 2644
rect 322072 2592 322078 2644
rect 327169 2635 327227 2641
rect 327169 2601 327181 2635
rect 327215 2632 327227 2635
rect 327215 2604 357434 2632
rect 327215 2601 327227 2604
rect 327169 2595 327227 2601
rect 313553 2527 313611 2533
rect 316420 2536 316908 2564
rect 311713 2499 311771 2505
rect 311713 2496 311725 2499
rect 306432 2468 308536 2496
rect 311176 2468 311725 2496
rect 306432 2456 306438 2468
rect 269945 2431 270003 2437
rect 269945 2397 269957 2431
rect 269991 2428 270003 2431
rect 270494 2428 270500 2440
rect 269991 2400 270500 2428
rect 269991 2397 270003 2400
rect 269945 2391 270003 2397
rect 270494 2388 270500 2400
rect 270552 2388 270558 2440
rect 272521 2431 272579 2437
rect 272521 2397 272533 2431
rect 272567 2428 272579 2431
rect 273070 2428 273076 2440
rect 272567 2400 273076 2428
rect 272567 2397 272579 2400
rect 272521 2391 272579 2397
rect 273070 2388 273076 2400
rect 273128 2388 273134 2440
rect 275097 2431 275155 2437
rect 275097 2397 275109 2431
rect 275143 2428 275155 2431
rect 275646 2428 275652 2440
rect 275143 2400 275652 2428
rect 275143 2397 275155 2400
rect 275097 2391 275155 2397
rect 275646 2388 275652 2400
rect 275704 2388 275710 2440
rect 277673 2431 277731 2437
rect 277673 2397 277685 2431
rect 277719 2428 277731 2431
rect 280249 2431 280307 2437
rect 277719 2400 278268 2428
rect 277719 2397 277731 2400
rect 277673 2391 277731 2397
rect 268028 2332 273254 2360
rect 251729 2295 251787 2301
rect 251729 2292 251741 2295
rect 251146 2264 251741 2292
rect 249153 2255 249211 2261
rect 251729 2261 251741 2264
rect 251775 2261 251787 2295
rect 251729 2255 251787 2261
rect 253842 2252 253848 2304
rect 253900 2292 253906 2304
rect 254305 2295 254363 2301
rect 254305 2292 254317 2295
rect 253900 2264 254317 2292
rect 253900 2252 253906 2264
rect 254305 2261 254317 2264
rect 254351 2261 254363 2295
rect 254305 2255 254363 2261
rect 255038 2252 255044 2304
rect 255096 2252 255102 2304
rect 255406 2252 255412 2304
rect 255464 2292 255470 2304
rect 256881 2295 256939 2301
rect 256881 2292 256893 2295
rect 255464 2264 256893 2292
rect 255464 2252 255470 2264
rect 256881 2261 256893 2264
rect 256927 2261 256939 2295
rect 256881 2255 256939 2261
rect 258074 2252 258080 2304
rect 258132 2292 258138 2304
rect 259457 2295 259515 2301
rect 259457 2292 259469 2295
rect 258132 2264 259469 2292
rect 258132 2252 258138 2264
rect 259457 2261 259469 2264
rect 259503 2261 259515 2295
rect 259457 2255 259515 2261
rect 260834 2252 260840 2304
rect 260892 2292 260898 2304
rect 262033 2295 262091 2301
rect 262033 2292 262045 2295
rect 260892 2264 262045 2292
rect 260892 2252 260898 2264
rect 262033 2261 262045 2264
rect 262079 2261 262091 2295
rect 262033 2255 262091 2261
rect 263594 2252 263600 2304
rect 263652 2292 263658 2304
rect 264609 2295 264667 2301
rect 264609 2292 264621 2295
rect 263652 2264 264621 2292
rect 263652 2252 263658 2264
rect 264609 2261 264621 2264
rect 264655 2261 264667 2295
rect 264609 2255 264667 2261
rect 267182 2252 267188 2304
rect 267240 2252 267246 2304
rect 267918 2252 267924 2304
rect 267976 2252 267982 2304
rect 268010 2252 268016 2304
rect 268068 2292 268074 2304
rect 269761 2295 269819 2301
rect 269761 2292 269773 2295
rect 268068 2264 269773 2292
rect 268068 2252 268074 2264
rect 269761 2261 269773 2264
rect 269807 2261 269819 2295
rect 269761 2255 269819 2261
rect 269850 2252 269856 2304
rect 269908 2292 269914 2304
rect 272337 2295 272395 2301
rect 272337 2292 272349 2295
rect 269908 2264 272349 2292
rect 269908 2252 269914 2264
rect 272337 2261 272349 2264
rect 272383 2261 272395 2295
rect 273226 2292 273254 2332
rect 278240 2304 278268 2400
rect 280249 2397 280261 2431
rect 280295 2428 280307 2431
rect 280798 2428 280804 2440
rect 280295 2400 280804 2428
rect 280295 2397 280307 2400
rect 280249 2391 280307 2397
rect 280798 2388 280804 2400
rect 280856 2388 280862 2440
rect 282825 2431 282883 2437
rect 282825 2397 282837 2431
rect 282871 2428 282883 2431
rect 283374 2428 283380 2440
rect 282871 2400 283380 2428
rect 282871 2397 282883 2400
rect 282825 2391 282883 2397
rect 283374 2388 283380 2400
rect 283432 2388 283438 2440
rect 285401 2431 285459 2437
rect 285401 2397 285413 2431
rect 285447 2428 285459 2431
rect 285950 2428 285956 2440
rect 285447 2400 285956 2428
rect 285447 2397 285459 2400
rect 285401 2391 285459 2397
rect 285950 2388 285956 2400
rect 286008 2388 286014 2440
rect 287977 2431 288035 2437
rect 287977 2397 287989 2431
rect 288023 2428 288035 2431
rect 288526 2428 288532 2440
rect 288023 2400 288532 2428
rect 288023 2397 288035 2400
rect 287977 2391 288035 2397
rect 288526 2388 288532 2400
rect 288584 2388 288590 2440
rect 290553 2431 290611 2437
rect 290553 2397 290565 2431
rect 290599 2428 290611 2431
rect 291102 2428 291108 2440
rect 290599 2400 291108 2428
rect 290599 2397 290611 2400
rect 290553 2391 290611 2397
rect 291102 2388 291108 2400
rect 291160 2388 291166 2440
rect 293129 2431 293187 2437
rect 293129 2397 293141 2431
rect 293175 2428 293187 2431
rect 293678 2428 293684 2440
rect 293175 2400 293684 2428
rect 293175 2397 293187 2400
rect 293129 2391 293187 2397
rect 293678 2388 293684 2400
rect 293736 2388 293742 2440
rect 295705 2431 295763 2437
rect 295705 2397 295717 2431
rect 295751 2428 295763 2431
rect 296254 2428 296260 2440
rect 295751 2400 296260 2428
rect 295751 2397 295763 2400
rect 295705 2391 295763 2397
rect 296254 2388 296260 2400
rect 296312 2388 296318 2440
rect 298281 2431 298339 2437
rect 298281 2397 298293 2431
rect 298327 2428 298339 2431
rect 298830 2428 298836 2440
rect 298327 2400 298836 2428
rect 298327 2397 298339 2400
rect 298281 2391 298339 2397
rect 298830 2388 298836 2400
rect 298888 2388 298894 2440
rect 300857 2431 300915 2437
rect 300857 2397 300869 2431
rect 300903 2428 300915 2431
rect 301406 2428 301412 2440
rect 300903 2400 301412 2428
rect 300903 2397 300915 2400
rect 300857 2391 300915 2397
rect 301406 2388 301412 2400
rect 301464 2388 301470 2440
rect 303433 2431 303491 2437
rect 303433 2397 303445 2431
rect 303479 2428 303491 2431
rect 303982 2428 303988 2440
rect 303479 2400 303988 2428
rect 303479 2397 303491 2400
rect 303433 2391 303491 2397
rect 303982 2388 303988 2400
rect 304040 2388 304046 2440
rect 306009 2431 306067 2437
rect 306009 2397 306021 2431
rect 306055 2428 306067 2431
rect 306558 2428 306564 2440
rect 306055 2400 306564 2428
rect 306055 2397 306067 2400
rect 306009 2391 306067 2397
rect 306558 2388 306564 2400
rect 306616 2388 306622 2440
rect 308585 2431 308643 2437
rect 308585 2397 308597 2431
rect 308631 2428 308643 2431
rect 309134 2428 309140 2440
rect 308631 2400 309140 2428
rect 308631 2397 308643 2400
rect 308585 2391 308643 2397
rect 309134 2388 309140 2400
rect 309192 2388 309198 2440
rect 311176 2437 311204 2468
rect 311713 2465 311725 2468
rect 311759 2496 311771 2499
rect 316420 2496 316448 2536
rect 311759 2468 316264 2496
rect 311759 2465 311771 2468
rect 311713 2459 311771 2465
rect 311161 2431 311219 2437
rect 311161 2397 311173 2431
rect 311207 2397 311219 2431
rect 311161 2391 311219 2397
rect 313737 2431 313795 2437
rect 313737 2397 313749 2431
rect 313783 2428 313795 2431
rect 314286 2428 314292 2440
rect 313783 2400 314292 2428
rect 313783 2397 313795 2400
rect 313737 2391 313795 2397
rect 314286 2388 314292 2400
rect 314344 2388 314350 2440
rect 302694 2320 302700 2372
rect 302752 2360 302758 2372
rect 302752 2332 309134 2360
rect 302752 2320 302758 2332
rect 274913 2295 274971 2301
rect 274913 2292 274925 2295
rect 273226 2264 274925 2292
rect 272337 2255 272395 2261
rect 274913 2261 274925 2264
rect 274959 2261 274971 2295
rect 274913 2255 274971 2261
rect 276014 2252 276020 2304
rect 276072 2292 276078 2304
rect 277489 2295 277547 2301
rect 277489 2292 277501 2295
rect 276072 2264 277501 2292
rect 276072 2252 276078 2264
rect 277489 2261 277501 2264
rect 277535 2261 277547 2295
rect 277489 2255 277547 2261
rect 278222 2252 278228 2304
rect 278280 2252 278286 2304
rect 278774 2252 278780 2304
rect 278832 2292 278838 2304
rect 280065 2295 280123 2301
rect 280065 2292 280077 2295
rect 278832 2264 280077 2292
rect 278832 2252 278838 2264
rect 280065 2261 280077 2264
rect 280111 2261 280123 2295
rect 280065 2255 280123 2261
rect 282638 2252 282644 2304
rect 282696 2252 282702 2304
rect 282730 2252 282736 2304
rect 282788 2292 282794 2304
rect 285217 2295 285275 2301
rect 285217 2292 285229 2295
rect 282788 2264 285229 2292
rect 282788 2252 282794 2264
rect 285217 2261 285229 2264
rect 285263 2261 285275 2295
rect 285217 2255 285275 2261
rect 285674 2252 285680 2304
rect 285732 2292 285738 2304
rect 287793 2295 287851 2301
rect 287793 2292 287805 2295
rect 285732 2264 287805 2292
rect 285732 2252 285738 2264
rect 287793 2261 287805 2264
rect 287839 2261 287851 2295
rect 287793 2255 287851 2261
rect 289906 2252 289912 2304
rect 289964 2292 289970 2304
rect 292945 2295 293003 2301
rect 292945 2292 292957 2295
rect 289964 2264 292957 2292
rect 289964 2252 289970 2264
rect 292945 2261 292957 2264
rect 292991 2261 293003 2295
rect 292945 2255 293003 2261
rect 295242 2252 295248 2304
rect 295300 2292 295306 2304
rect 298097 2295 298155 2301
rect 298097 2292 298109 2295
rect 295300 2264 298109 2292
rect 295300 2252 295306 2264
rect 298097 2261 298109 2264
rect 298143 2261 298155 2295
rect 298097 2255 298155 2261
rect 300854 2252 300860 2304
rect 300912 2292 300918 2304
rect 305825 2295 305883 2301
rect 305825 2292 305837 2295
rect 300912 2264 305837 2292
rect 300912 2252 300918 2264
rect 305825 2261 305837 2264
rect 305871 2261 305883 2295
rect 309106 2292 309134 2332
rect 309226 2320 309232 2372
rect 309284 2360 309290 2372
rect 316236 2360 316264 2468
rect 316328 2468 316448 2496
rect 316972 2468 325694 2496
rect 316328 2437 316356 2468
rect 316313 2431 316371 2437
rect 316313 2397 316325 2431
rect 316359 2397 316371 2431
rect 316972 2428 317000 2468
rect 316313 2391 316371 2397
rect 316420 2400 317000 2428
rect 318889 2431 318947 2437
rect 316420 2360 316448 2400
rect 318889 2397 318901 2431
rect 318935 2428 318947 2431
rect 319438 2428 319444 2440
rect 318935 2400 319444 2428
rect 318935 2397 318947 2400
rect 318889 2391 318947 2397
rect 319438 2388 319444 2400
rect 319496 2388 319502 2440
rect 321465 2431 321523 2437
rect 321465 2397 321477 2431
rect 321511 2428 321523 2431
rect 322014 2428 322020 2440
rect 321511 2400 322020 2428
rect 321511 2397 321523 2400
rect 321465 2391 321523 2397
rect 322014 2388 322020 2400
rect 322072 2388 322078 2440
rect 324041 2431 324099 2437
rect 324041 2397 324053 2431
rect 324087 2428 324099 2431
rect 324087 2400 324636 2428
rect 324087 2397 324099 2400
rect 324041 2391 324099 2397
rect 309284 2332 316172 2360
rect 316236 2332 316448 2360
rect 309284 2320 309290 2332
rect 310977 2295 311035 2301
rect 310977 2292 310989 2295
rect 309106 2264 310989 2292
rect 305825 2255 305883 2261
rect 310977 2261 310989 2264
rect 311023 2261 311035 2295
rect 310977 2255 311035 2261
rect 314286 2252 314292 2304
rect 314344 2252 314350 2304
rect 316144 2301 316172 2332
rect 316678 2320 316684 2372
rect 316736 2360 316742 2372
rect 316736 2332 323900 2360
rect 316736 2320 316742 2332
rect 316129 2295 316187 2301
rect 316129 2261 316141 2295
rect 316175 2261 316187 2295
rect 316129 2255 316187 2261
rect 318702 2252 318708 2304
rect 318760 2252 318766 2304
rect 319438 2252 319444 2304
rect 319496 2252 319502 2304
rect 321278 2252 321284 2304
rect 321336 2252 321342 2304
rect 323872 2301 323900 2332
rect 324608 2304 324636 2400
rect 325666 2360 325694 2468
rect 326617 2431 326675 2437
rect 326617 2397 326629 2431
rect 326663 2428 326675 2431
rect 327184 2428 327212 2595
rect 334894 2524 334900 2576
rect 334952 2524 334958 2576
rect 347777 2567 347835 2573
rect 347777 2533 347789 2567
rect 347823 2564 347835 2567
rect 349062 2564 349068 2576
rect 347823 2536 349068 2564
rect 347823 2533 347835 2536
rect 347777 2527 347835 2533
rect 326663 2400 327212 2428
rect 329193 2431 329251 2437
rect 326663 2397 326675 2400
rect 326617 2391 326675 2397
rect 329193 2397 329205 2431
rect 329239 2428 329251 2431
rect 329742 2428 329748 2440
rect 329239 2400 329748 2428
rect 329239 2397 329251 2400
rect 329193 2391 329251 2397
rect 329742 2388 329748 2400
rect 329800 2388 329806 2440
rect 331769 2431 331827 2437
rect 331769 2397 331781 2431
rect 331815 2428 331827 2431
rect 332318 2428 332324 2440
rect 331815 2400 332324 2428
rect 331815 2397 331827 2400
rect 331769 2391 331827 2397
rect 332318 2388 332324 2400
rect 332376 2388 332382 2440
rect 334345 2431 334403 2437
rect 334345 2397 334357 2431
rect 334391 2428 334403 2431
rect 334912 2428 334940 2524
rect 334391 2400 334940 2428
rect 336921 2431 336979 2437
rect 334391 2397 334403 2400
rect 334345 2391 334403 2397
rect 336921 2397 336933 2431
rect 336967 2428 336979 2431
rect 337470 2428 337476 2440
rect 336967 2400 337476 2428
rect 336967 2397 336979 2400
rect 336921 2391 336979 2397
rect 337470 2388 337476 2400
rect 337528 2388 337534 2440
rect 339497 2431 339555 2437
rect 339497 2397 339509 2431
rect 339543 2428 339555 2431
rect 340046 2428 340052 2440
rect 339543 2400 340052 2428
rect 339543 2397 339555 2400
rect 339497 2391 339555 2397
rect 340046 2388 340052 2400
rect 340104 2388 340110 2440
rect 342073 2431 342131 2437
rect 342073 2397 342085 2431
rect 342119 2428 342131 2431
rect 342622 2428 342628 2440
rect 342119 2400 342628 2428
rect 342119 2397 342131 2400
rect 342073 2391 342131 2397
rect 342622 2388 342628 2400
rect 342680 2388 342686 2440
rect 344649 2431 344707 2437
rect 344649 2397 344661 2431
rect 344695 2428 344707 2431
rect 345198 2428 345204 2440
rect 344695 2400 345204 2428
rect 344695 2397 344707 2400
rect 344649 2391 344707 2397
rect 345198 2388 345204 2400
rect 345256 2388 345262 2440
rect 347225 2431 347283 2437
rect 347225 2397 347237 2431
rect 347271 2428 347283 2431
rect 347792 2428 347820 2527
rect 349062 2524 349068 2536
rect 349120 2524 349126 2576
rect 349617 2567 349675 2573
rect 349617 2533 349629 2567
rect 349663 2564 349675 2567
rect 355410 2564 355416 2576
rect 349663 2536 355416 2564
rect 349663 2533 349675 2536
rect 349617 2527 349675 2533
rect 355410 2524 355416 2536
rect 355468 2524 355474 2576
rect 355502 2524 355508 2576
rect 355560 2524 355566 2576
rect 351914 2496 351920 2508
rect 347271 2400 347820 2428
rect 349724 2468 351920 2496
rect 347271 2397 347283 2400
rect 347225 2391 347283 2397
rect 349724 2360 349752 2468
rect 351914 2456 351920 2468
rect 351972 2456 351978 2508
rect 352926 2496 352932 2508
rect 352392 2468 352932 2496
rect 352392 2437 352420 2468
rect 352926 2456 352932 2468
rect 352984 2456 352990 2508
rect 349801 2431 349859 2437
rect 349801 2397 349813 2431
rect 349847 2397 349859 2431
rect 349801 2391 349859 2397
rect 352377 2431 352435 2437
rect 352377 2397 352389 2431
rect 352423 2397 352435 2431
rect 352377 2391 352435 2397
rect 354953 2431 355011 2437
rect 354953 2397 354965 2431
rect 354999 2428 355011 2431
rect 355520 2428 355548 2524
rect 357406 2496 357434 2604
rect 360654 2592 360660 2644
rect 360712 2592 360718 2644
rect 365070 2592 365076 2644
rect 365128 2592 365134 2644
rect 365254 2592 365260 2644
rect 365312 2632 365318 2644
rect 365809 2635 365867 2641
rect 365809 2632 365821 2635
rect 365312 2604 365821 2632
rect 365312 2592 365318 2604
rect 365809 2601 365821 2604
rect 365855 2632 365867 2635
rect 369854 2632 369860 2644
rect 365855 2604 369860 2632
rect 365855 2601 365867 2604
rect 365809 2595 365867 2601
rect 369854 2592 369860 2604
rect 369912 2592 369918 2644
rect 370225 2635 370283 2641
rect 370225 2601 370237 2635
rect 370271 2632 370283 2635
rect 373534 2632 373540 2644
rect 370271 2604 373540 2632
rect 370271 2601 370283 2604
rect 370225 2595 370283 2601
rect 373534 2592 373540 2604
rect 373592 2592 373598 2644
rect 376110 2592 376116 2644
rect 376168 2632 376174 2644
rect 378042 2632 378048 2644
rect 376168 2604 378048 2632
rect 376168 2592 376174 2604
rect 378042 2592 378048 2604
rect 378100 2592 378106 2644
rect 378134 2592 378140 2644
rect 378192 2632 378198 2644
rect 378689 2635 378747 2641
rect 378689 2632 378701 2635
rect 378192 2604 378701 2632
rect 378192 2592 378198 2604
rect 378689 2601 378701 2604
rect 378735 2632 378747 2635
rect 383194 2632 383200 2644
rect 378735 2604 383200 2632
rect 378735 2601 378747 2604
rect 378689 2595 378747 2601
rect 383194 2592 383200 2604
rect 383252 2592 383258 2644
rect 383286 2592 383292 2644
rect 383344 2632 383350 2644
rect 383838 2632 383844 2644
rect 383344 2604 383844 2632
rect 383344 2592 383350 2604
rect 383838 2592 383844 2604
rect 383896 2592 383902 2644
rect 385681 2635 385739 2641
rect 385681 2601 385693 2635
rect 385727 2632 385739 2635
rect 390646 2632 390652 2644
rect 385727 2604 390652 2632
rect 385727 2601 385739 2604
rect 385681 2595 385739 2601
rect 390646 2592 390652 2604
rect 390704 2592 390710 2644
rect 390833 2635 390891 2641
rect 390833 2601 390845 2635
rect 390879 2632 390891 2635
rect 394050 2632 394056 2644
rect 390879 2604 394056 2632
rect 390879 2601 390891 2604
rect 390833 2595 390891 2601
rect 394050 2592 394056 2604
rect 394108 2592 394114 2644
rect 398742 2592 398748 2644
rect 398800 2632 398806 2644
rect 399297 2635 399355 2641
rect 399297 2632 399309 2635
rect 398800 2604 399309 2632
rect 398800 2592 398806 2604
rect 399297 2601 399309 2604
rect 399343 2632 399355 2635
rect 408494 2632 408500 2644
rect 399343 2604 408500 2632
rect 399343 2601 399355 2604
rect 399297 2595 399355 2601
rect 408494 2592 408500 2604
rect 408552 2592 408558 2644
rect 412177 2635 412235 2641
rect 412177 2601 412189 2635
rect 412223 2632 412235 2635
rect 446582 2632 446588 2644
rect 412223 2604 446588 2632
rect 412223 2601 412235 2604
rect 412177 2595 412235 2601
rect 367649 2567 367707 2573
rect 367649 2533 367661 2567
rect 367695 2564 367707 2567
rect 373442 2564 373448 2576
rect 367695 2536 373448 2564
rect 367695 2533 367707 2536
rect 367649 2527 367707 2533
rect 373442 2524 373448 2536
rect 373500 2524 373506 2576
rect 375377 2567 375435 2573
rect 375377 2533 375389 2567
rect 375423 2564 375435 2567
rect 380894 2564 380900 2576
rect 375423 2536 380900 2564
rect 375423 2533 375435 2536
rect 375377 2527 375435 2533
rect 380894 2524 380900 2536
rect 380952 2524 380958 2576
rect 381078 2524 381084 2576
rect 381136 2564 381142 2576
rect 385034 2564 385040 2576
rect 381136 2536 385040 2564
rect 381136 2524 381142 2536
rect 385034 2524 385040 2536
rect 385092 2524 385098 2576
rect 388257 2567 388315 2573
rect 388257 2533 388269 2567
rect 388303 2564 388315 2567
rect 391934 2564 391940 2576
rect 388303 2536 391940 2564
rect 388303 2533 388315 2536
rect 388257 2527 388315 2533
rect 391934 2524 391940 2536
rect 391992 2524 391998 2576
rect 392026 2524 392032 2576
rect 392084 2564 392090 2576
rect 393314 2564 393320 2576
rect 392084 2536 393320 2564
rect 392084 2524 392090 2536
rect 393314 2524 393320 2536
rect 393372 2524 393378 2576
rect 393409 2567 393467 2573
rect 393409 2533 393421 2567
rect 393455 2564 393467 2567
rect 395246 2564 395252 2576
rect 393455 2536 395252 2564
rect 393455 2533 393467 2536
rect 393409 2527 393467 2533
rect 395246 2524 395252 2536
rect 395304 2524 395310 2576
rect 395985 2567 396043 2573
rect 395985 2533 395997 2567
rect 396031 2564 396043 2567
rect 397638 2564 397644 2576
rect 396031 2536 397644 2564
rect 396031 2533 396043 2536
rect 395985 2527 396043 2533
rect 397638 2524 397644 2536
rect 397696 2524 397702 2576
rect 398561 2567 398619 2573
rect 398561 2533 398573 2567
rect 398607 2564 398619 2567
rect 400214 2564 400220 2576
rect 398607 2536 400220 2564
rect 398607 2533 398619 2536
rect 398561 2527 398619 2533
rect 400214 2524 400220 2536
rect 400272 2524 400278 2576
rect 404354 2524 404360 2576
rect 404412 2524 404418 2576
rect 369946 2496 369952 2508
rect 357406 2468 369952 2496
rect 369946 2456 369952 2468
rect 370004 2456 370010 2508
rect 373537 2499 373595 2505
rect 373537 2465 373549 2499
rect 373583 2496 373595 2499
rect 400306 2496 400312 2508
rect 373583 2468 398144 2496
rect 373583 2465 373595 2468
rect 373537 2459 373595 2465
rect 354999 2400 355548 2428
rect 357529 2431 357587 2437
rect 354999 2397 355011 2400
rect 354953 2391 355011 2397
rect 357529 2397 357541 2431
rect 357575 2428 357587 2431
rect 360105 2431 360163 2437
rect 357575 2400 358124 2428
rect 357575 2397 357587 2400
rect 357529 2391 357587 2397
rect 325666 2332 349752 2360
rect 349816 2360 349844 2391
rect 350350 2360 350356 2372
rect 349816 2332 350356 2360
rect 350350 2320 350356 2332
rect 350408 2320 350414 2372
rect 357986 2360 357992 2372
rect 354784 2332 357992 2360
rect 323857 2295 323915 2301
rect 323857 2261 323869 2295
rect 323903 2261 323915 2295
rect 323857 2255 323915 2261
rect 324590 2252 324596 2304
rect 324648 2252 324654 2304
rect 326430 2252 326436 2304
rect 326488 2252 326494 2304
rect 329006 2252 329012 2304
rect 329064 2252 329070 2304
rect 329742 2252 329748 2304
rect 329800 2252 329806 2304
rect 331214 2252 331220 2304
rect 331272 2292 331278 2304
rect 331585 2295 331643 2301
rect 331585 2292 331597 2295
rect 331272 2264 331597 2292
rect 331272 2252 331278 2264
rect 331585 2261 331597 2264
rect 331631 2261 331643 2295
rect 331585 2255 331643 2261
rect 332318 2252 332324 2304
rect 332376 2252 332382 2304
rect 334158 2252 334164 2304
rect 334216 2252 334222 2304
rect 336734 2252 336740 2304
rect 336792 2252 336798 2304
rect 337470 2252 337476 2304
rect 337528 2252 337534 2304
rect 339310 2252 339316 2304
rect 339368 2252 339374 2304
rect 340046 2252 340052 2304
rect 340104 2252 340110 2304
rect 341886 2252 341892 2304
rect 341944 2252 341950 2304
rect 342622 2252 342628 2304
rect 342680 2252 342686 2304
rect 344462 2252 344468 2304
rect 344520 2252 344526 2304
rect 345198 2252 345204 2304
rect 345256 2252 345262 2304
rect 347038 2252 347044 2304
rect 347096 2252 347102 2304
rect 352190 2252 352196 2304
rect 352248 2252 352254 2304
rect 354784 2301 354812 2332
rect 357986 2320 357992 2332
rect 358044 2320 358050 2372
rect 358096 2304 358124 2400
rect 360105 2397 360117 2431
rect 360151 2428 360163 2431
rect 360654 2428 360660 2440
rect 360151 2400 360660 2428
rect 360151 2397 360163 2400
rect 360105 2391 360163 2397
rect 360654 2388 360660 2400
rect 360712 2388 360718 2440
rect 362681 2431 362739 2437
rect 362681 2397 362693 2431
rect 362727 2428 362739 2431
rect 362727 2400 363276 2428
rect 362727 2397 362739 2400
rect 362681 2391 362739 2397
rect 363248 2369 363276 2400
rect 365254 2388 365260 2440
rect 365312 2388 365318 2440
rect 367833 2431 367891 2437
rect 367833 2397 367845 2431
rect 367879 2428 367891 2431
rect 368382 2428 368388 2440
rect 367879 2400 368388 2428
rect 367879 2397 367891 2400
rect 367833 2391 367891 2397
rect 368382 2388 368388 2400
rect 368440 2388 368446 2440
rect 370409 2431 370467 2437
rect 370409 2397 370421 2431
rect 370455 2428 370467 2431
rect 370958 2428 370964 2440
rect 370455 2400 370964 2428
rect 370455 2397 370467 2400
rect 370409 2391 370467 2397
rect 370958 2388 370964 2400
rect 371016 2388 371022 2440
rect 372985 2431 373043 2437
rect 372985 2397 372997 2431
rect 373031 2428 373043 2431
rect 373552 2428 373580 2459
rect 373031 2400 373580 2428
rect 375561 2431 375619 2437
rect 373031 2397 373043 2400
rect 372985 2391 373043 2397
rect 375561 2397 375573 2431
rect 375607 2428 375619 2431
rect 376110 2428 376116 2440
rect 375607 2400 376116 2428
rect 375607 2397 375619 2400
rect 375561 2391 375619 2397
rect 376110 2388 376116 2400
rect 376168 2388 376174 2440
rect 378134 2388 378140 2440
rect 378192 2388 378198 2440
rect 380713 2431 380771 2437
rect 380713 2397 380725 2431
rect 380759 2428 380771 2431
rect 381262 2428 381268 2440
rect 380759 2400 381268 2428
rect 380759 2397 380771 2400
rect 380713 2391 380771 2397
rect 381262 2388 381268 2400
rect 381320 2388 381326 2440
rect 383289 2431 383347 2437
rect 383289 2397 383301 2431
rect 383335 2428 383347 2431
rect 383930 2428 383936 2440
rect 383335 2400 383936 2428
rect 383335 2397 383347 2400
rect 383289 2391 383347 2397
rect 383930 2388 383936 2400
rect 383988 2388 383994 2440
rect 385865 2431 385923 2437
rect 385865 2397 385877 2431
rect 385911 2428 385923 2431
rect 386414 2428 386420 2440
rect 385911 2400 386420 2428
rect 385911 2397 385923 2400
rect 385865 2391 385923 2397
rect 386414 2388 386420 2400
rect 386472 2388 386478 2440
rect 388441 2431 388499 2437
rect 388441 2397 388453 2431
rect 388487 2428 388499 2431
rect 388990 2428 388996 2440
rect 388487 2400 388996 2428
rect 388487 2397 388499 2400
rect 388441 2391 388499 2397
rect 388990 2388 388996 2400
rect 389048 2388 389054 2440
rect 391017 2431 391075 2437
rect 391017 2397 391029 2431
rect 391063 2428 391075 2431
rect 391566 2428 391572 2440
rect 391063 2400 391572 2428
rect 391063 2397 391075 2400
rect 391017 2391 391075 2397
rect 391566 2388 391572 2400
rect 391624 2388 391630 2440
rect 393314 2388 393320 2440
rect 393372 2428 393378 2440
rect 393593 2431 393651 2437
rect 393372 2400 393544 2428
rect 393372 2388 393378 2400
rect 363233 2363 363291 2369
rect 363233 2329 363245 2363
rect 363279 2360 363291 2363
rect 393516 2360 393544 2400
rect 393593 2397 393605 2431
rect 393639 2428 393651 2431
rect 394142 2428 394148 2440
rect 393639 2400 394148 2428
rect 393639 2397 393651 2400
rect 393593 2391 393651 2397
rect 394142 2388 394148 2400
rect 394200 2388 394206 2440
rect 396169 2431 396227 2437
rect 396169 2397 396181 2431
rect 396215 2428 396227 2431
rect 396718 2428 396724 2440
rect 396215 2400 396724 2428
rect 396215 2397 396227 2400
rect 396169 2391 396227 2397
rect 396718 2388 396724 2400
rect 396776 2388 396782 2440
rect 398116 2428 398144 2468
rect 398576 2468 400312 2496
rect 398576 2428 398604 2468
rect 400306 2456 400312 2468
rect 400364 2456 400370 2508
rect 401873 2499 401931 2505
rect 401873 2496 401885 2499
rect 401336 2468 401885 2496
rect 398116 2400 398604 2428
rect 398742 2388 398748 2440
rect 398800 2388 398806 2440
rect 401336 2437 401364 2468
rect 401873 2465 401885 2468
rect 401919 2496 401931 2499
rect 401919 2468 409736 2496
rect 401919 2465 401931 2468
rect 401873 2459 401931 2465
rect 401321 2431 401379 2437
rect 401321 2397 401333 2431
rect 401367 2397 401379 2431
rect 401321 2391 401379 2397
rect 403897 2431 403955 2437
rect 403897 2397 403909 2431
rect 403943 2428 403955 2431
rect 404354 2428 404360 2440
rect 403943 2400 404360 2428
rect 403943 2397 403955 2400
rect 403897 2391 403955 2397
rect 404354 2388 404360 2400
rect 404412 2388 404418 2440
rect 406473 2431 406531 2437
rect 406473 2397 406485 2431
rect 406519 2428 406531 2431
rect 409049 2431 409107 2437
rect 406519 2400 407068 2428
rect 406519 2397 406531 2400
rect 406473 2391 406531 2397
rect 403986 2360 403992 2372
rect 363279 2332 393314 2360
rect 393516 2332 403992 2360
rect 363279 2329 363291 2332
rect 363233 2323 363291 2329
rect 354769 2295 354827 2301
rect 354769 2261 354781 2295
rect 354815 2261 354827 2295
rect 354769 2255 354827 2261
rect 357342 2252 357348 2304
rect 357400 2252 357406 2304
rect 358078 2252 358084 2304
rect 358136 2252 358142 2304
rect 359918 2252 359924 2304
rect 359976 2252 359982 2304
rect 362497 2295 362555 2301
rect 362497 2261 362509 2295
rect 362543 2292 362555 2295
rect 367094 2292 367100 2304
rect 362543 2264 367100 2292
rect 362543 2261 362555 2264
rect 362497 2255 362555 2261
rect 367094 2252 367100 2264
rect 367152 2252 367158 2304
rect 368382 2252 368388 2304
rect 368440 2252 368446 2304
rect 370958 2252 370964 2304
rect 371016 2252 371022 2304
rect 372801 2295 372859 2301
rect 372801 2261 372813 2295
rect 372847 2292 372859 2295
rect 376386 2292 376392 2304
rect 372847 2264 376392 2292
rect 372847 2261 372859 2264
rect 372801 2255 372859 2261
rect 376386 2252 376392 2264
rect 376444 2252 376450 2304
rect 377950 2252 377956 2304
rect 378008 2252 378014 2304
rect 380529 2295 380587 2301
rect 380529 2261 380541 2295
rect 380575 2292 380587 2295
rect 381078 2292 381084 2304
rect 380575 2264 381084 2292
rect 380575 2261 380587 2264
rect 380529 2255 380587 2261
rect 381078 2252 381084 2264
rect 381136 2252 381142 2304
rect 381262 2252 381268 2304
rect 381320 2252 381326 2304
rect 383102 2252 383108 2304
rect 383160 2252 383166 2304
rect 383194 2252 383200 2304
rect 383252 2292 383258 2304
rect 383746 2292 383752 2304
rect 383252 2264 383752 2292
rect 383252 2252 383258 2264
rect 383746 2252 383752 2264
rect 383804 2252 383810 2304
rect 383841 2295 383899 2301
rect 383841 2261 383853 2295
rect 383887 2292 383899 2295
rect 383930 2292 383936 2304
rect 383887 2264 383936 2292
rect 383887 2261 383899 2264
rect 383841 2255 383899 2261
rect 383930 2252 383936 2264
rect 383988 2252 383994 2304
rect 386414 2252 386420 2304
rect 386472 2252 386478 2304
rect 388990 2252 388996 2304
rect 389048 2252 389054 2304
rect 391566 2252 391572 2304
rect 391624 2252 391630 2304
rect 393286 2292 393314 2332
rect 403986 2320 403992 2332
rect 404044 2320 404050 2372
rect 407040 2304 407068 2400
rect 409049 2397 409061 2431
rect 409095 2428 409107 2431
rect 409095 2400 409644 2428
rect 409095 2397 409107 2400
rect 409049 2391 409107 2397
rect 409616 2304 409644 2400
rect 409708 2360 409736 2468
rect 411625 2431 411683 2437
rect 411625 2397 411637 2431
rect 411671 2428 411683 2431
rect 412192 2428 412220 2595
rect 446582 2592 446588 2604
rect 446640 2592 446646 2644
rect 450814 2592 450820 2644
rect 450872 2592 450878 2644
rect 453393 2635 453451 2641
rect 453393 2632 453405 2635
rect 453316 2604 453405 2632
rect 414750 2524 414756 2576
rect 414808 2524 414814 2576
rect 419902 2524 419908 2576
rect 419960 2524 419966 2576
rect 425057 2567 425115 2573
rect 425057 2533 425069 2567
rect 425103 2564 425115 2567
rect 426158 2564 426164 2576
rect 425103 2536 426164 2564
rect 425103 2533 425115 2536
rect 425057 2527 425115 2533
rect 411671 2400 412220 2428
rect 414201 2431 414259 2437
rect 411671 2397 411683 2400
rect 411625 2391 411683 2397
rect 414201 2397 414213 2431
rect 414247 2428 414259 2431
rect 414768 2428 414796 2524
rect 414247 2400 414796 2428
rect 416777 2431 416835 2437
rect 414247 2397 414259 2400
rect 414201 2391 414259 2397
rect 416777 2397 416789 2431
rect 416823 2428 416835 2431
rect 417326 2428 417332 2440
rect 416823 2400 417332 2428
rect 416823 2397 416835 2400
rect 416777 2391 416835 2397
rect 417326 2388 417332 2400
rect 417384 2388 417390 2440
rect 419353 2431 419411 2437
rect 419353 2397 419365 2431
rect 419399 2428 419411 2431
rect 419920 2428 419948 2524
rect 419399 2400 419948 2428
rect 421929 2431 421987 2437
rect 419399 2397 419411 2400
rect 419353 2391 419411 2397
rect 421929 2397 421941 2431
rect 421975 2428 421987 2431
rect 422478 2428 422484 2440
rect 421975 2400 422484 2428
rect 421975 2397 421987 2400
rect 421929 2391 421987 2397
rect 422478 2388 422484 2400
rect 422536 2388 422542 2440
rect 424505 2431 424563 2437
rect 424505 2397 424517 2431
rect 424551 2428 424563 2431
rect 425072 2428 425100 2527
rect 426158 2524 426164 2536
rect 426216 2524 426222 2576
rect 430206 2524 430212 2576
rect 430264 2524 430270 2576
rect 431770 2524 431776 2576
rect 431828 2564 431834 2576
rect 434625 2567 434683 2573
rect 434625 2564 434637 2567
rect 431828 2536 434637 2564
rect 431828 2524 431834 2536
rect 434625 2533 434637 2536
rect 434671 2533 434683 2567
rect 434625 2527 434683 2533
rect 435358 2524 435364 2576
rect 435416 2524 435422 2576
rect 436830 2524 436836 2576
rect 436888 2564 436894 2576
rect 439777 2567 439835 2573
rect 439777 2564 439789 2567
rect 436888 2536 439789 2564
rect 436888 2524 436894 2536
rect 439777 2533 439789 2536
rect 439823 2533 439835 2567
rect 439777 2527 439835 2533
rect 441586 2536 451274 2564
rect 424551 2400 425100 2428
rect 427081 2431 427139 2437
rect 424551 2397 424563 2400
rect 424505 2391 424563 2397
rect 427081 2397 427093 2431
rect 427127 2428 427139 2431
rect 427630 2428 427636 2440
rect 427127 2400 427636 2428
rect 427127 2397 427139 2400
rect 427081 2391 427139 2397
rect 427630 2388 427636 2400
rect 427688 2388 427694 2440
rect 429657 2431 429715 2437
rect 429657 2397 429669 2431
rect 429703 2428 429715 2431
rect 430224 2428 430252 2524
rect 429703 2400 430252 2428
rect 432233 2431 432291 2437
rect 429703 2397 429715 2400
rect 429657 2391 429715 2397
rect 432233 2397 432245 2431
rect 432279 2428 432291 2431
rect 432782 2428 432788 2440
rect 432279 2400 432788 2428
rect 432279 2397 432291 2400
rect 432233 2391 432291 2397
rect 432782 2388 432788 2400
rect 432840 2388 432846 2440
rect 434809 2431 434867 2437
rect 434809 2397 434821 2431
rect 434855 2428 434867 2431
rect 435376 2428 435404 2524
rect 437937 2499 437995 2505
rect 437937 2465 437949 2499
rect 437983 2496 437995 2499
rect 441586 2496 441614 2536
rect 437983 2468 441614 2496
rect 437983 2465 437995 2468
rect 437937 2459 437995 2465
rect 434855 2400 435404 2428
rect 437385 2431 437443 2437
rect 434855 2397 434867 2400
rect 434809 2391 434867 2397
rect 437385 2397 437397 2431
rect 437431 2428 437443 2431
rect 437952 2428 437980 2459
rect 445662 2456 445668 2508
rect 445720 2456 445726 2508
rect 437431 2400 437980 2428
rect 439961 2431 440019 2437
rect 437431 2397 437443 2400
rect 437385 2391 437443 2397
rect 439961 2397 439973 2431
rect 440007 2428 440019 2431
rect 442537 2431 442595 2437
rect 440007 2400 440556 2428
rect 440007 2397 440019 2400
rect 439961 2391 440019 2397
rect 440234 2360 440240 2372
rect 409708 2332 440240 2360
rect 440234 2320 440240 2332
rect 440292 2320 440298 2372
rect 440528 2304 440556 2400
rect 442537 2397 442549 2431
rect 442583 2428 442595 2431
rect 445113 2431 445171 2437
rect 442583 2400 443132 2428
rect 442583 2397 442595 2400
rect 442537 2391 442595 2397
rect 443104 2304 443132 2400
rect 445113 2397 445125 2431
rect 445159 2428 445171 2431
rect 445680 2428 445708 2456
rect 445159 2400 445708 2428
rect 447689 2431 447747 2437
rect 445159 2397 445171 2400
rect 445113 2391 445171 2397
rect 447689 2397 447701 2431
rect 447735 2428 447747 2431
rect 450265 2431 450323 2437
rect 447735 2400 448284 2428
rect 447735 2397 447747 2400
rect 447689 2391 447747 2397
rect 448256 2304 448284 2400
rect 450265 2397 450277 2431
rect 450311 2428 450323 2431
rect 450814 2428 450820 2440
rect 450311 2400 450820 2428
rect 450311 2397 450323 2400
rect 450265 2391 450323 2397
rect 450814 2388 450820 2400
rect 450872 2388 450878 2440
rect 451246 2360 451274 2536
rect 452841 2431 452899 2437
rect 452841 2397 452853 2431
rect 452887 2428 452899 2431
rect 453316 2428 453344 2604
rect 453393 2601 453405 2604
rect 453439 2632 453451 2635
rect 464522 2632 464528 2644
rect 453439 2604 464528 2632
rect 453439 2601 453451 2604
rect 453393 2595 453451 2601
rect 464522 2592 464528 2604
rect 464580 2592 464586 2644
rect 466273 2635 466331 2641
rect 466273 2601 466285 2635
rect 466319 2632 466331 2635
rect 483566 2632 483572 2644
rect 466319 2604 483572 2632
rect 466319 2601 466331 2604
rect 466273 2595 466331 2601
rect 455414 2524 455420 2576
rect 455472 2564 455478 2576
rect 457809 2567 457867 2573
rect 457809 2564 457821 2567
rect 455472 2536 457821 2564
rect 455472 2524 455478 2536
rect 457809 2533 457821 2536
rect 457855 2533 457867 2567
rect 457809 2527 457867 2533
rect 461121 2567 461179 2573
rect 461121 2533 461133 2567
rect 461167 2564 461179 2567
rect 466086 2564 466092 2576
rect 461167 2536 466092 2564
rect 461167 2533 461179 2536
rect 461121 2527 461179 2533
rect 459554 2496 459560 2508
rect 452887 2400 453344 2428
rect 453500 2468 459560 2496
rect 452887 2397 452899 2400
rect 452841 2391 452899 2397
rect 453500 2360 453528 2468
rect 459554 2456 459560 2468
rect 459612 2456 459618 2508
rect 455417 2431 455475 2437
rect 455417 2397 455429 2431
rect 455463 2428 455475 2431
rect 455966 2428 455972 2440
rect 455463 2400 455972 2428
rect 455463 2397 455475 2400
rect 455417 2391 455475 2397
rect 455966 2388 455972 2400
rect 456024 2388 456030 2440
rect 457993 2431 458051 2437
rect 457993 2397 458005 2431
rect 458039 2428 458051 2431
rect 460569 2431 460627 2437
rect 458039 2400 458588 2428
rect 458039 2397 458051 2400
rect 457993 2391 458051 2397
rect 458560 2369 458588 2400
rect 460569 2397 460581 2431
rect 460615 2428 460627 2431
rect 461136 2428 461164 2527
rect 466086 2524 466092 2536
rect 466144 2524 466150 2576
rect 460615 2400 461164 2428
rect 463145 2431 463203 2437
rect 460615 2397 460627 2400
rect 460569 2391 460627 2397
rect 463145 2397 463157 2431
rect 463191 2428 463203 2431
rect 463694 2428 463700 2440
rect 463191 2400 463700 2428
rect 463191 2397 463203 2400
rect 463145 2391 463203 2397
rect 463694 2388 463700 2400
rect 463752 2388 463758 2440
rect 465721 2431 465779 2437
rect 465721 2397 465733 2431
rect 465767 2428 465779 2431
rect 466288 2428 466316 2595
rect 483566 2592 483572 2604
rect 483624 2592 483630 2644
rect 484302 2592 484308 2644
rect 484360 2592 484366 2644
rect 466362 2524 466368 2576
rect 466420 2564 466426 2576
rect 483014 2564 483020 2576
rect 466420 2536 483020 2564
rect 466420 2524 466426 2536
rect 483014 2524 483020 2536
rect 483072 2524 483078 2576
rect 476577 2499 476635 2505
rect 476577 2465 476589 2499
rect 476623 2496 476635 2499
rect 481634 2496 481640 2508
rect 476623 2468 481640 2496
rect 476623 2465 476635 2468
rect 476577 2459 476635 2465
rect 465767 2400 466316 2428
rect 468297 2431 468355 2437
rect 465767 2397 465779 2400
rect 465721 2391 465779 2397
rect 468297 2397 468309 2431
rect 468343 2428 468355 2431
rect 468846 2428 468852 2440
rect 468343 2400 468852 2428
rect 468343 2397 468355 2400
rect 468297 2391 468355 2397
rect 468846 2388 468852 2400
rect 468904 2388 468910 2440
rect 470873 2431 470931 2437
rect 470873 2397 470885 2431
rect 470919 2428 470931 2431
rect 471422 2428 471428 2440
rect 470919 2400 471428 2428
rect 470919 2397 470931 2400
rect 470873 2391 470931 2397
rect 471422 2388 471428 2400
rect 471480 2388 471486 2440
rect 473449 2431 473507 2437
rect 473449 2397 473461 2431
rect 473495 2428 473507 2431
rect 473906 2428 473912 2440
rect 473495 2400 473912 2428
rect 473495 2397 473507 2400
rect 473449 2391 473507 2397
rect 473906 2388 473912 2400
rect 473964 2388 473970 2440
rect 476025 2431 476083 2437
rect 476025 2397 476037 2431
rect 476071 2428 476083 2431
rect 476592 2428 476620 2459
rect 481634 2456 481640 2468
rect 481692 2456 481698 2508
rect 481726 2456 481732 2508
rect 481784 2456 481790 2508
rect 488534 2456 488540 2508
rect 488592 2496 488598 2508
rect 488592 2468 488948 2496
rect 488592 2456 488598 2468
rect 476071 2400 476620 2428
rect 478601 2431 478659 2437
rect 476071 2397 476083 2400
rect 476025 2391 476083 2397
rect 478601 2397 478613 2431
rect 478647 2397 478659 2431
rect 478601 2391 478659 2397
rect 481177 2431 481235 2437
rect 481177 2397 481189 2431
rect 481223 2428 481235 2431
rect 481744 2428 481772 2456
rect 481223 2400 481772 2428
rect 483753 2431 483811 2437
rect 481223 2397 481235 2400
rect 481177 2391 481235 2397
rect 483753 2397 483765 2431
rect 483799 2428 483811 2431
rect 484302 2428 484308 2440
rect 483799 2400 484308 2428
rect 483799 2397 483811 2400
rect 483753 2391 483811 2397
rect 451246 2332 453528 2360
rect 458545 2363 458603 2369
rect 458545 2329 458557 2363
rect 458591 2360 458603 2363
rect 475378 2360 475384 2372
rect 458591 2332 475384 2360
rect 458591 2329 458603 2332
rect 458545 2323 458603 2329
rect 475378 2320 475384 2332
rect 475436 2320 475442 2372
rect 478616 2360 478644 2391
rect 484302 2388 484308 2400
rect 484360 2388 484366 2440
rect 485774 2388 485780 2440
rect 485832 2428 485838 2440
rect 486329 2431 486387 2437
rect 486329 2428 486341 2431
rect 485832 2400 486341 2428
rect 485832 2388 485838 2400
rect 486329 2397 486341 2400
rect 486375 2397 486387 2431
rect 486329 2391 486387 2397
rect 488718 2388 488724 2440
rect 488776 2388 488782 2440
rect 488920 2437 488948 2468
rect 488905 2431 488963 2437
rect 488905 2397 488917 2431
rect 488951 2397 488963 2431
rect 488905 2391 488963 2397
rect 491018 2388 491024 2440
rect 491076 2428 491082 2440
rect 491481 2431 491539 2437
rect 491481 2428 491493 2431
rect 491076 2400 491493 2428
rect 491076 2388 491082 2400
rect 491481 2397 491493 2400
rect 491527 2397 491539 2431
rect 491481 2391 491539 2397
rect 493594 2388 493600 2440
rect 493652 2428 493658 2440
rect 494057 2431 494115 2437
rect 494057 2428 494069 2431
rect 493652 2400 494069 2428
rect 493652 2388 493658 2400
rect 494057 2397 494069 2400
rect 494103 2397 494115 2431
rect 494057 2391 494115 2397
rect 496170 2388 496176 2440
rect 496228 2428 496234 2440
rect 496633 2431 496691 2437
rect 496633 2428 496645 2431
rect 496228 2400 496645 2428
rect 496228 2388 496234 2400
rect 496633 2397 496645 2400
rect 496679 2397 496691 2431
rect 496633 2391 496691 2397
rect 498746 2388 498752 2440
rect 498804 2428 498810 2440
rect 499209 2431 499267 2437
rect 499209 2428 499221 2431
rect 498804 2400 499221 2428
rect 498804 2388 498810 2400
rect 499209 2397 499221 2400
rect 499255 2397 499267 2431
rect 499209 2391 499267 2397
rect 501322 2388 501328 2440
rect 501380 2428 501386 2440
rect 501785 2431 501843 2437
rect 501785 2428 501797 2431
rect 501380 2400 501797 2428
rect 501380 2388 501386 2400
rect 501785 2397 501797 2400
rect 501831 2397 501843 2431
rect 501785 2391 501843 2397
rect 503898 2388 503904 2440
rect 503956 2428 503962 2440
rect 504361 2431 504419 2437
rect 504361 2428 504373 2431
rect 503956 2400 504373 2428
rect 503956 2388 503962 2400
rect 504361 2397 504373 2400
rect 504407 2397 504419 2431
rect 504361 2391 504419 2397
rect 506474 2388 506480 2440
rect 506532 2428 506538 2440
rect 506937 2431 506995 2437
rect 506937 2428 506949 2431
rect 506532 2400 506949 2428
rect 506532 2388 506538 2400
rect 506937 2397 506949 2400
rect 506983 2397 506995 2431
rect 506937 2391 506995 2397
rect 509050 2388 509056 2440
rect 509108 2428 509114 2440
rect 509513 2431 509571 2437
rect 509513 2428 509525 2431
rect 509108 2400 509525 2428
rect 509108 2388 509114 2400
rect 509513 2397 509525 2400
rect 509559 2397 509571 2431
rect 509513 2391 509571 2397
rect 511626 2388 511632 2440
rect 511684 2428 511690 2440
rect 512089 2431 512147 2437
rect 512089 2428 512101 2431
rect 511684 2400 512101 2428
rect 511684 2388 511690 2400
rect 512089 2397 512101 2400
rect 512135 2397 512147 2431
rect 512089 2391 512147 2397
rect 514202 2388 514208 2440
rect 514260 2428 514266 2440
rect 514665 2431 514723 2437
rect 514665 2428 514677 2431
rect 514260 2400 514677 2428
rect 514260 2388 514266 2400
rect 514665 2397 514677 2400
rect 514711 2397 514723 2431
rect 514665 2391 514723 2397
rect 479153 2363 479211 2369
rect 479153 2360 479165 2363
rect 478616 2332 479165 2360
rect 479153 2329 479165 2332
rect 479199 2360 479211 2363
rect 484946 2360 484952 2372
rect 479199 2332 484952 2360
rect 479199 2329 479211 2332
rect 479153 2323 479211 2329
rect 484946 2320 484952 2332
rect 485004 2320 485010 2372
rect 488736 2360 488764 2388
rect 488736 2332 514524 2360
rect 398834 2292 398840 2304
rect 393286 2264 398840 2292
rect 398834 2252 398840 2264
rect 398892 2252 398898 2304
rect 401137 2295 401195 2301
rect 401137 2261 401149 2295
rect 401183 2292 401195 2295
rect 402422 2292 402428 2304
rect 401183 2264 402428 2292
rect 401183 2261 401195 2264
rect 401137 2255 401195 2261
rect 402422 2252 402428 2264
rect 402480 2252 402486 2304
rect 403713 2295 403771 2301
rect 403713 2261 403725 2295
rect 403759 2292 403771 2295
rect 405918 2292 405924 2304
rect 403759 2264 405924 2292
rect 403759 2261 403771 2264
rect 403713 2255 403771 2261
rect 405918 2252 405924 2264
rect 405976 2252 405982 2304
rect 406286 2252 406292 2304
rect 406344 2252 406350 2304
rect 407022 2252 407028 2304
rect 407080 2252 407086 2304
rect 408862 2252 408868 2304
rect 408920 2252 408926 2304
rect 409598 2252 409604 2304
rect 409656 2252 409662 2304
rect 411438 2252 411444 2304
rect 411496 2252 411502 2304
rect 414014 2252 414020 2304
rect 414072 2252 414078 2304
rect 416498 2252 416504 2304
rect 416556 2292 416562 2304
rect 416593 2295 416651 2301
rect 416593 2292 416605 2295
rect 416556 2264 416605 2292
rect 416556 2252 416562 2264
rect 416593 2261 416605 2264
rect 416639 2261 416651 2295
rect 416593 2255 416651 2261
rect 417326 2252 417332 2304
rect 417384 2252 417390 2304
rect 419166 2252 419172 2304
rect 419224 2252 419230 2304
rect 421742 2252 421748 2304
rect 421800 2252 421806 2304
rect 422478 2252 422484 2304
rect 422536 2252 422542 2304
rect 423582 2252 423588 2304
rect 423640 2292 423646 2304
rect 424321 2295 424379 2301
rect 424321 2292 424333 2295
rect 423640 2264 424333 2292
rect 423640 2252 423646 2264
rect 424321 2261 424333 2264
rect 424367 2261 424379 2295
rect 424321 2255 424379 2261
rect 426066 2252 426072 2304
rect 426124 2292 426130 2304
rect 426897 2295 426955 2301
rect 426897 2292 426909 2295
rect 426124 2264 426909 2292
rect 426124 2252 426130 2264
rect 426897 2261 426909 2264
rect 426943 2261 426955 2295
rect 426897 2255 426955 2261
rect 427630 2252 427636 2304
rect 427688 2252 427694 2304
rect 427722 2252 427728 2304
rect 427780 2292 427786 2304
rect 429473 2295 429531 2301
rect 429473 2292 429485 2295
rect 427780 2264 429485 2292
rect 427780 2252 427786 2264
rect 429473 2261 429485 2264
rect 429519 2261 429531 2295
rect 429473 2255 429531 2261
rect 430482 2252 430488 2304
rect 430540 2292 430546 2304
rect 432049 2295 432107 2301
rect 432049 2292 432061 2295
rect 430540 2264 432061 2292
rect 430540 2252 430546 2264
rect 432049 2261 432061 2264
rect 432095 2261 432107 2295
rect 432049 2255 432107 2261
rect 432782 2252 432788 2304
rect 432840 2252 432846 2304
rect 434622 2252 434628 2304
rect 434680 2292 434686 2304
rect 437201 2295 437259 2301
rect 437201 2292 437213 2295
rect 434680 2264 437213 2292
rect 434680 2252 434686 2264
rect 437201 2261 437213 2264
rect 437247 2261 437259 2295
rect 437201 2255 437259 2261
rect 440510 2252 440516 2304
rect 440568 2252 440574 2304
rect 442350 2252 442356 2304
rect 442408 2252 442414 2304
rect 443086 2252 443092 2304
rect 443144 2252 443150 2304
rect 444374 2252 444380 2304
rect 444432 2292 444438 2304
rect 444929 2295 444987 2301
rect 444929 2292 444941 2295
rect 444432 2264 444941 2292
rect 444432 2252 444438 2264
rect 444929 2261 444941 2264
rect 444975 2261 444987 2295
rect 444929 2255 444987 2261
rect 445754 2252 445760 2304
rect 445812 2292 445818 2304
rect 447505 2295 447563 2301
rect 447505 2292 447517 2295
rect 445812 2264 447517 2292
rect 445812 2252 445818 2264
rect 447505 2261 447517 2264
rect 447551 2261 447563 2295
rect 447505 2255 447563 2261
rect 448238 2252 448244 2304
rect 448296 2252 448302 2304
rect 448514 2252 448520 2304
rect 448572 2292 448578 2304
rect 450081 2295 450139 2301
rect 450081 2292 450093 2295
rect 448572 2264 450093 2292
rect 448572 2252 448578 2264
rect 450081 2261 450093 2264
rect 450127 2261 450139 2295
rect 450081 2255 450139 2261
rect 451366 2252 451372 2304
rect 451424 2292 451430 2304
rect 452657 2295 452715 2301
rect 452657 2292 452669 2295
rect 451424 2264 452669 2292
rect 451424 2252 451430 2264
rect 452657 2261 452669 2264
rect 452703 2261 452715 2295
rect 452657 2255 452715 2261
rect 453390 2252 453396 2304
rect 453448 2292 453454 2304
rect 455233 2295 455291 2301
rect 455233 2292 455245 2295
rect 453448 2264 455245 2292
rect 453448 2252 453454 2264
rect 455233 2261 455245 2264
rect 455279 2261 455291 2295
rect 455233 2255 455291 2261
rect 460382 2252 460388 2304
rect 460440 2252 460446 2304
rect 462314 2252 462320 2304
rect 462372 2292 462378 2304
rect 462961 2295 463019 2301
rect 462961 2292 462973 2295
rect 462372 2264 462973 2292
rect 462372 2252 462378 2264
rect 462961 2261 462973 2264
rect 463007 2261 463019 2295
rect 462961 2255 463019 2261
rect 463694 2252 463700 2304
rect 463752 2252 463758 2304
rect 463786 2252 463792 2304
rect 463844 2292 463850 2304
rect 465537 2295 465595 2301
rect 465537 2292 465549 2295
rect 463844 2264 465549 2292
rect 463844 2252 463850 2264
rect 465537 2261 465549 2264
rect 465583 2261 465595 2295
rect 465537 2255 465595 2261
rect 466454 2252 466460 2304
rect 466512 2292 466518 2304
rect 468113 2295 468171 2301
rect 468113 2292 468125 2295
rect 466512 2264 468125 2292
rect 466512 2252 466518 2264
rect 468113 2261 468125 2264
rect 468159 2261 468171 2295
rect 468113 2255 468171 2261
rect 468846 2252 468852 2304
rect 468904 2252 468910 2304
rect 469214 2252 469220 2304
rect 469272 2292 469278 2304
rect 470689 2295 470747 2301
rect 470689 2292 470701 2295
rect 469272 2264 470701 2292
rect 469272 2252 469278 2264
rect 470689 2261 470701 2264
rect 470735 2261 470747 2295
rect 470689 2255 470747 2261
rect 471422 2252 471428 2304
rect 471480 2252 471486 2304
rect 471882 2252 471888 2304
rect 471940 2292 471946 2304
rect 473265 2295 473323 2301
rect 473265 2292 473277 2295
rect 471940 2264 473277 2292
rect 471940 2252 471946 2264
rect 473265 2261 473277 2264
rect 473311 2261 473323 2295
rect 473265 2255 473323 2261
rect 473906 2252 473912 2304
rect 473964 2252 473970 2304
rect 473998 2252 474004 2304
rect 474056 2292 474062 2304
rect 475841 2295 475899 2301
rect 475841 2292 475853 2295
rect 474056 2264 475853 2292
rect 474056 2252 474062 2264
rect 475841 2261 475853 2264
rect 475887 2261 475899 2295
rect 475841 2255 475899 2261
rect 475930 2252 475936 2304
rect 475988 2292 475994 2304
rect 478417 2295 478475 2301
rect 478417 2292 478429 2295
rect 475988 2264 478429 2292
rect 475988 2252 475994 2264
rect 478417 2261 478429 2264
rect 478463 2261 478475 2295
rect 478417 2255 478475 2261
rect 478506 2252 478512 2304
rect 478564 2292 478570 2304
rect 480993 2295 481051 2301
rect 480993 2292 481005 2295
rect 478564 2264 481005 2292
rect 478564 2252 478570 2264
rect 480993 2261 481005 2264
rect 481039 2261 481051 2295
rect 480993 2255 481051 2261
rect 483566 2252 483572 2304
rect 483624 2252 483630 2304
rect 486142 2252 486148 2304
rect 486200 2252 486206 2304
rect 488718 2252 488724 2304
rect 488776 2252 488782 2304
rect 491294 2252 491300 2304
rect 491352 2252 491358 2304
rect 493870 2252 493876 2304
rect 493928 2252 493934 2304
rect 496446 2252 496452 2304
rect 496504 2252 496510 2304
rect 498194 2252 498200 2304
rect 498252 2292 498258 2304
rect 499025 2295 499083 2301
rect 499025 2292 499037 2295
rect 498252 2264 499037 2292
rect 498252 2252 498258 2264
rect 499025 2261 499037 2264
rect 499071 2261 499083 2295
rect 499025 2255 499083 2261
rect 500310 2252 500316 2304
rect 500368 2292 500374 2304
rect 501601 2295 501659 2301
rect 501601 2292 501613 2295
rect 500368 2264 501613 2292
rect 500368 2252 500374 2264
rect 501601 2261 501613 2264
rect 501647 2261 501659 2295
rect 501601 2255 501659 2261
rect 502334 2252 502340 2304
rect 502392 2292 502398 2304
rect 504177 2295 504235 2301
rect 504177 2292 504189 2295
rect 502392 2264 504189 2292
rect 502392 2252 502398 2264
rect 504177 2261 504189 2264
rect 504223 2261 504235 2295
rect 504177 2255 504235 2261
rect 505094 2252 505100 2304
rect 505152 2292 505158 2304
rect 506753 2295 506811 2301
rect 506753 2292 506765 2295
rect 505152 2264 506765 2292
rect 505152 2252 505158 2264
rect 506753 2261 506765 2264
rect 506799 2261 506811 2295
rect 506753 2255 506811 2261
rect 509326 2252 509332 2304
rect 509384 2252 509390 2304
rect 510522 2252 510528 2304
rect 510580 2292 510586 2304
rect 514496 2301 514524 2332
rect 511905 2295 511963 2301
rect 511905 2292 511917 2295
rect 510580 2264 511917 2292
rect 510580 2252 510586 2264
rect 511905 2261 511917 2264
rect 511951 2261 511963 2295
rect 511905 2255 511963 2261
rect 514481 2295 514539 2301
rect 514481 2261 514493 2295
rect 514527 2261 514539 2295
rect 514481 2255 514539 2261
rect 1104 2202 528816 2224
rect 1104 2150 67574 2202
rect 67626 2150 67638 2202
rect 67690 2150 67702 2202
rect 67754 2150 67766 2202
rect 67818 2150 67830 2202
rect 67882 2150 199502 2202
rect 199554 2150 199566 2202
rect 199618 2150 199630 2202
rect 199682 2150 199694 2202
rect 199746 2150 199758 2202
rect 199810 2150 331430 2202
rect 331482 2150 331494 2202
rect 331546 2150 331558 2202
rect 331610 2150 331622 2202
rect 331674 2150 331686 2202
rect 331738 2150 463358 2202
rect 463410 2150 463422 2202
rect 463474 2150 463486 2202
rect 463538 2150 463550 2202
rect 463602 2150 463614 2202
rect 463666 2150 528816 2202
rect 1104 2128 528816 2150
rect 37918 2048 37924 2100
rect 37976 2088 37982 2100
rect 98638 2088 98644 2100
rect 37976 2060 98644 2088
rect 37976 2048 37982 2060
rect 98638 2048 98644 2060
rect 98696 2048 98702 2100
rect 99742 2048 99748 2100
rect 99800 2088 99806 2100
rect 127710 2088 127716 2100
rect 99800 2060 127716 2088
rect 99800 2048 99806 2060
rect 127710 2048 127716 2060
rect 127768 2048 127774 2100
rect 127986 2048 127992 2100
rect 128044 2088 128050 2100
rect 136450 2088 136456 2100
rect 128044 2060 136456 2088
rect 128044 2048 128050 2060
rect 136450 2048 136456 2060
rect 136508 2048 136514 2100
rect 143442 2048 143448 2100
rect 143500 2088 143506 2100
rect 191098 2088 191104 2100
rect 143500 2060 191104 2088
rect 143500 2048 143506 2060
rect 191098 2048 191104 2060
rect 191156 2048 191162 2100
rect 195054 2048 195060 2100
rect 195112 2088 195118 2100
rect 263134 2088 263140 2100
rect 195112 2060 263140 2088
rect 195112 2048 195118 2060
rect 263134 2048 263140 2060
rect 263192 2048 263198 2100
rect 340046 2048 340052 2100
rect 340104 2088 340110 2100
rect 340104 2060 373948 2088
rect 340104 2048 340110 2060
rect 30190 1980 30196 2032
rect 30248 2020 30254 2032
rect 48774 2020 48780 2032
rect 30248 1992 48780 2020
rect 30248 1980 30254 1992
rect 48774 1980 48780 1992
rect 48832 1980 48838 2032
rect 53374 1980 53380 2032
rect 53432 2020 53438 2032
rect 108666 2020 108672 2032
rect 53432 1992 108672 2020
rect 53432 1980 53438 1992
rect 108666 1980 108672 1992
rect 108724 1980 108730 2032
rect 108758 1980 108764 2032
rect 108816 2020 108822 2032
rect 130654 2020 130660 2032
rect 108816 1992 130660 2020
rect 108816 1980 108822 1992
rect 130654 1980 130660 1992
rect 130712 1980 130718 2032
rect 139118 1980 139124 2032
rect 139176 2020 139182 2032
rect 143074 2020 143080 2032
rect 139176 1992 143080 2020
rect 139176 1980 139182 1992
rect 143074 1980 143080 1992
rect 143132 1980 143138 2032
rect 151998 1980 152004 2032
rect 152056 2020 152062 2032
rect 195606 2020 195612 2032
rect 152056 1992 195612 2020
rect 152056 1980 152062 1992
rect 195606 1980 195612 1992
rect 195664 1980 195670 2032
rect 200206 1980 200212 2032
rect 200264 2020 200270 2032
rect 264330 2020 264336 2032
rect 200264 1992 264336 2020
rect 200264 1980 200270 1992
rect 264330 1980 264336 1992
rect 264388 1980 264394 2032
rect 342622 1980 342628 2032
rect 342680 2020 342686 2032
rect 373920 2020 373948 2060
rect 377950 2048 377956 2100
rect 378008 2088 378014 2100
rect 383286 2088 383292 2100
rect 378008 2060 383292 2088
rect 378008 2048 378014 2060
rect 383286 2048 383292 2060
rect 383344 2048 383350 2100
rect 383930 2048 383936 2100
rect 383988 2088 383994 2100
rect 397362 2088 397368 2100
rect 383988 2060 397368 2088
rect 383988 2048 383994 2060
rect 397362 2048 397368 2060
rect 397420 2048 397426 2100
rect 409598 2048 409604 2100
rect 409656 2088 409662 2100
rect 443730 2088 443736 2100
rect 409656 2060 443736 2088
rect 409656 2048 409662 2060
rect 443730 2048 443736 2060
rect 443788 2048 443794 2100
rect 475378 2048 475384 2100
rect 475436 2088 475442 2100
rect 482738 2088 482744 2100
rect 475436 2060 482744 2088
rect 475436 2048 475442 2060
rect 482738 2048 482744 2060
rect 482796 2048 482802 2100
rect 342680 1992 373856 2020
rect 373920 1992 379514 2020
rect 342680 1980 342686 1992
rect 35342 1912 35348 1964
rect 35400 1952 35406 1964
rect 56502 1952 56508 1964
rect 35400 1924 56508 1952
rect 35400 1912 35406 1924
rect 56502 1912 56508 1924
rect 56560 1912 56566 1964
rect 58526 1912 58532 1964
rect 58584 1952 58590 1964
rect 115474 1952 115480 1964
rect 58584 1924 115480 1952
rect 58584 1912 58590 1924
rect 115474 1912 115480 1924
rect 115532 1912 115538 1964
rect 122926 1912 122932 1964
rect 122984 1952 122990 1964
rect 141694 1952 141700 1964
rect 122984 1924 141700 1952
rect 122984 1912 122990 1924
rect 141694 1912 141700 1924
rect 141752 1912 141758 1964
rect 157150 1912 157156 1964
rect 157208 1952 157214 1964
rect 196066 1952 196072 1964
rect 157208 1924 196072 1952
rect 157208 1912 157214 1924
rect 196066 1912 196072 1924
rect 196124 1912 196130 1964
rect 215662 1912 215668 1964
rect 215720 1952 215726 1964
rect 268378 1952 268384 1964
rect 215720 1924 268384 1952
rect 215720 1912 215726 1924
rect 268378 1912 268384 1924
rect 268436 1912 268442 1964
rect 302326 1912 302332 1964
rect 302384 1952 302390 1964
rect 321278 1952 321284 1964
rect 302384 1924 321284 1952
rect 302384 1912 302390 1924
rect 321278 1912 321284 1924
rect 321336 1912 321342 1964
rect 329742 1912 329748 1964
rect 329800 1952 329806 1964
rect 365622 1952 365628 1964
rect 329800 1924 365628 1952
rect 329800 1912 329806 1924
rect 365622 1912 365628 1924
rect 365680 1912 365686 1964
rect 66714 1844 66720 1896
rect 66772 1884 66778 1896
rect 70394 1884 70400 1896
rect 66772 1856 70400 1884
rect 66772 1844 66778 1856
rect 70394 1844 70400 1856
rect 70452 1844 70458 1896
rect 74902 1844 74908 1896
rect 74960 1884 74966 1896
rect 78674 1884 78680 1896
rect 74960 1856 78680 1884
rect 74960 1844 74966 1856
rect 78674 1844 78680 1856
rect 78732 1844 78738 1896
rect 80238 1844 80244 1896
rect 80296 1884 80302 1896
rect 89806 1884 89812 1896
rect 80296 1856 89812 1884
rect 80296 1844 80302 1856
rect 89806 1844 89812 1856
rect 89864 1844 89870 1896
rect 91830 1844 91836 1896
rect 91888 1884 91894 1896
rect 102134 1884 102140 1896
rect 91888 1856 102140 1884
rect 91888 1844 91894 1856
rect 102134 1844 102140 1856
rect 102192 1844 102198 1896
rect 102226 1844 102232 1896
rect 102284 1884 102290 1896
rect 107930 1884 107936 1896
rect 102284 1856 107936 1884
rect 102284 1844 102290 1856
rect 107930 1844 107936 1856
rect 107988 1844 107994 1896
rect 115290 1884 115296 1896
rect 109006 1856 115296 1884
rect 14734 1776 14740 1828
rect 14792 1816 14798 1828
rect 96798 1816 96804 1828
rect 14792 1788 96804 1816
rect 14792 1776 14798 1788
rect 96798 1776 96804 1788
rect 96856 1776 96862 1828
rect 97442 1776 97448 1828
rect 97500 1816 97506 1828
rect 109006 1816 109034 1856
rect 115290 1844 115296 1856
rect 115348 1844 115354 1896
rect 120350 1844 120356 1896
rect 120408 1884 120414 1896
rect 143166 1884 143172 1896
rect 120408 1856 143172 1884
rect 120408 1844 120414 1856
rect 143166 1844 143172 1856
rect 143224 1844 143230 1896
rect 148962 1844 148968 1896
rect 149020 1884 149026 1896
rect 157242 1884 157248 1896
rect 149020 1856 157248 1884
rect 149020 1844 149026 1856
rect 157242 1844 157248 1856
rect 157300 1844 157306 1896
rect 158990 1844 158996 1896
rect 159048 1884 159054 1896
rect 159048 1856 162072 1884
rect 159048 1844 159054 1856
rect 97500 1788 109034 1816
rect 97500 1776 97506 1788
rect 109218 1776 109224 1828
rect 109276 1816 109282 1828
rect 125502 1816 125508 1828
rect 109276 1788 125508 1816
rect 109276 1776 109282 1788
rect 125502 1776 125508 1788
rect 125560 1776 125566 1828
rect 130838 1776 130844 1828
rect 130896 1816 130902 1828
rect 148134 1816 148140 1828
rect 130896 1788 148140 1816
rect 130896 1776 130902 1788
rect 148134 1776 148140 1788
rect 148192 1776 148198 1828
rect 161934 1816 161940 1828
rect 148244 1788 161940 1816
rect 7006 1708 7012 1760
rect 7064 1748 7070 1760
rect 75546 1748 75552 1760
rect 7064 1720 75552 1748
rect 7064 1708 7070 1720
rect 75546 1708 75552 1720
rect 75604 1708 75610 1760
rect 75638 1708 75644 1760
rect 75696 1748 75702 1760
rect 80146 1748 80152 1760
rect 75696 1720 80152 1748
rect 75696 1708 75702 1720
rect 80146 1708 80152 1720
rect 80204 1708 80210 1760
rect 80330 1708 80336 1760
rect 80388 1748 80394 1760
rect 86954 1748 86960 1760
rect 80388 1720 86960 1748
rect 80388 1708 80394 1720
rect 86954 1708 86960 1720
rect 87012 1708 87018 1760
rect 87046 1708 87052 1760
rect 87104 1748 87110 1760
rect 92290 1748 92296 1760
rect 87104 1720 92296 1748
rect 87104 1708 87110 1720
rect 92290 1708 92296 1720
rect 92348 1708 92354 1760
rect 99558 1748 99564 1760
rect 94516 1720 99564 1748
rect 25038 1640 25044 1692
rect 25096 1680 25102 1692
rect 94516 1680 94544 1720
rect 99558 1708 99564 1720
rect 99616 1708 99622 1760
rect 103422 1748 103428 1760
rect 99760 1720 103428 1748
rect 25096 1652 94544 1680
rect 25096 1640 25102 1652
rect 94590 1640 94596 1692
rect 94648 1680 94654 1692
rect 99760 1680 99788 1720
rect 103422 1708 103428 1720
rect 103480 1708 103486 1760
rect 107470 1708 107476 1760
rect 107528 1748 107534 1760
rect 114922 1748 114928 1760
rect 107528 1720 114928 1748
rect 107528 1708 107534 1720
rect 114922 1708 114928 1720
rect 114980 1708 114986 1760
rect 118694 1708 118700 1760
rect 118752 1748 118758 1760
rect 127618 1748 127624 1760
rect 118752 1720 127624 1748
rect 118752 1708 118758 1720
rect 127618 1708 127624 1720
rect 127676 1708 127682 1760
rect 128170 1708 128176 1760
rect 128228 1748 128234 1760
rect 132586 1748 132592 1760
rect 128228 1720 132592 1748
rect 128228 1708 128234 1720
rect 132586 1708 132592 1720
rect 132644 1708 132650 1760
rect 141050 1748 141056 1760
rect 133156 1720 141056 1748
rect 111978 1680 111984 1692
rect 94648 1652 99788 1680
rect 101232 1652 111984 1680
rect 94648 1640 94654 1652
rect 50798 1572 50804 1624
rect 50856 1612 50862 1624
rect 101232 1612 101260 1652
rect 111978 1640 111984 1652
rect 112036 1640 112042 1692
rect 112806 1640 112812 1692
rect 112864 1680 112870 1692
rect 121454 1680 121460 1692
rect 112864 1652 121460 1680
rect 112864 1640 112870 1652
rect 121454 1640 121460 1652
rect 121512 1640 121518 1692
rect 121730 1640 121736 1692
rect 121788 1680 121794 1692
rect 132494 1680 132500 1692
rect 121788 1652 132500 1680
rect 121788 1640 121794 1652
rect 132494 1640 132500 1652
rect 132552 1640 132558 1692
rect 50856 1584 101260 1612
rect 50856 1572 50862 1584
rect 104894 1572 104900 1624
rect 104952 1612 104958 1624
rect 110782 1612 110788 1624
rect 104952 1584 110788 1612
rect 104952 1572 104958 1584
rect 110782 1572 110788 1584
rect 110840 1572 110846 1624
rect 115198 1572 115204 1624
rect 115256 1612 115262 1624
rect 133156 1612 133184 1720
rect 141050 1708 141056 1720
rect 141108 1708 141114 1760
rect 145834 1708 145840 1760
rect 145892 1748 145898 1760
rect 148244 1748 148272 1788
rect 161934 1776 161940 1788
rect 161992 1776 161998 1828
rect 162044 1816 162072 1856
rect 162302 1844 162308 1896
rect 162360 1884 162366 1896
rect 196710 1884 196716 1896
rect 162360 1856 196716 1884
rect 162360 1844 162366 1856
rect 196710 1844 196716 1856
rect 196768 1844 196774 1896
rect 220814 1844 220820 1896
rect 220872 1884 220878 1896
rect 269666 1884 269672 1896
rect 220872 1856 269672 1884
rect 220872 1844 220878 1856
rect 269666 1844 269672 1856
rect 269724 1844 269730 1896
rect 358078 1844 358084 1896
rect 358136 1884 358142 1896
rect 358136 1856 369854 1884
rect 358136 1844 358142 1856
rect 163682 1816 163688 1828
rect 162044 1788 163688 1816
rect 163682 1776 163688 1788
rect 163740 1776 163746 1828
rect 163958 1816 163964 1828
rect 163792 1788 163964 1816
rect 145892 1720 148272 1748
rect 145892 1708 145898 1720
rect 148502 1708 148508 1760
rect 148560 1748 148566 1760
rect 158530 1748 158536 1760
rect 148560 1720 158536 1748
rect 148560 1708 148566 1720
rect 158530 1708 158536 1720
rect 158588 1708 158594 1760
rect 161198 1708 161204 1760
rect 161256 1748 161262 1760
rect 163792 1748 163820 1788
rect 163958 1776 163964 1788
rect 164016 1776 164022 1828
rect 167454 1776 167460 1828
rect 167512 1816 167518 1828
rect 198734 1816 198740 1828
rect 167512 1788 198740 1816
rect 167512 1776 167518 1788
rect 198734 1776 198740 1788
rect 198792 1776 198798 1828
rect 225966 1776 225972 1828
rect 226024 1816 226030 1828
rect 270586 1816 270592 1828
rect 226024 1788 270592 1816
rect 226024 1776 226030 1788
rect 270586 1776 270592 1788
rect 270644 1776 270650 1828
rect 352190 1776 352196 1828
rect 352248 1816 352254 1828
rect 359826 1816 359832 1828
rect 352248 1788 359832 1816
rect 352248 1776 352254 1788
rect 359826 1776 359832 1788
rect 359884 1776 359890 1828
rect 369826 1816 369854 1856
rect 373828 1816 373856 1992
rect 379486 1952 379514 1992
rect 383102 1980 383108 2032
rect 383160 2020 383166 2032
rect 387794 2020 387800 2032
rect 383160 1992 387800 2020
rect 383160 1980 383166 1992
rect 387794 1980 387800 1992
rect 387852 1980 387858 2032
rect 391566 1980 391572 2032
rect 391624 2020 391630 2032
rect 420914 2020 420920 2032
rect 391624 1992 420920 2020
rect 391624 1980 391630 1992
rect 420914 1980 420920 1992
rect 420972 1980 420978 2032
rect 422478 1980 422484 2032
rect 422536 2020 422542 2032
rect 447686 2020 447692 2032
rect 422536 1992 447692 2020
rect 422536 1980 422542 1992
rect 447686 1980 447692 1992
rect 447744 1980 447750 2032
rect 463694 1980 463700 2032
rect 463752 2020 463758 2032
rect 481818 2020 481824 2032
rect 463752 1992 481824 2020
rect 463752 1980 463758 1992
rect 481818 1980 481824 1992
rect 481876 1980 481882 2032
rect 382274 1952 382280 1964
rect 379486 1924 382280 1952
rect 382274 1912 382280 1924
rect 382332 1912 382338 1964
rect 383746 1912 383752 1964
rect 383804 1952 383810 1964
rect 392026 1952 392032 1964
rect 383804 1924 392032 1952
rect 383804 1912 383810 1924
rect 392026 1912 392032 1924
rect 392084 1912 392090 1964
rect 417326 1912 417332 1964
rect 417384 1952 417390 1964
rect 447134 1952 447140 1964
rect 417384 1924 447140 1952
rect 417384 1912 417390 1924
rect 447134 1912 447140 1924
rect 447192 1912 447198 1964
rect 471422 1912 471428 1964
rect 471480 1952 471486 1964
rect 484118 1952 484124 1964
rect 471480 1924 484124 1952
rect 471480 1912 471486 1924
rect 484118 1912 484124 1924
rect 484176 1912 484182 1964
rect 443086 1844 443092 1896
rect 443144 1884 443150 1896
rect 481174 1884 481180 1896
rect 443144 1856 481180 1884
rect 443144 1844 443150 1856
rect 481174 1844 481180 1856
rect 481232 1844 481238 1896
rect 378686 1816 378692 1828
rect 369826 1788 372936 1816
rect 373828 1788 378692 1816
rect 172514 1748 172520 1760
rect 161256 1720 163820 1748
rect 163884 1720 172520 1748
rect 161256 1708 161262 1720
rect 133966 1640 133972 1692
rect 134024 1680 134030 1692
rect 163884 1680 163912 1720
rect 172514 1708 172520 1720
rect 172572 1708 172578 1760
rect 172606 1708 172612 1760
rect 172664 1748 172670 1760
rect 186866 1748 186872 1760
rect 172664 1720 186872 1748
rect 172664 1708 172670 1720
rect 186866 1708 186872 1720
rect 186924 1708 186930 1760
rect 188338 1708 188344 1760
rect 188396 1748 188402 1760
rect 192938 1748 192944 1760
rect 188396 1720 192944 1748
rect 188396 1708 188402 1720
rect 192938 1708 192944 1720
rect 192996 1708 193002 1760
rect 195974 1748 195980 1760
rect 193186 1720 195980 1748
rect 134024 1652 163912 1680
rect 134024 1640 134030 1652
rect 163958 1640 163964 1692
rect 164016 1680 164022 1692
rect 168098 1680 168104 1692
rect 164016 1652 168104 1680
rect 164016 1640 164022 1652
rect 168098 1640 168104 1652
rect 168156 1640 168162 1692
rect 168282 1640 168288 1692
rect 168340 1680 168346 1692
rect 185486 1680 185492 1692
rect 168340 1652 185492 1680
rect 168340 1640 168346 1652
rect 185486 1640 185492 1652
rect 185544 1640 185550 1692
rect 185854 1640 185860 1692
rect 185912 1680 185918 1692
rect 193186 1680 193214 1720
rect 195974 1708 195980 1720
rect 196032 1708 196038 1760
rect 337470 1708 337476 1760
rect 337528 1748 337534 1760
rect 372798 1748 372804 1760
rect 337528 1720 372804 1748
rect 337528 1708 337534 1720
rect 372798 1708 372804 1720
rect 372856 1708 372862 1760
rect 372908 1748 372936 1788
rect 378686 1776 378692 1788
rect 378744 1776 378750 1828
rect 388990 1776 388996 1828
rect 389048 1816 389054 1828
rect 432046 1816 432052 1828
rect 389048 1788 432052 1816
rect 389048 1776 389054 1788
rect 432046 1776 432052 1788
rect 432104 1776 432110 1828
rect 468846 1776 468852 1828
rect 468904 1816 468910 1828
rect 480254 1816 480260 1828
rect 468904 1788 480260 1816
rect 468904 1776 468910 1788
rect 480254 1776 480260 1788
rect 480312 1776 480318 1828
rect 381538 1748 381544 1760
rect 372908 1720 381544 1748
rect 381538 1708 381544 1720
rect 381596 1708 381602 1760
rect 394142 1708 394148 1760
rect 394200 1748 394206 1760
rect 440142 1748 440148 1760
rect 394200 1720 440148 1748
rect 394200 1708 394206 1720
rect 440142 1708 440148 1720
rect 440200 1708 440206 1760
rect 440510 1708 440516 1760
rect 440568 1748 440574 1760
rect 475286 1748 475292 1760
rect 440568 1720 475292 1748
rect 440568 1708 440574 1720
rect 475286 1708 475292 1720
rect 475344 1708 475350 1760
rect 185912 1652 193214 1680
rect 185912 1640 185918 1652
rect 282362 1640 282368 1692
rect 282420 1680 282426 1692
rect 291194 1680 291200 1692
rect 282420 1652 291200 1680
rect 282420 1640 282426 1652
rect 291194 1640 291200 1652
rect 291252 1640 291258 1692
rect 314286 1640 314292 1692
rect 314344 1680 314350 1692
rect 361574 1680 361580 1692
rect 314344 1652 361580 1680
rect 314344 1640 314350 1652
rect 361574 1640 361580 1652
rect 361632 1640 361638 1692
rect 368382 1640 368388 1692
rect 368440 1680 368446 1692
rect 400398 1680 400404 1692
rect 368440 1652 400404 1680
rect 368440 1640 368446 1652
rect 400398 1640 400404 1652
rect 400456 1640 400462 1692
rect 427630 1640 427636 1692
rect 427688 1680 427694 1692
rect 445570 1680 445576 1692
rect 427688 1652 445576 1680
rect 427688 1640 427694 1652
rect 445570 1640 445576 1652
rect 445628 1640 445634 1692
rect 448238 1640 448244 1692
rect 448296 1680 448302 1692
rect 477494 1680 477500 1692
rect 448296 1652 477500 1680
rect 448296 1640 448302 1652
rect 477494 1640 477500 1652
rect 477552 1640 477558 1692
rect 115256 1584 133184 1612
rect 115256 1572 115262 1584
rect 137002 1572 137008 1624
rect 137060 1612 137066 1624
rect 138106 1612 138112 1624
rect 137060 1584 138112 1612
rect 137060 1572 137066 1584
rect 138106 1572 138112 1584
rect 138164 1572 138170 1624
rect 144730 1612 144736 1624
rect 141344 1584 144736 1612
rect 63678 1544 63684 1556
rect 61120 1516 63684 1544
rect 50522 1476 50528 1488
rect 48884 1448 50528 1476
rect 42794 1408 42800 1420
rect 41386 1380 42800 1408
rect 19242 1340 19248 1352
rect 17420 1312 19248 1340
rect 14274 1136 14280 1148
rect 12056 1108 14280 1136
rect 4154 864 4160 876
rect 3252 836 4160 864
rect 74 796 130 800
rect 842 796 848 808
rect 74 768 848 796
rect 74 0 130 768
rect 842 756 848 768
rect 900 756 906 808
rect 1162 796 1218 800
rect 1302 796 1308 808
rect 1162 768 1308 796
rect 1162 0 1218 768
rect 1302 756 1308 768
rect 1360 756 1366 808
rect 2250 796 2306 800
rect 3252 796 3280 836
rect 4154 824 4160 836
rect 4212 824 4218 876
rect 5994 864 6000 876
rect 5184 836 6000 864
rect 2250 768 3280 796
rect 3338 796 3394 800
rect 3970 796 3976 808
rect 3338 768 3976 796
rect 2250 0 2306 768
rect 3338 0 3394 768
rect 3970 756 3976 768
rect 4028 756 4034 808
rect 4426 796 4482 800
rect 5184 796 5212 836
rect 5994 824 6000 836
rect 6052 824 6058 876
rect 11330 864 11336 876
rect 10888 836 11336 864
rect 4426 768 5212 796
rect 5514 796 5570 800
rect 6178 796 6184 808
rect 5514 768 6184 796
rect 4426 0 4482 768
rect 5514 0 5570 768
rect 6178 756 6184 768
rect 6236 756 6242 808
rect 6602 796 6658 800
rect 6730 796 6736 808
rect 6602 768 6736 796
rect 6602 0 6658 768
rect 6730 756 6736 768
rect 6788 756 6794 808
rect 7690 796 7746 800
rect 8478 796 8484 808
rect 7690 768 8484 796
rect 7690 0 7746 768
rect 8478 756 8484 768
rect 8536 756 8542 808
rect 8778 796 8834 800
rect 9582 796 9588 808
rect 8778 768 9588 796
rect 8778 0 8834 768
rect 9582 756 9588 768
rect 9640 756 9646 808
rect 9866 796 9922 800
rect 10888 796 10916 836
rect 11330 824 11336 836
rect 11388 824 11394 876
rect 12056 864 12084 1108
rect 14274 1096 14280 1108
rect 14332 1096 14338 1148
rect 17310 1000 17316 1012
rect 13924 972 17316 1000
rect 12056 836 12204 864
rect 9866 768 10916 796
rect 9866 0 9922 768
rect 10778 688 10784 740
rect 10836 728 10842 740
rect 10954 728 11010 800
rect 10836 700 11010 728
rect 10836 688 10842 700
rect 10954 0 11010 700
rect 12042 796 12098 800
rect 12176 796 12204 836
rect 12042 768 12204 796
rect 12042 0 12098 768
rect 13130 728 13186 800
rect 13924 728 13952 972
rect 17310 960 17316 972
rect 17368 960 17374 1012
rect 16574 932 16580 944
rect 14246 904 16580 932
rect 14246 864 14274 904
rect 16574 892 16580 904
rect 16632 892 16638 944
rect 17420 932 17448 1312
rect 19242 1300 19248 1312
rect 19300 1300 19306 1352
rect 29086 1300 29092 1352
rect 29144 1340 29150 1352
rect 29144 1312 33456 1340
rect 29144 1300 29150 1312
rect 20714 1272 20720 1284
rect 17328 904 17448 932
rect 17496 1244 20720 1272
rect 17496 932 17524 1244
rect 20714 1232 20720 1244
rect 20772 1232 20778 1284
rect 24762 1232 24768 1284
rect 24820 1272 24826 1284
rect 28258 1272 28264 1284
rect 24820 1244 28264 1272
rect 24820 1232 24826 1244
rect 28258 1232 28264 1244
rect 28316 1232 28322 1284
rect 33428 1272 33456 1312
rect 33502 1300 33508 1352
rect 33560 1340 33566 1352
rect 38654 1340 38660 1352
rect 33560 1312 38660 1340
rect 33560 1300 33566 1312
rect 38654 1300 38660 1312
rect 38712 1300 38718 1352
rect 34790 1272 34796 1284
rect 33428 1244 34796 1272
rect 34790 1232 34796 1244
rect 34848 1232 34854 1284
rect 35710 1232 35716 1284
rect 35768 1272 35774 1284
rect 41386 1272 41414 1380
rect 42794 1368 42800 1380
rect 42852 1368 42858 1420
rect 42150 1300 42156 1352
rect 42208 1340 42214 1352
rect 48884 1340 48912 1448
rect 50522 1436 50528 1448
rect 50580 1436 50586 1488
rect 51902 1436 51908 1488
rect 51960 1476 51966 1488
rect 57882 1476 57888 1488
rect 51960 1448 57888 1476
rect 51960 1436 51966 1448
rect 57882 1436 57888 1448
rect 57940 1436 57946 1488
rect 49694 1408 49700 1420
rect 42208 1312 48912 1340
rect 48976 1380 49700 1408
rect 42208 1300 42214 1312
rect 35768 1244 41414 1272
rect 35768 1232 35774 1244
rect 43254 1232 43260 1284
rect 43312 1272 43318 1284
rect 48976 1272 49004 1380
rect 49694 1368 49700 1380
rect 49752 1368 49758 1420
rect 53834 1408 53840 1420
rect 53760 1380 53840 1408
rect 49050 1300 49056 1352
rect 49108 1340 49114 1352
rect 53760 1340 53788 1380
rect 53834 1368 53840 1380
rect 53892 1368 53898 1420
rect 60550 1368 60556 1420
rect 60608 1408 60614 1420
rect 61120 1408 61148 1516
rect 63678 1504 63684 1516
rect 63736 1504 63742 1556
rect 69474 1504 69480 1556
rect 69532 1544 69538 1556
rect 74534 1544 74540 1556
rect 69532 1516 74540 1544
rect 69532 1504 69538 1516
rect 74534 1504 74540 1516
rect 74592 1504 74598 1556
rect 75730 1504 75736 1556
rect 75788 1544 75794 1556
rect 81526 1544 81532 1556
rect 75788 1516 81532 1544
rect 75788 1504 75794 1516
rect 81526 1504 81532 1516
rect 81584 1504 81590 1556
rect 84286 1504 84292 1556
rect 84344 1544 84350 1556
rect 118694 1544 118700 1556
rect 84344 1516 118700 1544
rect 84344 1504 84350 1516
rect 118694 1504 118700 1516
rect 118752 1504 118758 1556
rect 118786 1504 118792 1556
rect 118844 1544 118850 1556
rect 124214 1544 124220 1556
rect 118844 1516 124220 1544
rect 118844 1504 118850 1516
rect 124214 1504 124220 1516
rect 124272 1504 124278 1556
rect 136174 1544 136180 1556
rect 132420 1516 136180 1544
rect 62758 1436 62764 1488
rect 62816 1476 62822 1488
rect 64874 1476 64880 1488
rect 62816 1448 64880 1476
rect 62816 1436 62822 1448
rect 64874 1436 64880 1448
rect 64932 1436 64938 1488
rect 66254 1436 66260 1488
rect 66312 1476 66318 1488
rect 118878 1476 118884 1488
rect 66312 1448 118884 1476
rect 66312 1436 66318 1448
rect 118878 1436 118884 1448
rect 118936 1436 118942 1488
rect 119614 1436 119620 1488
rect 119672 1476 119678 1488
rect 125686 1476 125692 1488
rect 119672 1448 125692 1476
rect 119672 1436 119678 1448
rect 125686 1436 125692 1448
rect 125744 1436 125750 1488
rect 126146 1436 126152 1488
rect 126204 1476 126210 1488
rect 126974 1476 126980 1488
rect 126204 1448 126980 1476
rect 126204 1436 126210 1448
rect 126974 1436 126980 1448
rect 127032 1436 127038 1488
rect 128078 1436 128084 1488
rect 128136 1476 128142 1488
rect 132218 1476 132224 1488
rect 128136 1448 132224 1476
rect 128136 1436 128142 1448
rect 132218 1436 132224 1448
rect 132276 1436 132282 1488
rect 67910 1408 67916 1420
rect 60608 1380 61148 1408
rect 63328 1380 63540 1408
rect 60608 1368 60614 1380
rect 49108 1312 53788 1340
rect 49108 1300 49114 1312
rect 56134 1300 56140 1352
rect 56192 1340 56198 1352
rect 60642 1340 60648 1352
rect 56192 1312 60648 1340
rect 56192 1300 56198 1312
rect 60642 1300 60648 1312
rect 60700 1300 60706 1352
rect 60734 1300 60740 1352
rect 60792 1340 60798 1352
rect 63328 1340 63356 1380
rect 60792 1312 63356 1340
rect 63512 1340 63540 1380
rect 65260 1380 67916 1408
rect 65260 1340 65288 1380
rect 67910 1368 67916 1380
rect 67968 1368 67974 1420
rect 71424 1380 73568 1408
rect 63512 1312 65288 1340
rect 60792 1300 60798 1312
rect 66162 1300 66168 1352
rect 66220 1340 66226 1352
rect 71424 1340 71452 1380
rect 66220 1312 71452 1340
rect 66220 1300 66226 1312
rect 71498 1300 71504 1352
rect 71556 1340 71562 1352
rect 73338 1340 73344 1352
rect 71556 1312 73344 1340
rect 71556 1300 71562 1312
rect 73338 1300 73344 1312
rect 73396 1300 73402 1352
rect 43312 1244 49004 1272
rect 43312 1232 43318 1244
rect 49786 1232 49792 1284
rect 49844 1272 49850 1284
rect 53742 1272 53748 1284
rect 49844 1244 53748 1272
rect 49844 1232 49850 1244
rect 53742 1232 53748 1244
rect 53800 1232 53806 1284
rect 53944 1244 55444 1272
rect 21634 1204 21640 1216
rect 18570 1176 21640 1204
rect 17496 904 17632 932
rect 17328 864 17356 904
rect 14200 836 14274 864
rect 16546 836 17356 864
rect 14200 800 14228 836
rect 14200 768 14274 800
rect 13130 700 13952 728
rect 13130 0 13186 700
rect 14218 0 14274 768
rect 15306 796 15362 800
rect 15930 796 15936 808
rect 15306 768 15936 796
rect 15306 0 15362 768
rect 15930 756 15936 768
rect 15988 756 15994 808
rect 16394 796 16450 800
rect 16546 796 16574 836
rect 16394 768 16574 796
rect 17482 796 17538 800
rect 17604 796 17632 904
rect 18570 864 18598 1176
rect 21634 1164 21640 1176
rect 21692 1164 21698 1216
rect 27614 1204 27620 1216
rect 24044 1176 27620 1204
rect 23934 1136 23940 1148
rect 19674 1108 23940 1136
rect 19674 932 19702 1108
rect 23934 1096 23940 1108
rect 23992 1096 23998 1148
rect 23842 1068 23848 1080
rect 20760 1040 23848 1068
rect 19674 904 19840 932
rect 18570 836 18644 864
rect 18616 800 18644 836
rect 17482 768 17632 796
rect 18570 768 18644 800
rect 19658 796 19714 800
rect 19812 796 19840 904
rect 20760 864 20788 1040
rect 23842 1028 23848 1040
rect 23900 1028 23906 1080
rect 24044 932 24072 1176
rect 27614 1164 27620 1176
rect 27672 1164 27678 1216
rect 28902 1204 28908 1216
rect 27724 1176 28908 1204
rect 27724 1136 27752 1176
rect 28902 1164 28908 1176
rect 28960 1164 28966 1216
rect 53558 1204 53564 1216
rect 46584 1176 53564 1204
rect 32766 1136 32772 1148
rect 19658 768 19840 796
rect 20640 836 20788 864
rect 22066 904 24072 932
rect 25102 1108 27752 1136
rect 31726 1108 32772 1136
rect 20640 796 20668 836
rect 20746 796 20802 800
rect 20640 768 20802 796
rect 16394 0 16450 768
rect 17482 0 17538 768
rect 18570 0 18626 768
rect 19658 0 19714 768
rect 20746 0 20802 768
rect 21834 796 21890 800
rect 22066 796 22094 904
rect 24854 864 24860 876
rect 23308 836 24860 864
rect 21834 768 22094 796
rect 22922 796 22978 800
rect 23308 796 23336 836
rect 24854 824 24860 836
rect 24912 824 24918 876
rect 25102 864 25130 1108
rect 31726 1068 31754 1108
rect 32766 1096 32772 1108
rect 32824 1096 32830 1148
rect 37826 1096 37832 1148
rect 37884 1136 37890 1148
rect 44082 1136 44088 1148
rect 37884 1108 44088 1136
rect 37884 1096 37890 1108
rect 44082 1096 44088 1108
rect 44140 1096 44146 1148
rect 37458 1068 37464 1080
rect 26206 1040 31754 1068
rect 32324 1040 37464 1068
rect 26206 864 26234 1040
rect 31846 1000 31852 1012
rect 29472 972 31852 1000
rect 29362 932 29368 944
rect 25102 836 25176 864
rect 22922 768 23336 796
rect 24010 796 24066 800
rect 24762 796 24768 808
rect 24010 768 24768 796
rect 21834 0 21890 768
rect 22922 0 22978 768
rect 24010 0 24066 768
rect 24762 756 24768 768
rect 24820 756 24826 808
rect 25148 800 25176 836
rect 25098 768 25176 800
rect 26160 836 26234 864
rect 28000 904 29368 932
rect 26160 800 26188 836
rect 25098 0 25154 768
rect 26160 700 26242 800
rect 26186 0 26242 700
rect 27274 728 27330 800
rect 28000 728 28028 904
rect 29362 892 29368 904
rect 29420 892 29426 944
rect 29472 864 29500 972
rect 31846 960 31852 972
rect 31904 960 31910 1012
rect 32324 864 32352 1040
rect 37458 1028 37464 1040
rect 37516 1028 37522 1080
rect 39114 1068 39120 1080
rect 37660 1040 39120 1068
rect 33134 932 33140 944
rect 29472 836 29592 864
rect 27274 700 28028 728
rect 28362 796 28418 800
rect 29086 796 29092 808
rect 28362 768 29092 796
rect 27274 0 27330 700
rect 28362 0 28418 768
rect 29086 756 29092 768
rect 29144 756 29150 808
rect 29450 796 29506 800
rect 29564 796 29592 836
rect 31128 836 32352 864
rect 32416 904 33140 932
rect 29450 768 29592 796
rect 30538 796 30594 800
rect 31128 796 31156 836
rect 30538 768 31156 796
rect 31626 796 31682 800
rect 32416 796 32444 904
rect 33134 892 33140 904
rect 33192 892 33198 944
rect 36814 932 36820 944
rect 34624 904 36820 932
rect 31626 768 32444 796
rect 29450 0 29506 768
rect 30538 0 30594 768
rect 31626 0 31682 768
rect 32714 728 32770 800
rect 33802 796 33858 800
rect 34624 796 34652 904
rect 36814 892 36820 904
rect 36872 892 36878 944
rect 37660 932 37688 1040
rect 39114 1028 39120 1040
rect 39172 1028 39178 1080
rect 40862 1028 40868 1080
rect 40920 1068 40926 1080
rect 43162 1068 43168 1080
rect 40920 1040 43168 1068
rect 40920 1028 40926 1040
rect 43162 1028 43168 1040
rect 43220 1028 43226 1080
rect 41322 1000 41328 1012
rect 36924 904 37688 932
rect 38948 972 41328 1000
rect 33802 768 34652 796
rect 34890 796 34946 800
rect 35710 796 35716 808
rect 34890 768 35716 796
rect 33502 728 33508 740
rect 32714 700 33508 728
rect 32714 0 32770 700
rect 33502 688 33508 700
rect 33560 688 33566 740
rect 33802 0 33858 768
rect 34890 0 34946 768
rect 35710 756 35716 768
rect 35768 756 35774 808
rect 35978 796 36034 800
rect 36924 796 36952 904
rect 35978 768 36952 796
rect 37066 796 37122 800
rect 37826 796 37832 808
rect 37066 768 37832 796
rect 35978 0 36034 768
rect 37066 0 37122 768
rect 37826 756 37832 768
rect 37884 756 37890 808
rect 38154 728 38210 800
rect 38948 728 38976 972
rect 41322 960 41328 972
rect 41380 960 41386 1012
rect 46014 1000 46020 1012
rect 43364 972 46020 1000
rect 39270 904 41414 932
rect 39270 864 39298 904
rect 39224 836 39298 864
rect 41386 864 41414 904
rect 43364 864 43392 972
rect 46014 960 46020 972
rect 46072 960 46078 1012
rect 46584 932 46612 1176
rect 53558 1164 53564 1176
rect 53616 1164 53622 1216
rect 53944 1204 53972 1244
rect 53852 1176 53972 1204
rect 55416 1204 55444 1244
rect 56226 1232 56232 1284
rect 56284 1272 56290 1284
rect 58986 1272 58992 1284
rect 56284 1244 58992 1272
rect 56284 1232 56290 1244
rect 58986 1232 58992 1244
rect 59044 1232 59050 1284
rect 59630 1232 59636 1284
rect 59688 1272 59694 1284
rect 63218 1272 63224 1284
rect 59688 1244 63224 1272
rect 59688 1232 59694 1244
rect 63218 1232 63224 1244
rect 63276 1232 63282 1284
rect 68554 1272 68560 1284
rect 63420 1244 68560 1272
rect 57974 1204 57980 1216
rect 55416 1176 57980 1204
rect 47670 1096 47676 1148
rect 47728 1136 47734 1148
rect 48958 1136 48964 1148
rect 47728 1108 48964 1136
rect 47728 1096 47734 1108
rect 48958 1096 48964 1108
rect 49016 1096 49022 1148
rect 49050 1096 49056 1148
rect 49108 1136 49114 1148
rect 53852 1136 53880 1176
rect 57974 1164 57980 1176
rect 58032 1164 58038 1216
rect 58526 1164 58532 1216
rect 58584 1204 58590 1216
rect 62758 1204 62764 1216
rect 58584 1176 62764 1204
rect 58584 1164 58590 1176
rect 62758 1164 62764 1176
rect 62816 1164 62822 1216
rect 49108 1108 53880 1136
rect 49108 1096 49114 1108
rect 54018 1096 54024 1148
rect 54076 1136 54082 1148
rect 56686 1136 56692 1148
rect 54076 1108 56692 1136
rect 54076 1096 54082 1108
rect 56686 1096 56692 1108
rect 56744 1096 56750 1148
rect 57422 1096 57428 1148
rect 57480 1136 57486 1148
rect 63420 1136 63448 1244
rect 68554 1232 68560 1244
rect 68612 1232 68618 1284
rect 73430 1272 73436 1284
rect 69584 1244 73436 1272
rect 63586 1164 63592 1216
rect 63644 1204 63650 1216
rect 66714 1204 66720 1216
rect 63644 1176 66720 1204
rect 63644 1164 63650 1176
rect 66714 1164 66720 1176
rect 66772 1164 66778 1216
rect 66806 1164 66812 1216
rect 66864 1204 66870 1216
rect 69474 1204 69480 1216
rect 66864 1176 69480 1204
rect 66864 1164 66870 1176
rect 69474 1164 69480 1176
rect 69532 1164 69538 1216
rect 57480 1108 63448 1136
rect 57480 1096 57486 1108
rect 63954 1096 63960 1148
rect 64012 1136 64018 1148
rect 69584 1136 69612 1244
rect 73430 1232 73436 1244
rect 73488 1232 73494 1284
rect 69658 1164 69664 1216
rect 69716 1204 69722 1216
rect 73540 1204 73568 1380
rect 73614 1368 73620 1420
rect 73672 1368 73678 1420
rect 86770 1408 86776 1420
rect 77220 1380 86776 1408
rect 73632 1340 73660 1368
rect 74902 1340 74908 1352
rect 73632 1312 74908 1340
rect 74902 1300 74908 1312
rect 74960 1300 74966 1352
rect 74994 1300 75000 1352
rect 75052 1340 75058 1352
rect 77220 1340 77248 1380
rect 86770 1368 86776 1380
rect 86828 1368 86834 1420
rect 94130 1368 94136 1420
rect 94188 1408 94194 1420
rect 94188 1380 94360 1408
rect 94188 1368 94194 1380
rect 75052 1312 77248 1340
rect 75052 1300 75058 1312
rect 78030 1300 78036 1352
rect 78088 1340 78094 1352
rect 89714 1340 89720 1352
rect 78088 1312 89720 1340
rect 78088 1300 78094 1312
rect 89714 1300 89720 1312
rect 89772 1300 89778 1352
rect 89806 1300 89812 1352
rect 89864 1340 89870 1352
rect 92566 1340 92572 1352
rect 89864 1312 92572 1340
rect 89864 1300 89870 1312
rect 92566 1300 92572 1312
rect 92624 1300 92630 1352
rect 94332 1340 94360 1380
rect 95436 1380 101076 1408
rect 95436 1340 95464 1380
rect 94332 1312 95464 1340
rect 95510 1300 95516 1352
rect 95568 1340 95574 1352
rect 99006 1340 99012 1352
rect 95568 1312 99012 1340
rect 95568 1300 95574 1312
rect 99006 1300 99012 1312
rect 99064 1300 99070 1352
rect 73614 1232 73620 1284
rect 73672 1272 73678 1284
rect 75454 1272 75460 1284
rect 73672 1244 75460 1272
rect 73672 1232 73678 1244
rect 75454 1232 75460 1244
rect 75512 1232 75518 1284
rect 77202 1272 77208 1284
rect 76116 1244 77208 1272
rect 76116 1204 76144 1244
rect 77202 1232 77208 1244
rect 77260 1232 77266 1284
rect 79134 1232 79140 1284
rect 79192 1272 79198 1284
rect 79192 1244 80054 1272
rect 79192 1232 79198 1244
rect 69716 1176 73384 1204
rect 73540 1176 76144 1204
rect 80026 1204 80054 1244
rect 80146 1232 80152 1284
rect 80204 1272 80210 1284
rect 84102 1272 84108 1284
rect 80204 1244 84108 1272
rect 80204 1232 80210 1244
rect 84102 1232 84108 1244
rect 84160 1232 84166 1284
rect 85758 1232 85764 1284
rect 85816 1272 85822 1284
rect 85816 1244 89668 1272
rect 85816 1232 85822 1244
rect 87046 1204 87052 1216
rect 80026 1176 87052 1204
rect 69716 1164 69722 1176
rect 64012 1108 69612 1136
rect 64012 1096 64018 1108
rect 70486 1096 70492 1148
rect 70544 1136 70550 1148
rect 73356 1136 73384 1176
rect 87046 1164 87052 1176
rect 87104 1164 87110 1216
rect 89640 1204 89668 1244
rect 89898 1232 89904 1284
rect 89956 1272 89962 1284
rect 99098 1272 99104 1284
rect 89956 1244 99104 1272
rect 89956 1232 89962 1244
rect 99098 1232 99104 1244
rect 99156 1232 99162 1284
rect 101048 1272 101076 1380
rect 105262 1368 105268 1420
rect 105320 1408 105326 1420
rect 107746 1408 107752 1420
rect 105320 1380 107752 1408
rect 105320 1368 105326 1380
rect 107746 1368 107752 1380
rect 107804 1368 107810 1420
rect 110322 1408 110328 1420
rect 108960 1380 110328 1408
rect 101122 1300 101128 1352
rect 101180 1340 101186 1352
rect 108960 1340 108988 1380
rect 110322 1368 110328 1380
rect 110380 1368 110386 1420
rect 110782 1368 110788 1420
rect 110840 1408 110846 1420
rect 132420 1408 132448 1516
rect 136174 1504 136180 1516
rect 136232 1504 136238 1556
rect 132494 1436 132500 1488
rect 132552 1476 132558 1488
rect 141344 1476 141372 1584
rect 144730 1572 144736 1584
rect 144788 1572 144794 1624
rect 146202 1572 146208 1624
rect 146260 1612 146266 1624
rect 148502 1612 148508 1624
rect 146260 1584 148508 1612
rect 146260 1572 146266 1584
rect 148502 1572 148508 1584
rect 148560 1572 148566 1624
rect 148594 1572 148600 1624
rect 148652 1612 148658 1624
rect 252462 1612 252468 1624
rect 148652 1584 252468 1612
rect 148652 1572 148658 1584
rect 252462 1572 252468 1584
rect 252520 1572 252526 1624
rect 262398 1572 262404 1624
rect 262456 1612 262462 1624
rect 264974 1612 264980 1624
rect 262456 1584 264980 1612
rect 262456 1572 262462 1584
rect 264974 1572 264980 1584
rect 265032 1572 265038 1624
rect 278222 1572 278228 1624
rect 278280 1612 278286 1624
rect 283098 1612 283104 1624
rect 278280 1584 283104 1612
rect 278280 1572 278286 1584
rect 283098 1572 283104 1584
rect 283156 1572 283162 1624
rect 345198 1572 345204 1624
rect 345256 1612 345262 1624
rect 389174 1612 389180 1624
rect 345256 1584 389180 1612
rect 345256 1572 345262 1584
rect 389174 1572 389180 1584
rect 389232 1572 389238 1624
rect 396718 1572 396724 1624
rect 396776 1612 396782 1624
rect 440970 1612 440976 1624
rect 396776 1584 440976 1612
rect 396776 1572 396782 1584
rect 440970 1572 440976 1584
rect 441028 1572 441034 1624
rect 473906 1572 473912 1624
rect 473964 1612 473970 1624
rect 484210 1612 484216 1624
rect 473964 1584 484216 1612
rect 473964 1572 473970 1584
rect 484210 1572 484216 1584
rect 484268 1572 484274 1624
rect 141418 1504 141424 1556
rect 141476 1544 141482 1556
rect 148226 1544 148232 1556
rect 141476 1516 148232 1544
rect 141476 1504 141482 1516
rect 148226 1504 148232 1516
rect 148284 1504 148290 1556
rect 150342 1504 150348 1556
rect 150400 1544 150406 1556
rect 161566 1544 161572 1556
rect 150400 1516 161572 1544
rect 150400 1504 150406 1516
rect 161566 1504 161572 1516
rect 161624 1504 161630 1556
rect 161750 1504 161756 1556
rect 161808 1544 161814 1556
rect 166810 1544 166816 1556
rect 161808 1516 166816 1544
rect 161808 1504 161814 1516
rect 166810 1504 166816 1516
rect 166868 1504 166874 1556
rect 167454 1504 167460 1556
rect 167512 1544 167518 1556
rect 174630 1544 174636 1556
rect 167512 1516 174636 1544
rect 167512 1504 167518 1516
rect 174630 1504 174636 1516
rect 174688 1504 174694 1556
rect 174814 1504 174820 1556
rect 174872 1544 174878 1556
rect 179506 1544 179512 1556
rect 174872 1516 179512 1544
rect 174872 1504 174878 1516
rect 179506 1504 179512 1516
rect 179564 1504 179570 1556
rect 179598 1504 179604 1556
rect 179656 1544 179662 1556
rect 259914 1544 259920 1556
rect 179656 1516 259920 1544
rect 179656 1504 179662 1516
rect 259914 1504 259920 1516
rect 259972 1504 259978 1556
rect 273990 1504 273996 1556
rect 274048 1544 274054 1556
rect 282270 1544 282276 1556
rect 274048 1516 282276 1544
rect 274048 1504 274054 1516
rect 282270 1504 282276 1516
rect 282328 1504 282334 1556
rect 282546 1504 282552 1556
rect 282604 1544 282610 1556
rect 285674 1544 285680 1556
rect 282604 1516 285680 1544
rect 282604 1504 282610 1516
rect 285674 1504 285680 1516
rect 285732 1504 285738 1556
rect 293494 1504 293500 1556
rect 293552 1544 293558 1556
rect 300854 1544 300860 1556
rect 293552 1516 300860 1544
rect 293552 1504 293558 1516
rect 300854 1504 300860 1516
rect 300912 1504 300918 1556
rect 324590 1504 324596 1556
rect 324648 1544 324654 1556
rect 372614 1544 372620 1556
rect 324648 1516 372620 1544
rect 324648 1504 324654 1516
rect 372614 1504 372620 1516
rect 372672 1504 372678 1556
rect 381262 1504 381268 1556
rect 381320 1544 381326 1556
rect 417050 1544 417056 1556
rect 381320 1516 417056 1544
rect 381320 1504 381326 1516
rect 417050 1504 417056 1516
rect 417108 1504 417114 1556
rect 432782 1504 432788 1556
rect 432840 1544 432846 1556
rect 456794 1544 456800 1556
rect 432840 1516 456800 1544
rect 432840 1504 432846 1516
rect 456794 1504 456800 1516
rect 456852 1504 456858 1556
rect 132552 1448 141372 1476
rect 132552 1436 132558 1448
rect 143718 1436 143724 1488
rect 143776 1476 143782 1488
rect 147766 1476 147772 1488
rect 143776 1448 147772 1476
rect 143776 1436 143782 1448
rect 147766 1436 147772 1448
rect 147824 1436 147830 1488
rect 147858 1436 147864 1488
rect 147916 1476 147922 1488
rect 153378 1476 153384 1488
rect 147916 1448 153384 1476
rect 147916 1436 147922 1448
rect 153378 1436 153384 1448
rect 153436 1436 153442 1488
rect 154574 1436 154580 1488
rect 154632 1476 154638 1488
rect 156414 1476 156420 1488
rect 154632 1448 156420 1476
rect 154632 1436 154638 1448
rect 156414 1436 156420 1448
rect 156472 1436 156478 1488
rect 157306 1448 168620 1476
rect 110840 1380 132448 1408
rect 110840 1368 110846 1380
rect 132586 1368 132592 1420
rect 132644 1408 132650 1420
rect 144914 1408 144920 1420
rect 132644 1380 144920 1408
rect 132644 1368 132650 1380
rect 144914 1368 144920 1380
rect 144972 1368 144978 1420
rect 146662 1368 146668 1420
rect 146720 1408 146726 1420
rect 157306 1408 157334 1448
rect 146720 1380 157334 1408
rect 146720 1368 146726 1380
rect 157426 1368 157432 1420
rect 157484 1408 157490 1420
rect 166718 1408 166724 1420
rect 157484 1380 166724 1408
rect 157484 1368 157490 1380
rect 166718 1368 166724 1380
rect 166776 1368 166782 1420
rect 166810 1368 166816 1420
rect 166868 1408 166874 1420
rect 166994 1408 167000 1420
rect 166868 1380 167000 1408
rect 166868 1368 166874 1380
rect 166994 1368 167000 1380
rect 167052 1368 167058 1420
rect 168592 1408 168620 1448
rect 168650 1436 168656 1488
rect 168708 1476 168714 1488
rect 176746 1476 176752 1488
rect 168708 1448 176752 1476
rect 168708 1436 168714 1448
rect 176746 1436 176752 1448
rect 176804 1436 176810 1488
rect 176930 1436 176936 1488
rect 176988 1476 176994 1488
rect 181070 1476 181076 1488
rect 176988 1448 181076 1476
rect 176988 1436 176994 1448
rect 181070 1436 181076 1448
rect 181128 1436 181134 1488
rect 181346 1436 181352 1488
rect 181404 1476 181410 1488
rect 182174 1476 182180 1488
rect 181404 1448 182180 1476
rect 181404 1436 181410 1448
rect 182174 1436 182180 1448
rect 182232 1436 182238 1488
rect 183526 1448 184060 1476
rect 183526 1408 183554 1448
rect 167104 1380 167316 1408
rect 168592 1380 183554 1408
rect 101180 1312 108988 1340
rect 101180 1300 101186 1312
rect 109034 1300 109040 1352
rect 109092 1340 109098 1352
rect 113174 1340 113180 1352
rect 109092 1312 113180 1340
rect 109092 1300 109098 1312
rect 113174 1300 113180 1312
rect 113232 1300 113238 1352
rect 113634 1300 113640 1352
rect 113692 1340 113698 1352
rect 167104 1340 167132 1380
rect 113692 1312 167132 1340
rect 167288 1340 167316 1380
rect 183646 1368 183652 1420
rect 183704 1368 183710 1420
rect 184032 1408 184060 1448
rect 186682 1436 186688 1488
rect 186740 1476 186746 1488
rect 188338 1476 188344 1488
rect 186740 1448 188344 1476
rect 186740 1436 186746 1448
rect 188338 1436 188344 1448
rect 188396 1436 188402 1488
rect 190178 1436 190184 1488
rect 190236 1476 190242 1488
rect 195238 1476 195244 1488
rect 190236 1448 195244 1476
rect 190236 1436 190242 1448
rect 195238 1436 195244 1448
rect 195296 1436 195302 1488
rect 195330 1436 195336 1488
rect 195388 1476 195394 1488
rect 262306 1476 262312 1488
rect 195388 1448 262312 1476
rect 195388 1436 195394 1448
rect 262306 1436 262312 1448
rect 262364 1436 262370 1488
rect 271598 1436 271604 1488
rect 271656 1476 271662 1488
rect 273346 1476 273352 1488
rect 271656 1448 273352 1476
rect 271656 1436 271662 1448
rect 273346 1436 273352 1448
rect 273404 1436 273410 1488
rect 282914 1436 282920 1488
rect 282972 1476 282978 1488
rect 295242 1476 295248 1488
rect 282972 1448 295248 1476
rect 282972 1436 282978 1448
rect 295242 1436 295248 1448
rect 295300 1436 295306 1488
rect 302510 1436 302516 1488
rect 302568 1476 302574 1488
rect 306374 1476 306380 1488
rect 302568 1448 306380 1476
rect 302568 1436 302574 1448
rect 306374 1436 306380 1448
rect 306432 1436 306438 1488
rect 313366 1436 313372 1488
rect 313424 1476 313430 1488
rect 316678 1476 316684 1488
rect 313424 1448 316684 1476
rect 313424 1436 313430 1448
rect 316678 1436 316684 1448
rect 316736 1436 316742 1488
rect 319438 1436 319444 1488
rect 319496 1476 319502 1488
rect 367922 1476 367928 1488
rect 319496 1448 367928 1476
rect 319496 1436 319502 1448
rect 367922 1436 367928 1448
rect 367980 1436 367986 1488
rect 370958 1436 370964 1488
rect 371016 1476 371022 1488
rect 395430 1476 395436 1488
rect 371016 1448 395436 1476
rect 371016 1436 371022 1448
rect 395430 1436 395436 1448
rect 395488 1436 395494 1488
rect 407022 1436 407028 1488
rect 407080 1476 407086 1488
rect 442902 1476 442908 1488
rect 407080 1448 442908 1476
rect 407080 1436 407086 1448
rect 442902 1436 442908 1448
rect 442960 1436 442966 1488
rect 249518 1408 249524 1420
rect 184032 1380 249524 1408
rect 249518 1368 249524 1380
rect 249576 1368 249582 1420
rect 254946 1408 254952 1420
rect 254320 1380 254952 1408
rect 183664 1340 183692 1368
rect 167288 1312 183692 1340
rect 113692 1300 113698 1312
rect 183806 1300 183812 1352
rect 183864 1300 183870 1352
rect 184014 1300 184020 1352
rect 184072 1340 184078 1352
rect 208210 1340 208216 1352
rect 184072 1312 208216 1340
rect 184072 1300 184078 1312
rect 208210 1300 208216 1312
rect 208268 1300 208274 1352
rect 219618 1300 219624 1352
rect 219676 1340 219682 1352
rect 226058 1340 226064 1352
rect 219676 1312 226064 1340
rect 219676 1300 219682 1312
rect 226058 1300 226064 1312
rect 226116 1300 226122 1352
rect 228450 1300 228456 1352
rect 228508 1340 228514 1352
rect 233234 1340 233240 1352
rect 228508 1312 233240 1340
rect 228508 1300 228514 1312
rect 233234 1300 233240 1312
rect 233292 1300 233298 1352
rect 234982 1300 234988 1352
rect 235040 1340 235046 1352
rect 243998 1340 244004 1352
rect 235040 1312 244004 1340
rect 235040 1300 235046 1312
rect 243998 1300 244004 1312
rect 244056 1300 244062 1352
rect 254320 1340 254348 1380
rect 254946 1368 254952 1380
rect 255004 1368 255010 1420
rect 261202 1368 261208 1420
rect 261260 1408 261266 1420
rect 261260 1380 263548 1408
rect 261260 1368 261266 1380
rect 258074 1340 258080 1352
rect 246684 1312 254348 1340
rect 254412 1312 258080 1340
rect 106366 1272 106372 1284
rect 101048 1244 106372 1272
rect 106366 1232 106372 1244
rect 106424 1232 106430 1284
rect 106550 1232 106556 1284
rect 106608 1272 106614 1284
rect 118694 1272 118700 1284
rect 106608 1244 118700 1272
rect 106608 1232 106614 1244
rect 118694 1232 118700 1244
rect 118752 1232 118758 1284
rect 126882 1272 126888 1284
rect 123496 1244 126888 1272
rect 89806 1204 89812 1216
rect 89640 1176 89812 1204
rect 89806 1164 89812 1176
rect 89864 1164 89870 1216
rect 99190 1204 99196 1216
rect 89916 1176 99196 1204
rect 75730 1136 75736 1148
rect 70544 1108 73292 1136
rect 73356 1108 75736 1136
rect 70544 1096 70550 1108
rect 47854 1068 47860 1080
rect 41386 836 43392 864
rect 43594 904 46612 932
rect 46676 1040 47860 1068
rect 43594 864 43622 904
rect 46676 864 46704 1040
rect 47854 1028 47860 1040
rect 47912 1028 47918 1080
rect 59354 1068 59360 1080
rect 49988 1040 50844 1068
rect 48038 960 48044 1012
rect 48096 1000 48102 1012
rect 49988 1000 50016 1040
rect 48096 972 50016 1000
rect 50816 1000 50844 1040
rect 52932 1040 59360 1068
rect 52730 1000 52736 1012
rect 50816 972 52736 1000
rect 48096 960 48102 972
rect 52730 960 52736 972
rect 52788 960 52794 1012
rect 52638 932 52644 944
rect 48056 904 52644 932
rect 48056 864 48084 904
rect 52638 892 52644 904
rect 52696 892 52702 944
rect 48866 864 48872 876
rect 43594 836 43668 864
rect 39224 800 39252 836
rect 39224 768 39298 800
rect 38154 700 38976 728
rect 38154 0 38210 700
rect 39242 0 39298 768
rect 40330 796 40386 800
rect 40862 796 40868 808
rect 40330 768 40868 796
rect 40330 0 40386 768
rect 40862 756 40868 768
rect 40920 756 40926 808
rect 41418 796 41474 800
rect 42150 796 42156 808
rect 41418 768 42156 796
rect 41418 0 41474 768
rect 42150 756 42156 768
rect 42208 756 42214 808
rect 42506 796 42562 800
rect 43254 796 43260 808
rect 42506 768 43260 796
rect 42506 0 42562 768
rect 43254 756 43260 768
rect 43312 756 43318 808
rect 43640 800 43668 836
rect 45526 836 46704 864
rect 46768 836 48084 864
rect 48792 836 48872 864
rect 43594 768 43668 800
rect 44682 796 44738 800
rect 45526 796 45554 836
rect 44682 768 45554 796
rect 45770 796 45826 800
rect 46768 796 46796 836
rect 45770 768 46796 796
rect 46858 796 46914 800
rect 47670 796 47676 808
rect 46858 768 47676 796
rect 43594 0 43650 768
rect 44682 0 44738 768
rect 45770 0 45826 768
rect 46858 0 46914 768
rect 47670 756 47676 768
rect 47728 756 47734 808
rect 47946 796 48002 800
rect 48792 796 48820 836
rect 48866 824 48872 836
rect 48924 824 48930 876
rect 51902 864 51908 876
rect 50908 836 51908 864
rect 47946 768 48820 796
rect 49034 796 49090 800
rect 49786 796 49792 808
rect 49034 768 49792 796
rect 47946 0 48002 768
rect 49034 0 49090 768
rect 49786 756 49792 768
rect 49844 756 49850 808
rect 50122 728 50178 800
rect 50908 728 50936 836
rect 51902 824 51908 836
rect 51960 824 51966 876
rect 52932 864 52960 1040
rect 59354 1028 59360 1040
rect 59412 1028 59418 1080
rect 61838 1028 61844 1080
rect 61896 1068 61902 1080
rect 61896 1040 68232 1068
rect 61896 1028 61902 1040
rect 60550 1000 60556 1012
rect 54220 972 60556 1000
rect 54220 864 54248 972
rect 60550 960 60556 972
rect 60608 960 60614 1012
rect 63218 960 63224 1012
rect 63276 1000 63282 1012
rect 63276 972 64874 1000
rect 63276 960 63282 972
rect 56134 932 56140 944
rect 52012 836 52960 864
rect 53024 836 54248 864
rect 54312 904 56140 932
rect 50122 700 50936 728
rect 51210 796 51266 800
rect 52012 796 52040 836
rect 51210 768 52040 796
rect 52298 796 52354 800
rect 53024 796 53052 836
rect 52298 768 53052 796
rect 53386 796 53442 800
rect 54312 796 54340 904
rect 56134 892 56140 904
rect 56192 892 56198 944
rect 63494 932 63500 944
rect 56336 904 63500 932
rect 56226 864 56232 876
rect 55232 836 56232 864
rect 53386 768 54340 796
rect 54474 796 54530 800
rect 55232 796 55260 836
rect 56226 824 56232 836
rect 56284 824 56290 876
rect 54474 768 55260 796
rect 55562 796 55618 800
rect 56336 796 56364 904
rect 63494 892 63500 904
rect 63552 892 63558 944
rect 64846 932 64874 972
rect 65058 960 65064 1012
rect 65116 1000 65122 1012
rect 68094 1000 68100 1012
rect 65116 972 68100 1000
rect 65116 960 65122 972
rect 68094 960 68100 972
rect 68152 960 68158 1012
rect 68204 1000 68232 1040
rect 68278 1028 68284 1080
rect 68336 1068 68342 1080
rect 73154 1068 73160 1080
rect 68336 1040 73160 1068
rect 68336 1028 68342 1040
rect 73154 1028 73160 1040
rect 73212 1028 73218 1080
rect 73264 1068 73292 1108
rect 75730 1096 75736 1108
rect 75788 1096 75794 1148
rect 75822 1096 75828 1148
rect 75880 1136 75886 1148
rect 81342 1136 81348 1148
rect 75880 1108 81348 1136
rect 75880 1096 75886 1108
rect 81342 1096 81348 1108
rect 81400 1096 81406 1148
rect 84470 1136 84476 1148
rect 82372 1108 84476 1136
rect 75638 1068 75644 1080
rect 73264 1040 75644 1068
rect 75638 1028 75644 1040
rect 75696 1028 75702 1080
rect 80054 1068 80060 1080
rect 75748 1040 80060 1068
rect 68462 1000 68468 1012
rect 68204 972 68468 1000
rect 68462 960 68468 972
rect 68520 960 68526 1012
rect 68572 972 68784 1000
rect 68572 932 68600 972
rect 64846 904 68600 932
rect 68756 932 68784 972
rect 69842 960 69848 1012
rect 69900 1000 69906 1012
rect 71774 1000 71780 1012
rect 69900 972 71780 1000
rect 69900 960 69906 972
rect 71774 960 71780 972
rect 71832 960 71838 1012
rect 72878 960 72884 1012
rect 72936 960 72942 1012
rect 75748 1000 75776 1040
rect 80054 1028 80060 1040
rect 80112 1028 80118 1080
rect 82372 1000 82400 1108
rect 84470 1096 84476 1108
rect 84528 1096 84534 1148
rect 84654 1096 84660 1148
rect 84712 1136 84718 1148
rect 84712 1108 87092 1136
rect 84712 1096 84718 1108
rect 82446 1028 82452 1080
rect 82504 1068 82510 1080
rect 86862 1068 86868 1080
rect 82504 1040 86868 1068
rect 82504 1028 82510 1040
rect 86862 1028 86868 1040
rect 86920 1028 86926 1080
rect 86954 1000 86960 1012
rect 72988 972 75776 1000
rect 75932 972 82400 1000
rect 82556 972 86960 1000
rect 71406 932 71412 944
rect 68756 904 71412 932
rect 71406 892 71412 904
rect 71464 892 71470 944
rect 72896 932 72924 960
rect 72620 904 72924 932
rect 58986 824 58992 876
rect 59044 864 59050 876
rect 65242 864 65248 876
rect 59044 836 65248 864
rect 59044 824 59050 836
rect 65242 824 65248 836
rect 65300 824 65306 876
rect 68738 824 68744 876
rect 68796 864 68802 876
rect 72620 864 72648 904
rect 72878 864 72884 876
rect 68796 836 72648 864
rect 72712 836 72884 864
rect 68796 824 68802 836
rect 55562 768 56364 796
rect 50122 0 50178 700
rect 51210 0 51266 768
rect 52298 0 52354 768
rect 53386 0 53442 768
rect 54474 0 54530 768
rect 55562 0 55618 768
rect 56650 728 56706 800
rect 57738 796 57794 800
rect 58526 796 58532 808
rect 57738 768 58532 796
rect 57422 728 57428 740
rect 56650 700 57428 728
rect 56650 0 56706 700
rect 57422 688 57428 700
rect 57480 688 57486 740
rect 57738 0 57794 768
rect 58526 756 58532 768
rect 58584 756 58590 808
rect 58826 728 58882 800
rect 59914 796 59970 800
rect 60734 796 60740 808
rect 59914 768 60740 796
rect 59630 728 59636 740
rect 58826 700 59636 728
rect 58826 0 58882 700
rect 59630 688 59636 700
rect 59688 688 59694 740
rect 59914 0 59970 768
rect 60734 756 60740 768
rect 60792 756 60798 808
rect 61002 796 61058 800
rect 61838 796 61844 808
rect 61002 768 61844 796
rect 61002 0 61058 768
rect 61838 756 61844 768
rect 61896 756 61902 808
rect 62090 728 62146 800
rect 63178 796 63234 800
rect 63954 796 63960 808
rect 63178 768 63960 796
rect 62850 728 62856 740
rect 62090 700 62856 728
rect 62090 0 62146 700
rect 62850 688 62856 700
rect 62908 688 62914 740
rect 63178 0 63234 768
rect 63954 756 63960 768
rect 64012 756 64018 808
rect 64266 796 64322 800
rect 65058 796 65064 808
rect 64266 768 65064 796
rect 64266 0 64322 768
rect 65058 756 65064 768
rect 65116 756 65122 808
rect 65354 796 65410 800
rect 66162 796 66168 808
rect 65354 768 66168 796
rect 65354 0 65410 768
rect 66162 756 66168 768
rect 66220 756 66226 808
rect 66442 796 66498 800
rect 66806 796 66812 808
rect 66442 768 66812 796
rect 66442 0 66498 768
rect 66806 756 66812 768
rect 66864 756 66870 808
rect 67530 796 67586 800
rect 68278 796 68284 808
rect 67530 768 68284 796
rect 67530 0 67586 768
rect 68278 756 68284 768
rect 68336 756 68342 808
rect 68618 728 68674 800
rect 69382 728 69388 740
rect 68618 700 69388 728
rect 68618 0 68674 700
rect 69382 688 69388 700
rect 69440 688 69446 740
rect 69706 728 69762 800
rect 70794 796 70850 800
rect 71498 796 71504 808
rect 70794 768 71504 796
rect 70486 728 70492 740
rect 69706 700 70492 728
rect 69706 0 69762 700
rect 70486 688 70492 700
rect 70544 688 70550 740
rect 70794 0 70850 768
rect 71498 756 71504 768
rect 71556 756 71562 808
rect 71882 796 71938 800
rect 72712 796 72740 836
rect 72878 824 72884 836
rect 72936 824 72942 876
rect 72988 864 73016 972
rect 73062 892 73068 944
rect 73120 932 73126 944
rect 75932 932 75960 972
rect 80330 932 80336 944
rect 73120 904 75960 932
rect 76484 904 80336 932
rect 73120 892 73126 904
rect 72988 836 73108 864
rect 71882 768 72740 796
rect 72970 796 73026 800
rect 73080 796 73108 836
rect 73154 824 73160 876
rect 73212 864 73218 876
rect 75822 864 75828 876
rect 73212 836 75828 864
rect 73212 824 73218 836
rect 75822 824 75828 836
rect 75880 824 75886 876
rect 72970 768 73108 796
rect 71882 0 71938 768
rect 72970 0 73026 768
rect 74058 48 74114 800
rect 75146 796 75202 800
rect 75730 796 75736 808
rect 75146 768 75736 796
rect 74994 48 75000 60
rect 74058 20 75000 48
rect 74058 0 74114 20
rect 74994 8 75000 20
rect 75052 8 75058 60
rect 75146 0 75202 768
rect 75730 756 75736 768
rect 75788 756 75794 808
rect 76234 796 76290 800
rect 76484 796 76512 904
rect 80330 892 80336 904
rect 80388 892 80394 944
rect 81434 932 81440 944
rect 80440 904 81440 932
rect 76558 824 76564 876
rect 76616 864 76622 876
rect 80440 864 80468 904
rect 81434 892 81440 904
rect 81492 892 81498 944
rect 82556 864 82584 972
rect 86954 960 86960 972
rect 87012 960 87018 1012
rect 87064 1000 87092 1108
rect 87874 1028 87880 1080
rect 87932 1068 87938 1080
rect 89916 1068 89944 1176
rect 99190 1164 99196 1176
rect 99248 1164 99254 1216
rect 100018 1164 100024 1216
rect 100076 1204 100082 1216
rect 110690 1204 110696 1216
rect 100076 1176 110696 1204
rect 100076 1164 100082 1176
rect 110690 1164 110696 1176
rect 110748 1164 110754 1216
rect 110782 1164 110788 1216
rect 110840 1204 110846 1216
rect 112806 1204 112812 1216
rect 110840 1176 112812 1204
rect 110840 1164 110846 1176
rect 112806 1164 112812 1176
rect 112864 1164 112870 1216
rect 113082 1164 113088 1216
rect 113140 1204 113146 1216
rect 113140 1176 113772 1204
rect 113140 1164 113146 1176
rect 93302 1096 93308 1148
rect 93360 1136 93366 1148
rect 108850 1136 108856 1148
rect 93360 1108 108856 1136
rect 93360 1096 93366 1108
rect 108850 1096 108856 1108
rect 108908 1096 108914 1148
rect 108942 1096 108948 1148
rect 109000 1136 109006 1148
rect 113634 1136 113640 1148
rect 109000 1108 113640 1136
rect 109000 1096 109006 1108
rect 113634 1096 113640 1108
rect 113692 1096 113698 1148
rect 113744 1136 113772 1176
rect 113818 1164 113824 1216
rect 113876 1204 113882 1216
rect 115014 1204 115020 1216
rect 113876 1176 115020 1204
rect 113876 1164 113882 1176
rect 115014 1164 115020 1176
rect 115072 1164 115078 1216
rect 115106 1164 115112 1216
rect 115164 1204 115170 1216
rect 123496 1204 123524 1244
rect 126882 1232 126888 1244
rect 126940 1232 126946 1284
rect 126974 1232 126980 1284
rect 127032 1272 127038 1284
rect 133138 1272 133144 1284
rect 127032 1244 133144 1272
rect 127032 1232 127038 1244
rect 133138 1232 133144 1244
rect 133196 1232 133202 1284
rect 133230 1232 133236 1284
rect 133288 1272 133294 1284
rect 141418 1272 141424 1284
rect 133288 1244 137876 1272
rect 133288 1232 133294 1244
rect 115164 1176 123524 1204
rect 115164 1164 115170 1176
rect 123570 1164 123576 1216
rect 123628 1204 123634 1216
rect 126146 1204 126152 1216
rect 123628 1176 126152 1204
rect 123628 1164 123634 1176
rect 126146 1164 126152 1176
rect 126204 1164 126210 1216
rect 126238 1164 126244 1216
rect 126296 1204 126302 1216
rect 137738 1204 137744 1216
rect 126296 1176 137744 1204
rect 126296 1164 126302 1176
rect 137738 1164 137744 1176
rect 137796 1164 137802 1216
rect 137848 1204 137876 1244
rect 137986 1244 141424 1272
rect 137986 1204 138014 1244
rect 141418 1232 141424 1244
rect 141476 1232 141482 1284
rect 141510 1232 141516 1284
rect 141568 1272 141574 1284
rect 146478 1272 146484 1284
rect 141568 1244 146484 1272
rect 141568 1232 141574 1244
rect 146478 1232 146484 1244
rect 146536 1232 146542 1284
rect 147766 1232 147772 1284
rect 147824 1272 147830 1284
rect 151262 1272 151268 1284
rect 147824 1244 151268 1272
rect 147824 1232 147830 1244
rect 151262 1232 151268 1244
rect 151320 1232 151326 1284
rect 157150 1272 157156 1284
rect 151464 1244 157156 1272
rect 137848 1176 138014 1204
rect 139302 1164 139308 1216
rect 139360 1204 139366 1216
rect 147858 1204 147864 1216
rect 139360 1176 147864 1204
rect 139360 1164 139366 1176
rect 147858 1164 147864 1176
rect 147916 1164 147922 1216
rect 148134 1164 148140 1216
rect 148192 1204 148198 1216
rect 151354 1204 151360 1216
rect 148192 1176 151360 1204
rect 148192 1164 148198 1176
rect 151354 1164 151360 1176
rect 151412 1164 151418 1216
rect 113744 1108 114968 1136
rect 87932 1040 89944 1068
rect 87932 1028 87938 1040
rect 92198 1028 92204 1080
rect 92256 1068 92262 1080
rect 94314 1068 94320 1080
rect 92256 1040 94320 1068
rect 92256 1028 92262 1040
rect 94314 1028 94320 1040
rect 94372 1028 94378 1080
rect 94682 1028 94688 1080
rect 94740 1068 94746 1080
rect 102502 1068 102508 1080
rect 94740 1040 99604 1068
rect 94740 1028 94746 1040
rect 90174 1000 90180 1012
rect 87064 972 90180 1000
rect 90174 960 90180 972
rect 90232 960 90238 1012
rect 90266 960 90272 1012
rect 90324 1000 90330 1012
rect 94130 1000 94136 1012
rect 90324 972 94136 1000
rect 90324 960 90330 972
rect 94130 960 94136 972
rect 94188 960 94194 1012
rect 99374 1000 99380 1012
rect 94516 972 99380 1000
rect 91278 932 91284 944
rect 76616 836 80468 864
rect 81360 836 82584 864
rect 83568 904 91284 932
rect 76616 824 76622 836
rect 76234 768 76512 796
rect 77322 796 77378 800
rect 78030 796 78036 808
rect 77322 768 78036 796
rect 76234 0 76290 768
rect 77322 0 77378 768
rect 78030 756 78036 768
rect 78088 756 78094 808
rect 78410 796 78466 800
rect 79134 796 79140 808
rect 78410 768 79140 796
rect 78410 0 78466 768
rect 79134 756 79140 768
rect 79192 756 79198 808
rect 79498 796 79554 800
rect 80238 796 80244 808
rect 79498 768 80244 796
rect 79498 0 79554 768
rect 80238 756 80244 768
rect 80296 756 80302 808
rect 80586 796 80642 800
rect 81360 796 81388 836
rect 80586 768 81388 796
rect 81674 796 81730 800
rect 82446 796 82452 808
rect 81674 768 82452 796
rect 80586 0 80642 768
rect 81674 0 81730 768
rect 82446 756 82452 768
rect 82504 756 82510 808
rect 82762 728 82818 800
rect 83568 728 83596 904
rect 91278 892 91284 904
rect 91336 892 91342 944
rect 91370 892 91376 944
rect 91428 932 91434 944
rect 94314 932 94320 944
rect 91428 904 94320 932
rect 91428 892 91434 904
rect 94314 892 94320 904
rect 94372 892 94378 944
rect 84010 824 84016 876
rect 84068 864 84074 876
rect 86908 864 86914 876
rect 84068 836 86914 864
rect 84068 824 84074 836
rect 86908 824 86914 836
rect 86966 824 86972 876
rect 91830 864 91836 876
rect 87984 836 91836 864
rect 82762 700 83596 728
rect 83850 728 83906 800
rect 84938 796 84994 800
rect 85758 796 85764 808
rect 84938 768 85764 796
rect 84654 728 84660 740
rect 83850 700 84660 728
rect 82762 0 82818 700
rect 83850 0 83906 700
rect 84654 688 84660 700
rect 84712 688 84718 740
rect 84938 0 84994 768
rect 85758 756 85764 768
rect 85816 756 85822 808
rect 86026 592 86082 800
rect 87114 796 87170 800
rect 87874 796 87880 808
rect 87114 768 87880 796
rect 86862 592 86868 604
rect 86026 564 86868 592
rect 86026 0 86082 564
rect 86862 552 86868 564
rect 86920 552 86926 604
rect 87114 0 87170 768
rect 87874 756 87880 768
rect 87932 756 87938 808
rect 87230 688 87236 740
rect 87288 728 87294 740
rect 87984 728 88012 836
rect 91830 824 91836 836
rect 91888 824 91894 876
rect 87288 700 88012 728
rect 87288 688 87294 700
rect 88202 524 88258 800
rect 89290 796 89346 800
rect 90082 796 90088 808
rect 89290 768 90088 796
rect 89162 524 89168 536
rect 88202 496 89168 524
rect 88202 0 88258 496
rect 89162 484 89168 496
rect 89220 484 89226 536
rect 89290 0 89346 768
rect 90082 756 90088 768
rect 90140 756 90146 808
rect 90378 796 90434 800
rect 91370 796 91376 808
rect 90378 768 91376 796
rect 90378 0 90434 768
rect 91370 756 91376 768
rect 91428 756 91434 808
rect 91466 796 91522 800
rect 92198 796 92204 808
rect 91466 768 92204 796
rect 91466 0 91522 768
rect 92198 756 92204 768
rect 92256 756 92262 808
rect 92554 796 92610 800
rect 93302 796 93308 808
rect 92554 768 93308 796
rect 92554 0 92610 768
rect 93302 756 93308 768
rect 93360 756 93366 808
rect 93642 796 93698 800
rect 94516 796 94544 972
rect 99374 960 99380 972
rect 99432 960 99438 1012
rect 99576 1000 99604 1040
rect 99944 1040 102508 1068
rect 99944 1000 99972 1040
rect 102502 1028 102508 1040
rect 102560 1028 102566 1080
rect 104158 1028 104164 1080
rect 104216 1068 104222 1080
rect 110782 1068 110788 1080
rect 104216 1040 110788 1068
rect 104216 1028 104222 1040
rect 110782 1028 110788 1040
rect 110840 1028 110846 1080
rect 110874 1028 110880 1080
rect 110932 1068 110938 1080
rect 113818 1068 113824 1080
rect 110932 1040 113824 1068
rect 110932 1028 110938 1040
rect 113818 1028 113824 1040
rect 113876 1028 113882 1080
rect 113910 1028 113916 1080
rect 113968 1068 113974 1080
rect 114554 1068 114560 1080
rect 113968 1040 114560 1068
rect 113968 1028 113974 1040
rect 114554 1028 114560 1040
rect 114612 1028 114618 1080
rect 99576 972 99972 1000
rect 100938 960 100944 1012
rect 100996 1000 101002 1012
rect 113358 1000 113364 1012
rect 100996 972 113364 1000
rect 100996 960 101002 972
rect 113358 960 113364 972
rect 113416 960 113422 1012
rect 114940 1000 114968 1108
rect 115198 1096 115204 1148
rect 115256 1136 115262 1148
rect 121730 1136 121736 1148
rect 115256 1108 121736 1136
rect 115256 1096 115262 1108
rect 121730 1096 121736 1108
rect 121788 1096 121794 1148
rect 122098 1096 122104 1148
rect 122156 1136 122162 1148
rect 130746 1136 130752 1148
rect 122156 1108 130752 1136
rect 122156 1096 122162 1108
rect 130746 1096 130752 1108
rect 130804 1096 130810 1148
rect 132954 1096 132960 1148
rect 133012 1136 133018 1148
rect 139210 1136 139216 1148
rect 133012 1108 139216 1136
rect 133012 1096 133018 1108
rect 139210 1096 139216 1108
rect 139268 1096 139274 1148
rect 139394 1096 139400 1148
rect 139452 1136 139458 1148
rect 146386 1136 146392 1148
rect 139452 1108 146392 1136
rect 139452 1096 139458 1108
rect 146386 1096 146392 1108
rect 146444 1096 146450 1148
rect 148042 1096 148048 1148
rect 148100 1136 148106 1148
rect 150342 1136 150348 1148
rect 148100 1108 150348 1136
rect 148100 1096 148106 1108
rect 150342 1096 150348 1108
rect 150400 1096 150406 1148
rect 150434 1096 150440 1148
rect 150492 1136 150498 1148
rect 151464 1136 151492 1244
rect 157150 1232 157156 1244
rect 157208 1232 157214 1284
rect 157242 1232 157248 1284
rect 157300 1272 157306 1284
rect 183508 1272 183514 1284
rect 157300 1244 183514 1272
rect 157300 1232 157306 1244
rect 183508 1232 183514 1244
rect 183566 1232 183572 1284
rect 183824 1272 183852 1300
rect 186130 1272 186136 1284
rect 183824 1244 186136 1272
rect 186130 1232 186136 1244
rect 186188 1232 186194 1284
rect 186406 1232 186412 1284
rect 186464 1272 186470 1284
rect 244090 1272 244096 1284
rect 186464 1244 244096 1272
rect 186464 1232 186470 1244
rect 244090 1232 244096 1244
rect 244148 1232 244154 1284
rect 244366 1232 244372 1284
rect 244424 1272 244430 1284
rect 246684 1272 246712 1312
rect 244424 1244 246712 1272
rect 244424 1232 244430 1244
rect 247586 1232 247592 1284
rect 247644 1272 247650 1284
rect 254412 1272 254440 1312
rect 258074 1300 258080 1312
rect 258132 1300 258138 1352
rect 258902 1300 258908 1352
rect 258960 1340 258966 1352
rect 263410 1340 263416 1352
rect 258960 1312 263416 1340
rect 258960 1300 258966 1312
rect 263410 1300 263416 1312
rect 263468 1300 263474 1352
rect 263520 1340 263548 1380
rect 267826 1368 267832 1420
rect 267884 1408 267890 1420
rect 269850 1408 269856 1420
rect 267884 1380 269856 1408
rect 267884 1368 267890 1380
rect 269850 1368 269856 1380
rect 269908 1368 269914 1420
rect 274266 1368 274272 1420
rect 274324 1408 274330 1420
rect 282638 1408 282644 1420
rect 274324 1380 282644 1408
rect 274324 1368 274330 1380
rect 282638 1368 282644 1380
rect 282696 1368 282702 1420
rect 282840 1380 282960 1408
rect 282840 1340 282868 1380
rect 263520 1312 282868 1340
rect 282932 1340 282960 1380
rect 283190 1368 283196 1420
rect 283248 1408 283254 1420
rect 289906 1408 289912 1420
rect 283248 1380 289912 1408
rect 283248 1368 283254 1380
rect 289906 1368 289912 1380
rect 289964 1368 289970 1420
rect 295794 1368 295800 1420
rect 295852 1408 295858 1420
rect 298186 1408 298192 1420
rect 295852 1380 298192 1408
rect 295852 1368 295858 1380
rect 298186 1368 298192 1380
rect 298244 1368 298250 1420
rect 300210 1368 300216 1420
rect 300268 1408 300274 1420
rect 303522 1408 303528 1420
rect 300268 1380 303528 1408
rect 300268 1368 300274 1380
rect 303522 1368 303528 1380
rect 303580 1368 303586 1420
rect 306558 1368 306564 1420
rect 306616 1408 306622 1420
rect 318702 1408 318708 1420
rect 306616 1380 318708 1408
rect 306616 1368 306622 1380
rect 318702 1368 318708 1380
rect 318760 1368 318766 1420
rect 332318 1368 332324 1420
rect 332376 1408 332382 1420
rect 375558 1408 375564 1420
rect 332376 1380 375564 1408
rect 332376 1368 332382 1380
rect 375558 1368 375564 1380
rect 375616 1368 375622 1420
rect 386414 1368 386420 1420
rect 386472 1408 386478 1420
rect 426986 1408 426992 1420
rect 386472 1380 426992 1408
rect 386472 1368 386478 1380
rect 426986 1368 426992 1380
rect 427044 1368 427050 1420
rect 360194 1340 360200 1352
rect 282932 1312 360200 1340
rect 360194 1300 360200 1312
rect 360252 1300 360258 1352
rect 372706 1340 372712 1352
rect 369826 1312 372712 1340
rect 255406 1272 255412 1284
rect 247644 1244 254440 1272
rect 254504 1244 255412 1272
rect 247644 1232 247650 1244
rect 151538 1164 151544 1216
rect 151596 1204 151602 1216
rect 156874 1204 156880 1216
rect 151596 1176 156880 1204
rect 151596 1164 151602 1176
rect 156874 1164 156880 1176
rect 156932 1164 156938 1216
rect 156966 1164 156972 1216
rect 157024 1204 157030 1216
rect 166994 1204 167000 1216
rect 157024 1176 167000 1204
rect 157024 1164 157030 1176
rect 166994 1164 167000 1176
rect 167052 1164 167058 1216
rect 167086 1164 167092 1216
rect 167144 1204 167150 1216
rect 176378 1204 176384 1216
rect 167144 1176 176384 1204
rect 167144 1164 167150 1176
rect 176378 1164 176384 1176
rect 176436 1164 176442 1216
rect 176562 1164 176568 1216
rect 176620 1204 176626 1216
rect 176620 1176 181576 1204
rect 176620 1164 176626 1176
rect 150492 1108 151492 1136
rect 150492 1096 150498 1108
rect 152366 1096 152372 1148
rect 152424 1136 152430 1148
rect 156782 1136 156788 1148
rect 152424 1108 156788 1136
rect 152424 1096 152430 1108
rect 156782 1096 156788 1108
rect 156840 1096 156846 1148
rect 158898 1096 158904 1148
rect 158956 1136 158962 1148
rect 166718 1136 166724 1148
rect 158956 1108 166724 1136
rect 158956 1096 158962 1108
rect 166718 1096 166724 1108
rect 166776 1096 166782 1148
rect 166810 1096 166816 1148
rect 166868 1136 166874 1148
rect 167178 1136 167184 1148
rect 166868 1108 167184 1136
rect 166868 1096 166874 1108
rect 167178 1096 167184 1108
rect 167236 1096 167242 1148
rect 168098 1096 168104 1148
rect 168156 1136 168162 1148
rect 170858 1136 170864 1148
rect 168156 1108 170864 1136
rect 168156 1096 168162 1108
rect 170858 1096 170864 1108
rect 170916 1096 170922 1148
rect 170950 1096 170956 1148
rect 171008 1136 171014 1148
rect 173250 1136 173256 1148
rect 171008 1108 173256 1136
rect 171008 1096 171014 1108
rect 173250 1096 173256 1108
rect 173308 1096 173314 1148
rect 173342 1096 173348 1148
rect 173400 1136 173406 1148
rect 181548 1136 181576 1176
rect 181622 1164 181628 1216
rect 181680 1204 181686 1216
rect 183646 1204 183652 1216
rect 181680 1176 183652 1204
rect 181680 1164 181686 1176
rect 183646 1164 183652 1176
rect 183704 1164 183710 1216
rect 183830 1164 183836 1216
rect 183888 1204 183894 1216
rect 183888 1176 186084 1204
rect 183888 1164 183894 1176
rect 183922 1136 183928 1148
rect 173400 1108 181484 1136
rect 181548 1108 183928 1136
rect 173400 1096 173406 1108
rect 115014 1028 115020 1080
rect 115072 1068 115078 1080
rect 118602 1068 118608 1080
rect 115072 1040 118608 1068
rect 115072 1028 115078 1040
rect 118602 1028 118608 1040
rect 118660 1028 118666 1080
rect 118786 1028 118792 1080
rect 118844 1068 118850 1080
rect 142706 1068 142712 1080
rect 118844 1040 142712 1068
rect 118844 1028 118850 1040
rect 142706 1028 142712 1040
rect 142764 1028 142770 1080
rect 156690 1068 156696 1080
rect 142816 1040 156696 1068
rect 115198 1000 115204 1012
rect 114940 972 115204 1000
rect 115198 960 115204 972
rect 115256 960 115262 1012
rect 116486 960 116492 1012
rect 116544 1000 116550 1012
rect 133046 1000 133052 1012
rect 116544 972 128492 1000
rect 116544 960 116550 972
rect 94590 892 94596 944
rect 94648 932 94654 944
rect 97534 932 97540 944
rect 94648 904 97540 932
rect 94648 892 94654 904
rect 97534 892 97540 904
rect 97592 892 97598 944
rect 113910 932 113916 944
rect 103532 904 113916 932
rect 97442 864 97448 876
rect 96586 836 97448 864
rect 93642 768 94544 796
rect 94730 796 94786 800
rect 95510 796 95516 808
rect 94730 768 95516 796
rect 93642 0 93698 768
rect 94730 0 94786 768
rect 95510 756 95516 768
rect 95568 756 95574 808
rect 95818 796 95874 800
rect 96586 796 96614 836
rect 97442 824 97448 836
rect 97500 824 97506 876
rect 103532 864 103560 904
rect 113910 892 113916 904
rect 113968 892 113974 944
rect 114002 892 114008 944
rect 114060 932 114066 944
rect 128262 932 128268 944
rect 114060 904 128268 932
rect 114060 892 114066 904
rect 128262 892 128268 904
rect 128320 892 128326 944
rect 128464 932 128492 972
rect 130672 972 133052 1000
rect 128464 904 128860 932
rect 103348 836 103560 864
rect 95818 768 96614 796
rect 95818 0 95874 768
rect 96906 456 96962 800
rect 97994 796 98050 800
rect 98822 796 98828 808
rect 97994 768 98828 796
rect 97902 456 97908 468
rect 96906 428 97908 456
rect 96906 0 96962 428
rect 97902 416 97908 428
rect 97960 416 97966 468
rect 97994 0 98050 768
rect 98822 756 98828 768
rect 98880 756 98886 808
rect 99082 796 99138 800
rect 99742 796 99748 808
rect 99082 768 99748 796
rect 99082 0 99138 768
rect 99742 756 99748 768
rect 99800 756 99806 808
rect 100170 728 100226 800
rect 101258 796 101314 800
rect 102042 796 102048 808
rect 101258 768 102048 796
rect 100938 728 100944 740
rect 100170 700 100944 728
rect 100170 0 100226 700
rect 100938 688 100944 700
rect 100996 688 101002 740
rect 101258 0 101314 768
rect 102042 756 102048 768
rect 102100 756 102106 808
rect 102346 796 102402 800
rect 103348 796 103376 836
rect 103606 824 103612 876
rect 103664 864 103670 876
rect 108298 864 108304 876
rect 103664 836 108304 864
rect 103664 824 103670 836
rect 108298 824 108304 836
rect 108356 824 108362 876
rect 119614 864 119620 876
rect 108408 836 113864 864
rect 102346 768 103376 796
rect 103434 796 103490 800
rect 104158 796 104164 808
rect 103434 768 104164 796
rect 102346 0 102402 768
rect 103434 0 103490 768
rect 104158 756 104164 768
rect 104216 756 104222 808
rect 104522 796 104578 800
rect 105262 796 105268 808
rect 104522 768 105268 796
rect 104522 0 104578 768
rect 105262 756 105268 768
rect 105320 756 105326 808
rect 105610 796 105666 800
rect 106550 796 106556 808
rect 105610 768 106556 796
rect 105610 0 105666 768
rect 106550 756 106556 768
rect 106608 756 106614 808
rect 106698 796 106754 800
rect 107470 796 107476 808
rect 106698 768 107476 796
rect 106698 0 106754 768
rect 107470 756 107476 768
rect 107528 756 107534 808
rect 107786 796 107842 800
rect 108408 796 108436 836
rect 107786 768 108436 796
rect 107786 0 107842 768
rect 108758 756 108764 808
rect 108816 796 108822 808
rect 108874 796 108930 800
rect 108816 768 108930 796
rect 108816 756 108822 768
rect 108874 0 108930 768
rect 109962 796 110018 800
rect 110874 796 110880 808
rect 109962 768 110880 796
rect 109962 0 110018 768
rect 110874 756 110880 768
rect 110932 756 110938 808
rect 111050 796 111106 800
rect 111886 796 111892 808
rect 111050 768 111892 796
rect 111050 0 111106 768
rect 111886 756 111892 768
rect 111944 756 111950 808
rect 112138 796 112194 800
rect 113082 796 113088 808
rect 112138 768 113088 796
rect 112138 0 112194 768
rect 113082 756 113088 768
rect 113140 756 113146 808
rect 113226 660 113282 800
rect 113836 728 113864 836
rect 114112 836 119620 864
rect 114112 728 114140 836
rect 119614 824 119620 836
rect 119672 824 119678 876
rect 123570 864 123576 876
rect 119724 836 123576 864
rect 113836 700 114140 728
rect 114314 796 114370 800
rect 116486 796 116492 808
rect 114314 768 116492 796
rect 114002 660 114008 672
rect 113226 632 114008 660
rect 113226 0 113282 632
rect 114002 620 114008 632
rect 114060 620 114066 672
rect 113358 552 113364 604
rect 113416 592 113422 604
rect 114186 592 114192 604
rect 113416 564 114192 592
rect 113416 552 113422 564
rect 114186 552 114192 564
rect 114244 552 114250 604
rect 114314 0 114370 768
rect 116486 756 116492 768
rect 116544 756 116550 808
rect 114738 688 114744 740
rect 114796 728 114802 740
rect 119724 728 119752 836
rect 123570 824 123576 836
rect 123628 824 123634 876
rect 127986 864 127992 876
rect 124048 836 127992 864
rect 114796 700 119752 728
rect 120026 796 120082 800
rect 122098 796 122104 808
rect 120026 768 122104 796
rect 114796 688 114802 700
rect 115382 620 115388 672
rect 115440 660 115446 672
rect 118510 660 118516 672
rect 115440 632 118516 660
rect 115440 620 115446 632
rect 118510 620 118516 632
rect 118568 620 118574 672
rect 118602 620 118608 672
rect 118660 660 118666 672
rect 119522 660 119528 672
rect 118660 632 119528 660
rect 118660 620 118666 632
rect 119522 620 119528 632
rect 119580 620 119586 672
rect 114462 552 114468 604
rect 114520 592 114526 604
rect 119706 592 119712 604
rect 114520 564 119712 592
rect 114520 552 114526 564
rect 119706 552 119712 564
rect 119764 552 119770 604
rect 114922 484 114928 536
rect 114980 524 114986 536
rect 118602 524 118608 536
rect 114980 496 118608 524
rect 114980 484 114986 496
rect 118602 484 118608 496
rect 118660 484 118666 536
rect 114738 416 114744 468
rect 114796 456 114802 468
rect 117498 456 117504 468
rect 114796 428 117504 456
rect 114796 416 114802 428
rect 117498 416 117504 428
rect 117556 416 117562 468
rect 114554 212 114560 264
rect 114612 252 114618 264
rect 119430 252 119436 264
rect 114612 224 119436 252
rect 114612 212 114618 224
rect 119430 212 119436 224
rect 119488 212 119494 264
rect 120026 0 120082 768
rect 122098 756 122104 768
rect 122156 756 122162 808
rect 122202 728 122258 800
rect 124048 728 124076 836
rect 127986 824 127992 836
rect 128044 824 128050 876
rect 128832 864 128860 904
rect 130470 864 130476 876
rect 128832 836 130476 864
rect 130470 824 130476 836
rect 130528 824 130534 876
rect 122202 700 124076 728
rect 124378 796 124434 800
rect 126238 796 126244 808
rect 124378 768 126244 796
rect 122202 0 122258 700
rect 124378 0 124434 768
rect 126238 756 126244 768
rect 126296 756 126302 808
rect 126554 796 126610 800
rect 128170 796 128176 808
rect 126554 768 128176 796
rect 124490 212 124496 264
rect 124548 252 124554 264
rect 126422 252 126428 264
rect 124548 224 126428 252
rect 124548 212 124554 224
rect 126422 212 126428 224
rect 126480 212 126486 264
rect 126554 0 126610 768
rect 128170 756 128176 768
rect 128228 756 128234 808
rect 128730 796 128786 800
rect 130672 796 130700 972
rect 133046 960 133052 972
rect 133104 960 133110 1012
rect 133138 960 133144 1012
rect 133196 1000 133202 1012
rect 133196 972 133368 1000
rect 133196 960 133202 972
rect 131022 892 131028 944
rect 131080 932 131086 944
rect 133340 932 133368 972
rect 134886 960 134892 1012
rect 134944 1000 134950 1012
rect 139302 1000 139308 1012
rect 134944 972 139308 1000
rect 134944 960 134950 972
rect 139302 960 139308 972
rect 139360 960 139366 1012
rect 142816 1000 142844 1040
rect 156690 1028 156696 1040
rect 156748 1028 156754 1080
rect 157518 1028 157524 1080
rect 157576 1068 157582 1080
rect 172238 1068 172244 1080
rect 157576 1040 171272 1068
rect 157576 1028 157582 1040
rect 139412 972 142844 1000
rect 139412 932 139440 972
rect 142890 960 142896 1012
rect 142948 1000 142954 1012
rect 156966 1000 156972 1012
rect 142948 972 156972 1000
rect 142948 960 142954 972
rect 156966 960 156972 972
rect 157024 960 157030 1012
rect 157334 1000 157340 1012
rect 157260 972 157340 1000
rect 131080 904 133276 932
rect 133340 904 139440 932
rect 131080 892 131086 904
rect 133248 864 133276 904
rect 139486 892 139492 944
rect 139544 932 139550 944
rect 146202 932 146208 944
rect 139544 904 146208 932
rect 139544 892 139550 904
rect 146202 892 146208 904
rect 146260 892 146266 944
rect 146478 892 146484 944
rect 146536 932 146542 944
rect 148042 932 148048 944
rect 146536 904 148048 932
rect 146536 892 146542 904
rect 148042 892 148048 904
rect 148100 892 148106 944
rect 150434 932 150440 944
rect 148152 904 150440 932
rect 137002 864 137008 876
rect 133248 836 137008 864
rect 137002 824 137008 836
rect 137060 824 137066 876
rect 137112 836 137784 864
rect 128730 768 130700 796
rect 130906 796 130962 800
rect 132954 796 132960 808
rect 130906 768 132960 796
rect 126882 620 126888 672
rect 126940 660 126946 672
rect 128354 660 128360 672
rect 126940 632 128360 660
rect 126940 620 126946 632
rect 128354 620 128360 632
rect 128412 620 128418 672
rect 128730 0 128786 768
rect 130906 0 130962 768
rect 132954 756 132960 768
rect 133012 756 133018 808
rect 133082 796 133138 800
rect 134886 796 134892 808
rect 133082 768 134892 796
rect 133082 0 133138 768
rect 134886 756 134892 768
rect 134944 756 134950 808
rect 135258 796 135314 800
rect 137112 796 137140 836
rect 135258 768 137140 796
rect 135258 0 135314 768
rect 137434 592 137490 800
rect 137756 728 137784 836
rect 137830 824 137836 876
rect 137888 864 137894 876
rect 139118 864 139124 876
rect 137888 836 139124 864
rect 137888 824 137894 836
rect 139118 824 139124 836
rect 139176 824 139182 876
rect 139210 824 139216 876
rect 139268 864 139274 876
rect 143718 864 143724 876
rect 139268 836 143724 864
rect 139268 824 139274 836
rect 143718 824 143724 836
rect 143776 824 143782 876
rect 146294 864 146300 876
rect 143828 836 146300 864
rect 139610 796 139666 800
rect 141510 796 141516 808
rect 139610 768 141516 796
rect 139394 728 139400 740
rect 137756 700 139400 728
rect 139394 688 139400 700
rect 139452 688 139458 740
rect 139302 592 139308 604
rect 137434 564 139308 592
rect 137434 0 137490 564
rect 139302 552 139308 564
rect 139360 552 139366 604
rect 139610 0 139666 768
rect 141510 756 141516 768
rect 141568 756 141574 808
rect 141786 796 141842 800
rect 143828 796 143856 836
rect 146294 824 146300 836
rect 146352 824 146358 876
rect 141786 768 143856 796
rect 141786 0 141842 768
rect 143962 660 144018 800
rect 146138 796 146194 800
rect 148152 796 148180 904
rect 150434 892 150440 904
rect 150492 892 150498 944
rect 150526 892 150532 944
rect 150584 932 150590 944
rect 154574 932 154580 944
rect 150584 904 154580 932
rect 150584 892 150590 904
rect 154574 892 154580 904
rect 154632 892 154638 944
rect 157260 932 157288 972
rect 157334 960 157340 972
rect 157392 960 157398 1012
rect 157426 960 157432 1012
rect 157484 1000 157490 1012
rect 157484 972 167040 1000
rect 157484 960 157490 972
rect 154776 904 157288 932
rect 159008 904 166672 932
rect 150360 836 154574 864
rect 146138 768 148180 796
rect 148314 796 148370 800
rect 150360 796 150388 836
rect 154546 808 154574 836
rect 148314 768 150388 796
rect 145834 660 145840 672
rect 143962 632 145840 660
rect 143962 0 144018 632
rect 145834 620 145840 632
rect 145892 620 145898 672
rect 146138 0 146194 768
rect 146386 8 146392 60
rect 146444 48 146450 60
rect 147950 48 147956 60
rect 146444 20 147956 48
rect 146444 8 146450 20
rect 147950 8 147956 20
rect 148008 8 148014 60
rect 148314 0 148370 768
rect 150490 728 150546 800
rect 152366 728 152372 740
rect 150490 700 152372 728
rect 150490 0 150546 700
rect 152366 688 152372 700
rect 152424 688 152430 740
rect 152666 660 152722 800
rect 154546 768 154580 808
rect 154574 756 154580 768
rect 154632 756 154638 808
rect 154776 660 154804 904
rect 159008 864 159036 904
rect 156800 836 159036 864
rect 152666 632 154804 660
rect 154842 796 154898 800
rect 156800 796 156828 836
rect 159082 824 159088 876
rect 159140 864 159146 876
rect 159140 836 166580 864
rect 159140 824 159146 836
rect 154842 768 156828 796
rect 152666 0 152722 632
rect 154842 0 154898 768
rect 157018 456 157074 800
rect 159194 728 159250 800
rect 161370 796 161426 800
rect 161750 796 161756 808
rect 161370 768 161756 796
rect 161198 728 161204 740
rect 159194 700 161204 728
rect 157150 552 157156 604
rect 157208 592 157214 604
rect 158990 592 158996 604
rect 157208 564 158996 592
rect 157208 552 157214 564
rect 158990 552 158996 564
rect 159048 552 159054 604
rect 157242 484 157248 536
rect 157300 524 157306 536
rect 158898 524 158904 536
rect 157300 496 158904 524
rect 157300 484 157306 496
rect 158898 484 158904 496
rect 158956 484 158962 536
rect 158990 456 158996 468
rect 157018 428 158996 456
rect 157018 0 157074 428
rect 158990 416 158996 428
rect 159048 416 159054 468
rect 159194 0 159250 700
rect 161198 688 161204 700
rect 161256 688 161262 740
rect 161370 0 161426 768
rect 161750 756 161756 768
rect 161808 756 161814 808
rect 162050 728 162106 800
rect 162050 700 162854 728
rect 162050 0 162106 700
rect 162826 660 162854 700
rect 164050 660 164056 672
rect 162826 632 164056 660
rect 164050 620 164056 632
rect 164108 620 164114 672
rect 164226 524 164282 800
rect 164326 620 164332 672
rect 164384 660 164390 672
rect 166258 660 166264 672
rect 164384 632 166264 660
rect 164384 620 164390 632
rect 166258 620 166264 632
rect 166316 620 166322 672
rect 166258 524 166264 536
rect 164226 496 166264 524
rect 164226 0 164282 496
rect 166258 484 166264 496
rect 166316 484 166322 536
rect 166402 388 166458 800
rect 166552 592 166580 836
rect 166644 796 166672 904
rect 167012 864 167040 972
rect 167178 960 167184 1012
rect 167236 1000 167242 1012
rect 171134 1000 171140 1012
rect 167236 972 171140 1000
rect 167236 960 167242 972
rect 171134 960 171140 972
rect 171192 960 171198 1012
rect 171244 1000 171272 1040
rect 171888 1040 172244 1068
rect 171888 1000 171916 1040
rect 172238 1028 172244 1040
rect 172296 1028 172302 1080
rect 172330 1028 172336 1080
rect 172388 1068 172394 1080
rect 176470 1068 176476 1080
rect 172388 1040 176476 1068
rect 172388 1028 172394 1040
rect 176470 1028 176476 1040
rect 176528 1028 176534 1080
rect 176746 1028 176752 1080
rect 176804 1068 176810 1080
rect 181346 1068 181352 1080
rect 176804 1040 181352 1068
rect 176804 1028 176810 1040
rect 181346 1028 181352 1040
rect 181404 1028 181410 1080
rect 181456 1068 181484 1108
rect 183922 1096 183928 1108
rect 183980 1096 183986 1148
rect 184014 1096 184020 1148
rect 184072 1136 184078 1148
rect 185854 1136 185860 1148
rect 184072 1108 185860 1136
rect 184072 1096 184078 1108
rect 185854 1096 185860 1108
rect 185912 1096 185918 1148
rect 181456 1040 183876 1068
rect 177482 1000 177488 1012
rect 171244 972 171916 1000
rect 171980 972 177488 1000
rect 168098 892 168104 944
rect 168156 932 168162 944
rect 170950 932 170956 944
rect 168156 904 170956 932
rect 168156 892 168162 904
rect 170950 892 170956 904
rect 171008 892 171014 944
rect 168282 864 168288 876
rect 167012 836 168288 864
rect 168282 824 168288 836
rect 168340 824 168346 876
rect 171980 864 172008 972
rect 177482 960 177488 972
rect 177540 960 177546 1012
rect 183508 1000 183514 1012
rect 177592 972 183514 1000
rect 172238 892 172244 944
rect 172296 932 172302 944
rect 176930 932 176936 944
rect 172296 904 176936 932
rect 172296 892 172302 904
rect 176930 892 176936 904
rect 176988 892 176994 944
rect 177592 864 177620 972
rect 183508 960 183514 972
rect 183566 960 183572 1012
rect 183848 1000 183876 1040
rect 184106 1028 184112 1080
rect 184164 1068 184170 1080
rect 185946 1068 185952 1080
rect 184164 1040 185952 1068
rect 184164 1028 184170 1040
rect 185946 1028 185952 1040
rect 186004 1028 186010 1080
rect 186056 1068 186084 1176
rect 186222 1164 186228 1216
rect 186280 1204 186286 1216
rect 213086 1204 213092 1216
rect 186280 1176 213092 1204
rect 186280 1164 186286 1176
rect 213086 1164 213092 1176
rect 213144 1164 213150 1216
rect 224310 1164 224316 1216
rect 224368 1204 224374 1216
rect 224368 1176 224954 1204
rect 224368 1164 224374 1176
rect 186774 1096 186780 1148
rect 186832 1136 186838 1148
rect 195054 1136 195060 1148
rect 186832 1108 195060 1136
rect 186832 1096 186838 1108
rect 195054 1096 195060 1108
rect 195112 1096 195118 1148
rect 215386 1136 215392 1148
rect 195164 1108 215392 1136
rect 186682 1068 186688 1080
rect 186056 1040 186688 1068
rect 186682 1028 186688 1040
rect 186740 1028 186746 1080
rect 186866 1028 186872 1080
rect 186924 1068 186930 1080
rect 195164 1068 195192 1108
rect 215386 1096 215392 1108
rect 215444 1096 215450 1148
rect 219710 1096 219716 1148
rect 219768 1136 219774 1148
rect 223390 1136 223396 1148
rect 219768 1108 223396 1136
rect 219768 1096 219774 1108
rect 223390 1096 223396 1108
rect 223448 1096 223454 1148
rect 224926 1136 224954 1176
rect 226426 1164 226432 1216
rect 226484 1204 226490 1216
rect 236270 1204 236276 1216
rect 226484 1176 236276 1204
rect 226484 1164 226490 1176
rect 236270 1164 236276 1176
rect 236328 1164 236334 1216
rect 238478 1164 238484 1216
rect 238536 1204 238542 1216
rect 243906 1204 243912 1216
rect 238536 1176 243912 1204
rect 238536 1164 238542 1176
rect 243906 1164 243912 1176
rect 243964 1164 243970 1216
rect 244642 1164 244648 1216
rect 244700 1204 244706 1216
rect 254504 1204 254532 1244
rect 255406 1232 255412 1244
rect 255464 1232 255470 1284
rect 256878 1232 256884 1284
rect 256936 1272 256942 1284
rect 267826 1272 267832 1284
rect 256936 1244 267832 1272
rect 256936 1232 256942 1244
rect 267826 1232 267832 1244
rect 267884 1232 267890 1284
rect 267918 1232 267924 1284
rect 267976 1272 267982 1284
rect 282822 1272 282828 1284
rect 267976 1244 282828 1272
rect 267976 1232 267982 1244
rect 282822 1232 282828 1244
rect 282880 1232 282886 1284
rect 283006 1232 283012 1284
rect 283064 1272 283070 1284
rect 369826 1272 369854 1312
rect 372706 1300 372712 1312
rect 372764 1300 372770 1352
rect 460382 1340 460388 1352
rect 376726 1312 379514 1340
rect 376726 1272 376754 1312
rect 283064 1244 369854 1272
rect 371896 1244 376754 1272
rect 283064 1232 283070 1244
rect 244700 1176 254532 1204
rect 244700 1164 244706 1176
rect 254762 1164 254768 1216
rect 254820 1204 254826 1216
rect 268010 1204 268016 1216
rect 254820 1176 268016 1204
rect 254820 1164 254826 1176
rect 268010 1164 268016 1176
rect 268068 1164 268074 1216
rect 268654 1164 268660 1216
rect 268712 1204 268718 1216
rect 273254 1204 273260 1216
rect 268712 1176 273260 1204
rect 268712 1164 268718 1176
rect 273254 1164 273260 1176
rect 273312 1164 273318 1216
rect 273346 1164 273352 1216
rect 273404 1204 273410 1216
rect 276014 1204 276020 1216
rect 273404 1176 276020 1204
rect 273404 1164 273410 1176
rect 276014 1164 276020 1176
rect 276072 1164 276078 1216
rect 278038 1164 278044 1216
rect 278096 1204 278102 1216
rect 282546 1204 282552 1216
rect 278096 1176 282552 1204
rect 278096 1164 278102 1176
rect 282546 1164 282552 1176
rect 282604 1164 282610 1216
rect 371896 1204 371924 1244
rect 287164 1176 371924 1204
rect 379486 1204 379514 1312
rect 457824 1312 460388 1340
rect 448514 1272 448520 1284
rect 446784 1244 448520 1272
rect 383010 1204 383016 1216
rect 379486 1176 383016 1204
rect 224926 1108 229232 1136
rect 186924 1040 195192 1068
rect 186924 1028 186930 1040
rect 195238 1028 195244 1080
rect 195296 1068 195302 1080
rect 220538 1068 220544 1080
rect 195296 1040 220544 1068
rect 195296 1028 195302 1040
rect 220538 1028 220544 1040
rect 220596 1028 220602 1080
rect 222102 1028 222108 1080
rect 222160 1068 222166 1080
rect 229094 1068 229100 1080
rect 222160 1040 229100 1068
rect 222160 1028 222166 1040
rect 229094 1028 229100 1040
rect 229152 1028 229158 1080
rect 229204 1068 229232 1108
rect 230566 1096 230572 1148
rect 230624 1136 230630 1148
rect 230624 1108 234614 1136
rect 230624 1096 230630 1108
rect 233694 1068 233700 1080
rect 229204 1040 233700 1068
rect 233694 1028 233700 1040
rect 233752 1028 233758 1080
rect 234586 1068 234614 1108
rect 237282 1096 237288 1148
rect 237340 1136 237346 1148
rect 237340 1108 244504 1136
rect 237340 1096 237346 1108
rect 241422 1068 241428 1080
rect 234586 1040 241428 1068
rect 241422 1028 241428 1040
rect 241480 1028 241486 1080
rect 241514 1028 241520 1080
rect 241572 1068 241578 1080
rect 242894 1068 242900 1080
rect 241572 1040 242900 1068
rect 241572 1028 241578 1040
rect 242894 1028 242900 1040
rect 242952 1028 242958 1080
rect 242986 1028 242992 1080
rect 243044 1068 243050 1080
rect 244366 1068 244372 1080
rect 243044 1040 244372 1068
rect 243044 1028 243050 1040
rect 244366 1028 244372 1040
rect 244424 1028 244430 1080
rect 244476 1068 244504 1108
rect 245746 1096 245752 1148
rect 245804 1136 245810 1148
rect 253842 1136 253848 1148
rect 245804 1108 253848 1136
rect 245804 1096 245810 1108
rect 253842 1096 253848 1108
rect 253900 1096 253906 1148
rect 253934 1096 253940 1148
rect 253992 1136 253998 1148
rect 267182 1136 267188 1148
rect 253992 1108 267188 1136
rect 253992 1096 253998 1108
rect 267182 1096 267188 1108
rect 267240 1096 267246 1148
rect 267734 1096 267740 1148
rect 267792 1136 267798 1148
rect 282730 1136 282736 1148
rect 267792 1108 282736 1136
rect 267792 1096 267798 1108
rect 282730 1096 282736 1108
rect 282788 1096 282794 1148
rect 247034 1068 247040 1080
rect 244476 1040 247040 1068
rect 247034 1028 247040 1040
rect 247092 1028 247098 1080
rect 248046 1028 248052 1080
rect 248104 1068 248110 1080
rect 254946 1068 254952 1080
rect 248104 1040 254952 1068
rect 248104 1028 248110 1040
rect 254946 1028 254952 1040
rect 255004 1028 255010 1080
rect 255038 1028 255044 1080
rect 255096 1068 255102 1080
rect 261202 1068 261208 1080
rect 255096 1040 261208 1068
rect 255096 1028 255102 1040
rect 261202 1028 261208 1040
rect 261260 1028 261266 1080
rect 261294 1028 261300 1080
rect 261352 1068 261358 1080
rect 271598 1068 271604 1080
rect 261352 1040 271604 1068
rect 261352 1028 261358 1040
rect 271598 1028 271604 1040
rect 271656 1028 271662 1080
rect 271690 1028 271696 1080
rect 271748 1068 271754 1080
rect 282454 1068 282460 1080
rect 271748 1040 282460 1068
rect 271748 1028 271754 1040
rect 282454 1028 282460 1040
rect 282512 1028 282518 1080
rect 283098 1028 283104 1080
rect 283156 1068 283162 1080
rect 287164 1068 287192 1176
rect 383010 1164 383016 1176
rect 383068 1164 383074 1216
rect 287238 1096 287244 1148
rect 287296 1136 287302 1148
rect 292206 1136 292212 1148
rect 287296 1108 292212 1136
rect 287296 1096 287302 1108
rect 292206 1096 292212 1108
rect 292264 1096 292270 1148
rect 292298 1096 292304 1148
rect 292356 1136 292362 1148
rect 293494 1136 293500 1148
rect 292356 1108 293500 1136
rect 292356 1096 292362 1108
rect 293494 1096 293500 1108
rect 293552 1096 293558 1148
rect 302510 1136 302516 1148
rect 297376 1108 302516 1136
rect 283156 1040 287192 1068
rect 283156 1028 283162 1040
rect 287790 1028 287796 1080
rect 287848 1068 287854 1080
rect 291010 1068 291016 1080
rect 287848 1040 291016 1068
rect 287848 1028 287854 1040
rect 291010 1028 291016 1040
rect 291068 1028 291074 1080
rect 291102 1028 291108 1080
rect 291160 1068 291166 1080
rect 297376 1068 297404 1108
rect 302510 1096 302516 1108
rect 302568 1096 302574 1148
rect 304810 1096 304816 1148
rect 304868 1136 304874 1148
rect 311894 1136 311900 1148
rect 304868 1108 311900 1136
rect 304868 1096 304874 1108
rect 311894 1096 311900 1108
rect 311952 1096 311958 1148
rect 311986 1096 311992 1148
rect 312044 1136 312050 1148
rect 336734 1136 336740 1148
rect 312044 1108 336740 1136
rect 312044 1096 312050 1108
rect 336734 1096 336740 1108
rect 336792 1096 336798 1148
rect 365070 1096 365076 1148
rect 365128 1136 365134 1148
rect 365128 1108 373166 1136
rect 365128 1096 365134 1108
rect 302694 1068 302700 1080
rect 291160 1040 297404 1068
rect 297468 1040 302700 1068
rect 291160 1028 291166 1040
rect 183848 972 187004 1000
rect 177942 892 177948 944
rect 178000 932 178006 944
rect 181530 932 181536 944
rect 178000 904 181536 932
rect 178000 892 178006 904
rect 181530 892 181536 904
rect 181588 892 181594 944
rect 183646 932 183652 944
rect 181732 904 183652 932
rect 168392 836 172008 864
rect 172256 836 177620 864
rect 168190 796 168196 808
rect 166644 768 168196 796
rect 168190 756 168196 768
rect 168248 756 168254 808
rect 166718 688 166724 740
rect 166776 728 166782 740
rect 168282 728 168288 740
rect 166776 700 168288 728
rect 166776 688 166782 700
rect 168282 688 168288 700
rect 168340 688 168346 740
rect 166626 620 166632 672
rect 166684 660 166690 672
rect 168392 660 168420 836
rect 166684 632 168420 660
rect 166684 620 166690 632
rect 168466 592 168472 604
rect 166552 564 168472 592
rect 168466 552 168472 564
rect 168524 552 168530 604
rect 166534 484 166540 536
rect 166592 524 166598 536
rect 168098 524 168104 536
rect 166592 496 168104 524
rect 166592 484 166598 496
rect 168098 484 168104 496
rect 168156 484 168162 536
rect 168578 524 168634 800
rect 170754 728 170810 800
rect 171042 756 171048 808
rect 171100 796 171106 808
rect 172256 796 172284 836
rect 177666 824 177672 876
rect 177724 864 177730 876
rect 178678 864 178684 876
rect 177724 836 178684 864
rect 177724 824 177730 836
rect 178678 824 178684 836
rect 178736 824 178742 876
rect 181732 864 181760 904
rect 183646 892 183652 904
rect 183704 892 183710 944
rect 185670 892 185676 944
rect 185728 932 185734 944
rect 186866 932 186872 944
rect 185728 904 186872 932
rect 185728 892 185734 904
rect 186866 892 186872 904
rect 186924 892 186930 944
rect 186976 932 187004 972
rect 187878 960 187884 1012
rect 187936 1000 187942 1012
rect 218238 1000 218244 1012
rect 187936 972 218244 1000
rect 187936 960 187942 972
rect 218238 960 218244 972
rect 218296 960 218302 1012
rect 228542 1000 228548 1012
rect 219406 972 228548 1000
rect 186976 904 194916 932
rect 179340 836 181760 864
rect 171100 768 172284 796
rect 172930 796 172986 800
rect 173342 796 173348 808
rect 172930 768 173348 796
rect 171100 756 171106 768
rect 172330 728 172336 740
rect 170754 700 172336 728
rect 170398 524 170404 536
rect 168578 496 170404 524
rect 166902 388 166908 400
rect 166402 360 166908 388
rect 166402 0 166458 360
rect 166902 348 166908 360
rect 166960 348 166966 400
rect 168578 0 168634 496
rect 170398 484 170404 496
rect 170456 484 170462 536
rect 170754 0 170810 700
rect 172330 688 172336 700
rect 172388 688 172394 740
rect 170858 620 170864 672
rect 170916 660 170922 672
rect 172790 660 172796 672
rect 170916 632 172796 660
rect 170916 620 170922 632
rect 172790 620 172796 632
rect 172848 620 172854 672
rect 172930 0 172986 768
rect 173342 756 173348 768
rect 173400 756 173406 808
rect 175106 796 175162 800
rect 177022 796 177028 808
rect 175106 768 177028 796
rect 173158 688 173164 740
rect 173216 728 173222 740
rect 174998 728 175004 740
rect 173216 700 175004 728
rect 173216 688 173222 700
rect 174998 688 175004 700
rect 175056 688 175062 740
rect 173066 552 173072 604
rect 173124 592 173130 604
rect 173986 592 173992 604
rect 173124 564 173992 592
rect 173124 552 173130 564
rect 173986 552 173992 564
rect 174044 552 174050 604
rect 173250 8 173256 60
rect 173308 48 173314 60
rect 174814 48 174820 60
rect 173308 20 174820 48
rect 173308 8 173314 20
rect 174814 8 174820 20
rect 174872 8 174878 60
rect 175106 0 175162 768
rect 177022 756 177028 768
rect 177080 756 177086 808
rect 177282 796 177338 800
rect 179340 796 179368 836
rect 183922 824 183928 876
rect 183980 864 183986 876
rect 194888 864 194916 904
rect 198734 892 198740 944
rect 198792 932 198798 944
rect 219406 932 219434 972
rect 228542 960 228548 972
rect 228600 960 228606 1012
rect 231670 960 231676 1012
rect 231728 1000 231734 1012
rect 231728 972 239260 1000
rect 231728 960 231734 972
rect 198792 904 219434 932
rect 198792 892 198798 904
rect 219526 892 219532 944
rect 219584 932 219590 944
rect 239122 932 239128 944
rect 219584 904 239128 932
rect 219584 892 219590 904
rect 239122 892 239128 904
rect 239180 892 239186 944
rect 239232 932 239260 972
rect 239398 960 239404 1012
rect 239456 1000 239462 1012
rect 262398 1000 262404 1012
rect 239456 972 262404 1000
rect 239456 960 239462 972
rect 262398 960 262404 972
rect 262456 960 262462 1012
rect 262490 960 262496 1012
rect 262548 1000 262554 1012
rect 274082 1000 274088 1012
rect 262548 972 263548 1000
rect 262548 960 262554 972
rect 239950 932 239956 944
rect 239232 904 239956 932
rect 239950 892 239956 904
rect 240008 892 240014 944
rect 241606 932 241612 944
rect 240060 904 241612 932
rect 195238 864 195244 876
rect 183980 836 194824 864
rect 194888 836 195244 864
rect 183980 824 183986 836
rect 177282 768 179368 796
rect 177282 0 177338 768
rect 179458 592 179514 800
rect 181634 796 181690 800
rect 183508 796 183514 808
rect 181634 768 183514 796
rect 181254 592 181260 604
rect 179458 564 181260 592
rect 179458 0 179514 564
rect 181254 552 181260 564
rect 181312 552 181318 604
rect 179782 144 179788 196
rect 179840 184 179846 196
rect 181254 184 181260 196
rect 179840 156 181260 184
rect 179840 144 179846 156
rect 181254 144 181260 156
rect 181312 144 181318 196
rect 181634 0 181690 768
rect 183508 756 183514 768
rect 183566 756 183572 808
rect 183810 796 183866 800
rect 185670 796 185676 808
rect 183810 768 185676 796
rect 181898 552 181904 604
rect 181956 592 181962 604
rect 183554 592 183560 604
rect 181956 564 183560 592
rect 181956 552 181962 564
rect 183554 552 183560 564
rect 183612 552 183618 604
rect 181898 144 181904 196
rect 181956 184 181962 196
rect 183646 184 183652 196
rect 181956 156 183652 184
rect 181956 144 181962 156
rect 183646 144 183652 156
rect 183704 144 183710 196
rect 183810 0 183866 768
rect 185670 756 185676 768
rect 185728 756 185734 808
rect 185986 728 186042 800
rect 188162 796 188218 800
rect 190178 796 190184 808
rect 188162 768 190184 796
rect 187878 728 187884 740
rect 185986 700 187884 728
rect 185986 0 186042 700
rect 187878 688 187884 700
rect 187936 688 187942 740
rect 188162 0 188218 768
rect 190178 756 190184 768
rect 190236 756 190242 808
rect 190338 320 190394 800
rect 192514 660 192570 800
rect 194594 660 194600 672
rect 192514 632 194600 660
rect 192202 320 192208 332
rect 190338 292 192208 320
rect 190338 0 190394 292
rect 192202 280 192208 292
rect 192260 280 192266 332
rect 192514 0 192570 632
rect 194594 620 194600 632
rect 194652 620 194658 672
rect 192846 484 192852 536
rect 192904 524 192910 536
rect 194318 524 194324 536
rect 192904 496 194324 524
rect 192904 484 192910 496
rect 194318 484 194324 496
rect 194376 484 194382 536
rect 194690 388 194746 800
rect 194796 796 194824 836
rect 195238 824 195244 836
rect 195296 824 195302 876
rect 197998 824 198004 876
rect 198056 864 198062 876
rect 219618 864 219624 876
rect 198056 836 219624 864
rect 198056 824 198062 836
rect 219618 824 219624 836
rect 219676 824 219682 876
rect 240060 864 240088 904
rect 241606 892 241612 904
rect 241664 892 241670 944
rect 241698 892 241704 944
rect 241756 932 241762 944
rect 245746 932 245752 944
rect 241756 904 245752 932
rect 241756 892 241762 904
rect 245746 892 245752 904
rect 245804 892 245810 944
rect 246022 892 246028 944
rect 246080 932 246086 944
rect 247586 932 247592 944
rect 246080 904 247592 932
rect 246080 892 246086 904
rect 247586 892 247592 904
rect 247644 892 247650 944
rect 247696 904 250560 932
rect 219912 836 240088 864
rect 194962 796 194968 808
rect 194796 768 194968 796
rect 194962 756 194968 768
rect 195020 756 195026 808
rect 196342 756 196348 808
rect 196400 796 196406 808
rect 212074 796 212080 808
rect 196400 768 212080 796
rect 196400 756 196406 768
rect 212074 756 212080 768
rect 212132 756 212138 808
rect 219912 728 219940 836
rect 241974 824 241980 876
rect 242032 864 242038 876
rect 247696 864 247724 904
rect 242032 836 247724 864
rect 250532 864 250560 904
rect 250806 892 250812 944
rect 250864 932 250870 944
rect 253750 932 253756 944
rect 250864 904 253756 932
rect 250864 892 250870 904
rect 253750 892 253756 904
rect 253808 892 253814 944
rect 263520 932 263548 972
rect 265360 972 274088 1000
rect 265360 932 265388 972
rect 274082 960 274088 972
rect 274140 960 274146 1012
rect 276474 960 276480 1012
rect 276532 1000 276538 1012
rect 282362 1000 282368 1012
rect 276532 972 282368 1000
rect 276532 960 276538 972
rect 282362 960 282368 972
rect 282420 960 282426 1012
rect 282822 960 282828 1012
rect 282880 1000 282886 1012
rect 282880 972 293816 1000
rect 282880 960 282886 972
rect 254044 904 263456 932
rect 263520 904 265388 932
rect 254044 864 254072 904
rect 250532 836 254072 864
rect 242032 824 242038 836
rect 254118 824 254124 876
rect 254176 864 254182 876
rect 263428 864 263456 904
rect 265434 892 265440 944
rect 265492 932 265498 944
rect 267826 932 267832 944
rect 265492 904 267832 932
rect 265492 892 265498 904
rect 267826 892 267832 904
rect 267884 892 267890 944
rect 273162 932 273168 944
rect 267936 904 273168 932
rect 265618 864 265624 876
rect 254176 836 262628 864
rect 263428 836 265624 864
rect 254176 824 254182 836
rect 200086 700 219940 728
rect 220054 796 220110 800
rect 222102 796 222108 808
rect 220054 768 222108 796
rect 195146 620 195152 672
rect 195204 660 195210 672
rect 200086 660 200114 700
rect 219526 660 219532 672
rect 195204 632 200114 660
rect 209746 632 219532 660
rect 195204 620 195210 632
rect 194962 552 194968 604
rect 195020 592 195026 604
rect 195974 592 195980 604
rect 195020 564 195980 592
rect 195020 552 195026 564
rect 195974 552 195980 564
rect 196032 552 196038 604
rect 196066 552 196072 604
rect 196124 592 196130 604
rect 209746 592 209774 632
rect 219526 620 219532 632
rect 219584 620 219590 672
rect 196124 564 209774 592
rect 196124 552 196130 564
rect 195054 484 195060 536
rect 195112 524 195118 536
rect 196342 524 196348 536
rect 195112 496 196348 524
rect 195112 484 195118 496
rect 196342 484 196348 496
rect 196400 484 196406 536
rect 194870 416 194876 468
rect 194928 456 194934 468
rect 197998 456 198004 468
rect 194928 428 198004 456
rect 194928 416 194934 428
rect 197998 416 198004 428
rect 198056 416 198062 468
rect 198734 388 198740 400
rect 194690 360 198740 388
rect 192938 76 192944 128
rect 192996 116 193002 128
rect 194594 116 194600 128
rect 192996 88 194600 116
rect 192996 76 193002 88
rect 194594 76 194600 88
rect 194652 76 194658 128
rect 192846 8 192852 60
rect 192904 48 192910 60
rect 194502 48 194508 60
rect 192904 20 194508 48
rect 192904 8 192910 20
rect 194502 8 194508 20
rect 194560 8 194566 60
rect 194690 0 194746 360
rect 198734 348 198740 360
rect 198792 348 198798 400
rect 195238 280 195244 332
rect 195296 320 195302 332
rect 202782 320 202788 332
rect 195296 292 202788 320
rect 195296 280 195302 292
rect 202782 280 202788 292
rect 202840 280 202846 332
rect 194962 212 194968 264
rect 195020 252 195026 264
rect 210234 252 210240 264
rect 195020 224 210240 252
rect 195020 212 195026 224
rect 210234 212 210240 224
rect 210292 212 210298 264
rect 195974 144 195980 196
rect 196032 184 196038 196
rect 207934 184 207940 196
rect 196032 156 207940 184
rect 196032 144 196038 156
rect 207934 144 207940 156
rect 207992 144 207998 196
rect 194778 76 194784 128
rect 194836 116 194842 128
rect 205082 116 205088 128
rect 194836 88 205088 116
rect 194836 76 194842 88
rect 205082 76 205088 88
rect 205140 76 205146 128
rect 194870 8 194876 60
rect 194928 48 194934 60
rect 219710 48 219716 60
rect 194928 20 219716 48
rect 194928 8 194934 20
rect 219710 8 219716 20
rect 219768 8 219774 60
rect 220054 0 220110 768
rect 222102 756 222108 768
rect 222160 756 222166 808
rect 222230 796 222286 800
rect 224310 796 224316 808
rect 222230 768 224316 796
rect 222230 0 222286 768
rect 224310 756 224316 768
rect 224368 756 224374 808
rect 224406 796 224462 800
rect 226426 796 226432 808
rect 224406 768 226432 796
rect 224406 0 224462 768
rect 226426 756 226432 768
rect 226484 756 226490 808
rect 226582 796 226638 800
rect 228450 796 228456 808
rect 226582 768 228456 796
rect 226582 0 226638 768
rect 228450 756 228456 768
rect 228508 756 228514 808
rect 228758 796 228814 800
rect 230566 796 230572 808
rect 228758 768 230572 796
rect 228758 0 228814 768
rect 230566 756 230572 768
rect 230624 756 230630 808
rect 230934 796 230990 800
rect 231670 796 231676 808
rect 230934 768 231676 796
rect 230934 0 230990 768
rect 231670 756 231676 768
rect 231728 756 231734 808
rect 233110 796 233166 800
rect 234982 796 234988 808
rect 233110 768 234988 796
rect 233110 0 233166 768
rect 234982 756 234988 768
rect 235040 756 235046 808
rect 235286 796 235342 800
rect 237282 796 237288 808
rect 235286 768 237288 796
rect 235286 0 235342 768
rect 237282 756 237288 768
rect 237340 756 237346 808
rect 237462 796 237518 800
rect 238478 796 238484 808
rect 237462 768 238484 796
rect 237462 0 237518 768
rect 238478 756 238484 768
rect 238536 756 238542 808
rect 239638 796 239694 800
rect 241698 796 241704 808
rect 239638 768 241704 796
rect 239638 0 239694 768
rect 241698 756 241704 768
rect 241756 756 241762 808
rect 241814 796 241870 800
rect 242986 796 242992 808
rect 241814 768 242992 796
rect 239950 688 239956 740
rect 240008 728 240014 740
rect 241514 728 241520 740
rect 240008 700 241520 728
rect 240008 688 240014 700
rect 241514 688 241520 700
rect 241572 688 241578 740
rect 241814 0 241870 768
rect 242986 756 242992 768
rect 243044 756 243050 808
rect 243990 660 244046 800
rect 246166 796 246222 800
rect 248046 796 248052 808
rect 246166 768 248052 796
rect 246022 660 246028 672
rect 243990 632 246028 660
rect 243990 0 244046 632
rect 246022 620 246028 632
rect 246080 620 246086 672
rect 246166 0 246222 768
rect 248046 756 248052 768
rect 248104 756 248110 808
rect 248342 184 248398 800
rect 250518 660 250574 800
rect 250806 660 250812 672
rect 250518 632 250812 660
rect 250346 184 250352 196
rect 248342 156 250352 184
rect 248342 0 248398 156
rect 250346 144 250352 156
rect 250404 144 250410 196
rect 250518 0 250574 632
rect 250806 620 250812 632
rect 250864 620 250870 672
rect 252694 660 252750 800
rect 254870 796 254926 800
rect 256878 796 256884 808
rect 254870 768 256884 796
rect 254762 660 254768 672
rect 252694 632 254768 660
rect 250622 212 250628 264
rect 250680 252 250686 264
rect 252554 252 252560 264
rect 250680 224 252560 252
rect 250680 212 250686 224
rect 252554 212 252560 224
rect 252612 212 252618 264
rect 252694 0 252750 632
rect 254762 620 254768 632
rect 254820 620 254826 672
rect 254870 0 254926 768
rect 256878 756 256884 768
rect 256936 756 256942 808
rect 257046 796 257102 800
rect 258902 796 258908 808
rect 257046 768 258908 796
rect 257046 0 257102 768
rect 258902 756 258908 768
rect 258960 756 258966 808
rect 259222 796 259278 800
rect 261294 796 261300 808
rect 259222 768 261300 796
rect 259222 0 259278 768
rect 261294 756 261300 768
rect 261352 756 261358 808
rect 261398 796 261454 800
rect 262490 796 262496 808
rect 261398 768 262496 796
rect 259362 416 259368 468
rect 259420 456 259426 468
rect 260834 456 260840 468
rect 259420 428 260840 456
rect 259420 416 259426 428
rect 260834 416 260840 428
rect 260892 416 260898 468
rect 261398 0 261454 768
rect 262490 756 262496 768
rect 262548 756 262554 808
rect 262600 796 262628 836
rect 265618 824 265624 836
rect 265676 824 265682 876
rect 265894 824 265900 876
rect 265952 864 265958 876
rect 267936 864 267964 904
rect 273162 892 273168 904
rect 273220 892 273226 944
rect 273346 892 273352 944
rect 273404 932 273410 944
rect 278038 932 278044 944
rect 273404 904 274404 932
rect 273404 892 273410 904
rect 265952 836 267964 864
rect 265952 824 265958 836
rect 268194 824 268200 876
rect 268252 864 268258 876
rect 274266 864 274272 876
rect 268252 836 274272 864
rect 268252 824 268258 836
rect 274266 824 274272 836
rect 274324 824 274330 876
rect 274376 864 274404 904
rect 274652 904 278044 932
rect 274652 864 274680 904
rect 278038 892 278044 904
rect 278096 892 278102 944
rect 278590 932 278596 944
rect 278148 904 278596 932
rect 274376 836 274680 864
rect 274818 824 274824 876
rect 274876 864 274882 876
rect 278148 864 278176 904
rect 278590 892 278596 904
rect 278648 892 278654 944
rect 278682 892 278688 944
rect 278740 932 278746 944
rect 278740 904 280568 932
rect 278740 892 278746 904
rect 274876 836 278176 864
rect 274876 824 274882 836
rect 278958 824 278964 876
rect 279016 864 279022 876
rect 280338 864 280344 876
rect 279016 836 280344 864
rect 279016 824 279022 836
rect 280338 824 280344 836
rect 280396 824 280402 876
rect 280540 864 280568 904
rect 280890 892 280896 944
rect 280948 932 280954 944
rect 283006 932 283012 944
rect 280948 904 283012 932
rect 280948 892 280954 904
rect 283006 892 283012 904
rect 283064 892 283070 944
rect 283190 892 283196 944
rect 283248 932 283254 944
rect 283248 904 289676 932
rect 283248 892 283254 904
rect 282914 864 282920 876
rect 280540 836 282920 864
rect 282914 824 282920 836
rect 282972 824 282978 876
rect 287790 864 287796 876
rect 285048 836 287796 864
rect 263410 796 263416 808
rect 262600 768 263416 796
rect 263410 756 263416 768
rect 263468 756 263474 808
rect 263574 660 263630 800
rect 265750 728 265806 800
rect 267734 728 267740 740
rect 265750 700 267740 728
rect 265434 660 265440 672
rect 263574 632 265440 660
rect 263574 0 263630 632
rect 265434 620 265440 632
rect 265492 620 265498 672
rect 265750 0 265806 700
rect 267734 688 267740 700
rect 267792 688 267798 740
rect 267926 728 267982 800
rect 270102 796 270158 800
rect 271690 796 271696 808
rect 270102 768 271696 796
rect 268654 728 268660 740
rect 267926 700 268660 728
rect 267926 0 267982 700
rect 268654 688 268660 700
rect 268712 688 268718 740
rect 270102 0 270158 768
rect 271690 756 271696 768
rect 271748 756 271754 808
rect 272278 728 272334 800
rect 274454 796 274510 800
rect 276474 796 276480 808
rect 274454 768 276480 796
rect 273990 728 273996 740
rect 272278 700 273996 728
rect 272278 0 272334 700
rect 273990 688 273996 700
rect 274048 688 274054 740
rect 274454 0 274510 768
rect 276474 756 276480 768
rect 276532 756 276538 808
rect 276630 796 276686 800
rect 278590 796 278596 808
rect 276630 768 278596 796
rect 276630 0 276686 768
rect 278590 756 278596 768
rect 278648 756 278654 808
rect 278806 592 278862 800
rect 280982 796 281038 800
rect 282822 796 282828 808
rect 280982 768 282828 796
rect 280890 592 280896 604
rect 278806 564 280896 592
rect 278806 0 278862 564
rect 280890 552 280896 564
rect 280948 552 280954 604
rect 280982 0 281038 768
rect 282822 756 282828 768
rect 282880 756 282886 808
rect 283158 728 283214 800
rect 285048 796 285076 836
rect 287790 824 287796 836
rect 287848 824 287854 876
rect 289538 864 289544 876
rect 289372 836 289544 864
rect 284956 768 285076 796
rect 285334 796 285390 800
rect 287238 796 287244 808
rect 285334 768 287244 796
rect 284956 728 284984 768
rect 283158 700 284984 728
rect 283158 0 283214 700
rect 285334 0 285390 768
rect 287238 756 287244 768
rect 287296 756 287302 808
rect 287510 796 287566 800
rect 289372 796 289400 836
rect 289538 824 289544 836
rect 289596 824 289602 876
rect 289648 864 289676 904
rect 289722 892 289728 944
rect 289780 932 289786 944
rect 293788 932 293816 972
rect 293862 960 293868 1012
rect 293920 1000 293926 1012
rect 297468 1000 297496 1040
rect 302694 1028 302700 1040
rect 302752 1028 302758 1080
rect 306926 1028 306932 1080
rect 306984 1068 306990 1080
rect 334158 1068 334164 1080
rect 306984 1040 315436 1068
rect 306984 1028 306990 1040
rect 293920 972 297496 1000
rect 293920 960 293926 972
rect 297542 960 297548 1012
rect 297600 1000 297606 1012
rect 300210 1000 300216 1012
rect 297600 972 300216 1000
rect 297600 960 297606 972
rect 300210 960 300216 972
rect 300268 960 300274 1012
rect 300394 960 300400 1012
rect 300452 1000 300458 1012
rect 300452 972 302556 1000
rect 300452 960 300458 972
rect 295794 932 295800 944
rect 289780 904 292160 932
rect 293788 904 295800 932
rect 289780 892 289786 904
rect 291746 864 291752 876
rect 289648 836 291752 864
rect 291746 824 291752 836
rect 291804 824 291810 876
rect 287510 768 289400 796
rect 289686 796 289742 800
rect 291102 796 291108 808
rect 289686 768 291108 796
rect 287510 0 287566 768
rect 289686 0 289742 768
rect 291102 756 291108 768
rect 291160 756 291166 808
rect 291862 524 291918 800
rect 292132 796 292160 904
rect 295794 892 295800 904
rect 295852 892 295858 944
rect 302528 932 302556 972
rect 302786 960 302792 1012
rect 302844 1000 302850 1012
rect 315298 1000 315304 1012
rect 302844 972 315304 1000
rect 302844 960 302850 972
rect 315298 960 315304 972
rect 315356 960 315362 1012
rect 315408 1000 315436 1040
rect 316788 1040 334164 1068
rect 316494 1000 316500 1012
rect 315408 972 316500 1000
rect 316494 960 316500 972
rect 316552 960 316558 1012
rect 295996 904 302464 932
rect 302528 904 306696 932
rect 293862 796 293868 808
rect 292132 768 293868 796
rect 293862 756 293868 768
rect 293920 756 293926 808
rect 294038 796 294094 800
rect 295996 796 296024 904
rect 302326 864 302332 876
rect 297836 836 302332 864
rect 294038 768 296024 796
rect 296214 796 296270 800
rect 297836 796 297864 836
rect 302326 824 302332 836
rect 302384 824 302390 876
rect 302436 864 302464 904
rect 306558 864 306564 876
rect 302436 836 306564 864
rect 306558 824 306564 836
rect 306616 824 306622 876
rect 306668 864 306696 904
rect 308122 892 308128 944
rect 308180 932 308186 944
rect 316788 932 316816 1040
rect 334158 1028 334164 1040
rect 334216 1028 334222 1080
rect 357986 1028 357992 1080
rect 358044 1068 358050 1080
rect 362586 1068 362592 1080
rect 358044 1040 362592 1068
rect 358044 1028 358050 1040
rect 362586 1028 362592 1040
rect 362644 1028 362650 1080
rect 364352 1040 367048 1068
rect 316862 960 316868 1012
rect 316920 1000 316926 1012
rect 331214 1000 331220 1012
rect 316920 972 331220 1000
rect 316920 960 316926 972
rect 331214 960 331220 972
rect 331272 960 331278 1012
rect 359918 960 359924 1012
rect 359976 1000 359982 1012
rect 364352 1000 364380 1040
rect 359976 972 364380 1000
rect 367020 1000 367048 1040
rect 367094 1028 367100 1080
rect 367152 1068 367158 1080
rect 367152 1040 370988 1068
rect 367152 1028 367158 1040
rect 367020 972 368812 1000
rect 359976 960 359982 972
rect 308180 904 316816 932
rect 308180 892 308186 904
rect 316954 892 316960 944
rect 317012 932 317018 944
rect 341886 932 341892 944
rect 317012 904 341892 932
rect 317012 892 317018 904
rect 341886 892 341892 904
rect 341944 892 341950 944
rect 357342 892 357348 944
rect 357400 932 357406 944
rect 357400 904 364104 932
rect 357400 892 357406 904
rect 307202 864 307208 876
rect 306668 836 307208 864
rect 307202 824 307208 836
rect 307260 824 307266 876
rect 307386 824 307392 876
rect 307444 864 307450 876
rect 313366 864 313372 876
rect 307444 836 313372 864
rect 307444 824 307450 836
rect 313366 824 313372 836
rect 313424 824 313430 876
rect 339310 864 339316 876
rect 313476 836 321554 864
rect 296214 768 297864 796
rect 298390 796 298446 800
rect 300394 796 300400 808
rect 298390 768 300400 796
rect 293862 524 293868 536
rect 291862 496 293868 524
rect 291862 0 291918 496
rect 293862 484 293868 496
rect 293920 484 293926 536
rect 294038 0 294094 768
rect 296214 0 296270 768
rect 298390 0 298446 768
rect 300394 756 300400 768
rect 300452 756 300458 808
rect 300566 796 300622 800
rect 302602 796 302608 808
rect 300566 768 302608 796
rect 298554 76 298560 128
rect 298612 116 298618 128
rect 300394 116 300400 128
rect 298612 88 300400 116
rect 298612 76 298618 88
rect 300394 76 300400 88
rect 300452 76 300458 128
rect 300566 0 300622 768
rect 302602 756 302608 768
rect 302660 756 302666 808
rect 302742 796 302798 800
rect 304810 796 304816 808
rect 302742 768 304816 796
rect 302742 0 302798 768
rect 304810 756 304816 768
rect 304868 756 304874 808
rect 304918 796 304974 800
rect 306926 796 306932 808
rect 304918 768 306932 796
rect 304918 0 304974 768
rect 306926 756 306932 768
rect 306984 756 306990 808
rect 307094 796 307150 800
rect 308122 796 308128 808
rect 307094 768 308128 796
rect 307094 0 307150 768
rect 308122 756 308128 768
rect 308180 756 308186 808
rect 309270 796 309326 800
rect 311066 796 311072 808
rect 309270 768 311072 796
rect 309270 0 309326 768
rect 311066 756 311072 768
rect 311124 756 311130 808
rect 311446 660 311502 800
rect 313476 660 313504 836
rect 311446 632 313504 660
rect 313622 796 313678 800
rect 315666 796 315672 808
rect 313622 768 315672 796
rect 311446 0 311502 632
rect 313622 0 313678 768
rect 315666 756 315672 768
rect 315724 756 315730 808
rect 315798 48 315854 800
rect 315942 756 315948 808
rect 316000 796 316006 808
rect 316954 796 316960 808
rect 316000 768 316960 796
rect 316000 756 316006 768
rect 316954 756 316960 768
rect 317012 756 317018 808
rect 317974 116 318030 800
rect 321526 796 321554 836
rect 325666 836 339316 864
rect 325666 796 325694 836
rect 339310 824 339316 836
rect 339368 824 339374 876
rect 359826 824 359832 876
rect 359884 864 359890 876
rect 364076 864 364104 904
rect 368784 864 368812 972
rect 370960 864 370988 1040
rect 373138 864 373166 1108
rect 376386 1096 376392 1148
rect 376444 1136 376450 1148
rect 376444 1108 379698 1136
rect 376444 1096 376450 1108
rect 373534 1028 373540 1080
rect 373592 1068 373598 1080
rect 373592 1040 377516 1068
rect 373592 1028 373598 1040
rect 377488 864 377516 1040
rect 379670 864 379698 1108
rect 442350 1068 442356 1080
rect 359884 836 360194 864
rect 364076 836 364840 864
rect 368784 836 368888 864
rect 359884 824 359890 836
rect 321526 768 325694 796
rect 355410 756 355416 808
rect 355468 796 355474 808
rect 360066 796 360122 800
rect 355468 768 360122 796
rect 360166 796 360194 836
rect 362242 796 362298 800
rect 360166 768 362298 796
rect 355468 756 355474 768
rect 318058 212 318064 264
rect 318116 252 318122 264
rect 329006 252 329012 264
rect 318116 224 329012 252
rect 318116 212 318122 224
rect 329006 212 329012 224
rect 329064 212 329070 264
rect 318242 144 318248 196
rect 318300 184 318306 196
rect 326430 184 326436 196
rect 318300 156 326436 184
rect 318300 144 318306 156
rect 326430 144 326436 156
rect 326488 144 326494 196
rect 347038 116 347044 128
rect 317974 88 347044 116
rect 317874 48 317880 60
rect 315798 20 317880 48
rect 315798 0 315854 20
rect 317874 8 317880 20
rect 317932 8 317938 60
rect 317974 0 318030 88
rect 347038 76 347044 88
rect 347096 76 347102 128
rect 318058 8 318064 60
rect 318116 48 318122 60
rect 344462 48 344468 60
rect 318116 20 344468 48
rect 318116 8 318122 20
rect 344462 8 344468 20
rect 344520 8 344526 60
rect 360066 0 360122 768
rect 362242 0 362298 768
rect 362586 756 362592 808
rect 362644 796 362650 808
rect 364418 796 364474 800
rect 362644 768 364474 796
rect 362644 756 362650 768
rect 364418 0 364474 768
rect 364812 728 364840 836
rect 366594 728 366650 800
rect 364812 700 366650 728
rect 366594 0 366650 700
rect 368770 796 368826 800
rect 368860 796 368888 836
rect 368770 768 368888 796
rect 370884 836 370988 864
rect 373000 836 373166 864
rect 377416 836 377516 864
rect 379624 836 379698 864
rect 438412 1040 442356 1068
rect 438412 864 438440 1040
rect 442350 1028 442356 1040
rect 442408 1028 442414 1080
rect 444374 932 444380 944
rect 441586 904 444380 932
rect 438412 836 438532 864
rect 370884 796 370912 836
rect 370946 796 371002 800
rect 370884 768 371002 796
rect 368770 0 368826 768
rect 370946 0 371002 768
rect 373000 660 373028 836
rect 373122 660 373178 800
rect 373442 756 373448 808
rect 373500 796 373506 808
rect 375298 796 375354 800
rect 373500 768 375354 796
rect 377416 796 377444 836
rect 379624 800 379652 836
rect 377474 796 377530 800
rect 377416 768 377530 796
rect 379624 768 379706 800
rect 373500 756 373506 768
rect 373000 632 373178 660
rect 373122 0 373178 632
rect 375298 0 375354 768
rect 377474 0 377530 768
rect 379650 0 379706 768
rect 380894 756 380900 808
rect 380952 796 380958 808
rect 381826 796 381882 800
rect 380952 768 381882 796
rect 380952 756 380958 768
rect 381826 0 381882 768
rect 383838 756 383844 808
rect 383896 796 383902 808
rect 384002 796 384058 800
rect 383896 768 384058 796
rect 383896 756 383902 768
rect 384002 0 384058 768
rect 385034 756 385040 808
rect 385092 796 385098 808
rect 386178 796 386234 800
rect 385092 768 386234 796
rect 385092 756 385098 768
rect 386178 0 386234 768
rect 387794 756 387800 808
rect 387852 796 387858 808
rect 388354 796 388410 800
rect 387852 768 388410 796
rect 387852 756 387858 768
rect 388354 0 388410 768
rect 390530 796 390586 800
rect 390646 796 390652 808
rect 390530 768 390652 796
rect 390530 0 390586 768
rect 390646 756 390652 768
rect 390704 756 390710 808
rect 391934 756 391940 808
rect 391992 796 391998 808
rect 392706 796 392762 800
rect 391992 768 392762 796
rect 391992 756 391998 768
rect 392706 0 392762 768
rect 394050 756 394056 808
rect 394108 796 394114 808
rect 394882 796 394938 800
rect 394108 768 394938 796
rect 394108 756 394114 768
rect 394882 0 394938 768
rect 395246 756 395252 808
rect 395304 796 395310 808
rect 397058 796 397114 800
rect 395304 768 397114 796
rect 395304 756 395310 768
rect 397058 0 397114 768
rect 397638 756 397644 808
rect 397696 796 397702 808
rect 399234 796 399290 800
rect 397696 768 399290 796
rect 397696 756 397702 768
rect 399234 0 399290 768
rect 400214 756 400220 808
rect 400272 796 400278 808
rect 401410 796 401466 800
rect 400272 768 401466 796
rect 400272 756 400278 768
rect 401410 0 401466 768
rect 402422 756 402428 808
rect 402480 796 402486 808
rect 403586 796 403642 800
rect 402480 768 403642 796
rect 402480 756 402486 768
rect 403586 0 403642 768
rect 405762 728 405818 800
rect 406286 756 406292 808
rect 406344 796 406350 808
rect 407938 796 407994 800
rect 406344 768 407994 796
rect 406344 756 406350 768
rect 405918 728 405924 740
rect 405762 700 405924 728
rect 405762 0 405818 700
rect 405918 688 405924 700
rect 405976 688 405982 740
rect 407938 0 407994 768
rect 408862 756 408868 808
rect 408920 796 408926 808
rect 410114 796 410170 800
rect 408920 768 410170 796
rect 408920 756 408926 768
rect 410114 0 410170 768
rect 411438 756 411444 808
rect 411496 796 411502 808
rect 412290 796 412346 800
rect 411496 768 412346 796
rect 411496 756 411502 768
rect 412290 0 412346 768
rect 414014 756 414020 808
rect 414072 796 414078 808
rect 414466 796 414522 800
rect 414072 768 414522 796
rect 414072 756 414078 768
rect 414466 0 414522 768
rect 416498 756 416504 808
rect 416556 796 416562 808
rect 416642 796 416698 800
rect 416556 768 416698 796
rect 416556 756 416562 768
rect 416642 0 416698 768
rect 418818 796 418874 800
rect 419166 796 419172 808
rect 418818 768 419172 796
rect 418818 0 418874 768
rect 419166 756 419172 768
rect 419224 756 419230 808
rect 420994 796 421050 800
rect 421742 796 421748 808
rect 420994 768 421748 796
rect 420994 0 421050 768
rect 421742 756 421748 768
rect 421800 756 421806 808
rect 423170 796 423226 800
rect 423582 796 423588 808
rect 423170 768 423588 796
rect 423170 0 423226 768
rect 423582 756 423588 768
rect 423640 756 423646 808
rect 425346 796 425402 800
rect 426066 796 426072 808
rect 425346 768 426072 796
rect 425346 0 425402 768
rect 426066 756 426072 768
rect 426124 756 426130 808
rect 427522 796 427578 800
rect 427722 796 427728 808
rect 427522 768 427728 796
rect 427522 0 427578 768
rect 427722 756 427728 768
rect 427780 756 427786 808
rect 429698 796 429754 800
rect 430482 796 430488 808
rect 429698 768 430488 796
rect 429698 0 429754 768
rect 430482 756 430488 768
rect 430540 756 430546 808
rect 431770 756 431776 808
rect 431828 796 431834 808
rect 431874 796 431930 800
rect 431828 768 431930 796
rect 431828 756 431834 768
rect 431874 0 431930 768
rect 434050 796 434106 800
rect 434622 796 434628 808
rect 434050 768 434628 796
rect 434050 0 434106 768
rect 434622 756 434628 768
rect 434680 756 434686 808
rect 436226 796 436282 800
rect 436830 796 436836 808
rect 436226 768 436836 796
rect 436226 0 436282 768
rect 436830 756 436836 768
rect 436888 756 436894 808
rect 438402 796 438458 800
rect 438504 796 438532 836
rect 438402 768 438532 796
rect 440578 796 440634 800
rect 441586 796 441614 904
rect 444374 892 444380 904
rect 444432 892 444438 944
rect 445754 864 445760 876
rect 442920 836 445760 864
rect 440578 768 441614 796
rect 442754 796 442810 800
rect 442920 796 442948 836
rect 445754 824 445760 836
rect 445812 824 445818 876
rect 442754 768 442948 796
rect 444930 796 444986 800
rect 446784 796 446812 1244
rect 448514 1232 448520 1244
rect 448572 1232 448578 1284
rect 451366 1204 451372 1216
rect 447106 1176 451372 1204
rect 447106 864 447134 1176
rect 451366 1164 451372 1176
rect 451424 1164 451430 1216
rect 457824 1204 457852 1312
rect 460382 1300 460388 1312
rect 460440 1300 460446 1352
rect 481542 1300 481548 1352
rect 481600 1340 481606 1352
rect 491294 1340 491300 1352
rect 481600 1312 491300 1340
rect 481600 1300 481606 1312
rect 491294 1300 491300 1312
rect 491352 1300 491358 1352
rect 462314 1272 462320 1284
rect 455524 1176 457852 1204
rect 457916 1244 462320 1272
rect 453390 1136 453396 1148
rect 449296 1108 453396 1136
rect 449296 864 449324 1108
rect 453390 1096 453396 1108
rect 453448 1096 453454 1148
rect 455414 864 455420 876
rect 447106 836 447180 864
rect 447152 800 447180 836
rect 444930 768 446812 796
rect 447106 768 447180 800
rect 449176 836 449324 864
rect 453500 836 455420 864
rect 438402 0 438458 768
rect 440578 0 440634 768
rect 442754 0 442810 768
rect 444930 0 444986 768
rect 447106 0 447162 768
rect 449176 728 449204 836
rect 449282 728 449338 800
rect 449176 700 449338 728
rect 449282 0 449338 700
rect 451458 796 451514 800
rect 453500 796 453528 836
rect 455414 824 455420 836
rect 455472 824 455478 876
rect 451458 768 453528 796
rect 453634 796 453690 800
rect 455524 796 455552 1176
rect 457916 1136 457944 1244
rect 462314 1232 462320 1244
rect 462372 1232 462378 1284
rect 470594 1232 470600 1284
rect 470652 1272 470658 1284
rect 473998 1272 474004 1284
rect 470652 1244 474004 1272
rect 470652 1232 470658 1244
rect 473998 1232 474004 1244
rect 474056 1232 474062 1284
rect 485958 1232 485964 1284
rect 486016 1272 486022 1284
rect 496446 1272 496452 1284
rect 486016 1244 496452 1272
rect 486016 1232 486022 1244
rect 496446 1232 496452 1244
rect 496504 1232 496510 1284
rect 499206 1272 499212 1284
rect 496556 1244 499212 1272
rect 463786 1204 463792 1216
rect 460492 1176 463792 1204
rect 460492 1136 460520 1176
rect 463786 1164 463792 1176
rect 463844 1164 463850 1216
rect 472894 1164 472900 1216
rect 472952 1204 472958 1216
rect 478506 1204 478512 1216
rect 472952 1176 478512 1204
rect 472952 1164 472958 1176
rect 478506 1164 478512 1176
rect 478564 1164 478570 1216
rect 483750 1164 483756 1216
rect 483808 1204 483814 1216
rect 493870 1204 493876 1216
rect 483808 1176 493876 1204
rect 483808 1164 483814 1176
rect 493870 1164 493876 1176
rect 493928 1164 493934 1216
rect 455824 1108 457944 1136
rect 458008 1108 460520 1136
rect 455824 864 455852 1108
rect 453634 768 455552 796
rect 455708 836 455852 864
rect 458008 864 458036 1108
rect 464246 1096 464252 1148
rect 464304 1136 464310 1148
rect 469214 1136 469220 1148
rect 464304 1108 469220 1136
rect 464304 1096 464310 1108
rect 469214 1096 469220 1108
rect 469272 1096 469278 1148
rect 476040 1108 477724 1136
rect 466454 1068 466460 1080
rect 462516 1040 466460 1068
rect 462516 1000 462544 1040
rect 466454 1028 466460 1040
rect 466512 1028 466518 1080
rect 471882 1000 471888 1012
rect 460170 972 462544 1000
rect 464540 972 471888 1000
rect 460170 864 460198 972
rect 464540 864 464568 972
rect 471882 960 471888 972
rect 471940 960 471946 1012
rect 475930 932 475936 944
rect 470796 904 475936 932
rect 470594 864 470600 876
rect 458008 836 458128 864
rect 460170 836 460244 864
rect 464540 836 464660 864
rect 455708 796 455736 836
rect 455810 796 455866 800
rect 455708 768 455866 796
rect 451458 0 451514 768
rect 453634 0 453690 768
rect 455810 0 455866 768
rect 457986 796 458042 800
rect 458100 796 458128 836
rect 460216 800 460244 836
rect 457986 768 458128 796
rect 460162 768 460244 800
rect 462338 796 462394 800
rect 464246 796 464252 808
rect 462338 768 464252 796
rect 457986 0 458042 768
rect 460162 0 460218 768
rect 462338 0 462394 768
rect 464246 756 464252 768
rect 464304 756 464310 808
rect 464514 796 464570 800
rect 464632 796 464660 836
rect 468588 836 470600 864
rect 464514 768 464660 796
rect 464514 0 464570 768
rect 466690 728 466746 800
rect 468588 728 468616 836
rect 470594 824 470600 836
rect 470652 824 470658 876
rect 466690 700 468616 728
rect 468866 796 468922 800
rect 470796 796 470824 904
rect 475930 892 475936 904
rect 475988 892 475994 944
rect 476040 864 476068 1108
rect 477696 1000 477724 1108
rect 478874 1096 478880 1148
rect 478932 1136 478938 1148
rect 488718 1136 488724 1148
rect 478932 1108 488724 1136
rect 478932 1096 478938 1108
rect 488718 1096 488724 1108
rect 488776 1096 488782 1148
rect 489886 1108 490788 1136
rect 483566 1000 483572 1012
rect 477696 972 483572 1000
rect 483566 960 483572 972
rect 483624 960 483630 1012
rect 489886 932 489914 1108
rect 490760 1068 490788 1108
rect 491110 1096 491116 1148
rect 491168 1136 491174 1148
rect 496556 1136 496584 1244
rect 499206 1232 499212 1244
rect 499264 1232 499270 1284
rect 498286 1164 498292 1216
rect 498344 1204 498350 1216
rect 510522 1204 510528 1216
rect 498344 1176 510528 1204
rect 498344 1164 498350 1176
rect 510522 1164 510528 1176
rect 510580 1164 510586 1216
rect 491168 1108 496584 1136
rect 491168 1096 491174 1108
rect 499114 1096 499120 1148
rect 499172 1136 499178 1148
rect 505094 1136 505100 1148
rect 499172 1108 505100 1136
rect 499172 1096 499178 1108
rect 505094 1096 505100 1108
rect 505152 1096 505158 1148
rect 498194 1068 498200 1080
rect 490760 1040 498200 1068
rect 498194 1028 498200 1040
rect 498252 1028 498258 1080
rect 499206 1028 499212 1080
rect 499264 1068 499270 1080
rect 502334 1068 502340 1080
rect 499264 1040 502340 1068
rect 499264 1028 499270 1040
rect 502334 1028 502340 1040
rect 502392 1028 502398 1080
rect 500310 1000 500316 1012
rect 490760 972 500316 1000
rect 490760 932 490788 972
rect 500310 960 500316 972
rect 500368 960 500374 1012
rect 499114 932 499120 944
rect 475120 836 476068 864
rect 476960 904 480254 932
rect 468866 768 470824 796
rect 471042 796 471098 800
rect 472894 796 472900 808
rect 471042 768 472900 796
rect 466690 0 466746 700
rect 468866 0 468922 768
rect 471042 0 471098 768
rect 472894 756 472900 768
rect 472952 756 472958 808
rect 473218 728 473274 800
rect 475120 728 475148 836
rect 473218 700 475148 728
rect 475394 796 475450 800
rect 476960 796 476988 904
rect 480226 864 480254 904
rect 486298 904 489914 932
rect 490392 904 490788 932
rect 492830 904 499120 932
rect 486142 864 486148 876
rect 480226 836 486148 864
rect 486142 824 486148 836
rect 486200 824 486206 876
rect 486298 864 486326 904
rect 486252 836 486326 864
rect 475394 768 476988 796
rect 477570 796 477626 800
rect 478874 796 478880 808
rect 477570 768 478880 796
rect 473218 0 473274 700
rect 475394 0 475450 768
rect 477570 0 477626 768
rect 478874 756 478880 768
rect 478932 756 478938 808
rect 479746 796 479802 800
rect 481542 796 481548 808
rect 479746 768 481548 796
rect 479746 0 479802 768
rect 481542 756 481548 768
rect 481600 756 481606 808
rect 481922 796 481978 800
rect 483750 796 483756 808
rect 481922 768 483756 796
rect 481922 0 481978 768
rect 483750 756 483756 768
rect 483808 756 483814 808
rect 484098 796 484154 800
rect 485958 796 485964 808
rect 484098 768 485964 796
rect 484098 0 484154 768
rect 485958 756 485964 768
rect 486016 756 486022 808
rect 486252 800 486280 836
rect 486252 700 486330 800
rect 486274 0 486330 700
rect 488450 796 488506 800
rect 490392 796 490420 904
rect 492830 864 492858 904
rect 499114 892 499120 904
rect 499172 892 499178 944
rect 509326 864 509332 876
rect 492784 836 492858 864
rect 497016 836 509332 864
rect 492784 800 492812 836
rect 488450 768 490420 796
rect 488450 0 488506 768
rect 490626 728 490682 800
rect 491110 728 491116 740
rect 490626 700 491116 728
rect 490626 0 490682 700
rect 491110 688 491116 700
rect 491168 688 491174 740
rect 492784 700 492858 800
rect 492802 0 492858 700
rect 494978 796 495034 800
rect 497016 796 497044 836
rect 509326 824 509332 836
rect 509384 824 509390 876
rect 494978 768 497044 796
rect 497154 796 497210 800
rect 498286 796 498292 808
rect 497154 768 498292 796
rect 494978 0 495034 768
rect 497154 0 497210 768
rect 498286 756 498292 768
rect 498344 756 498350 808
rect 499330 48 499386 800
rect 514202 48 514208 60
rect 499330 20 514208 48
rect 499330 0 499386 20
rect 514202 8 514208 20
rect 514260 8 514266 60
<< via1 >>
rect 92204 11908 92256 11960
rect 199936 11908 199988 11960
rect 100668 11840 100720 11892
rect 199200 11840 199252 11892
rect 175464 11772 175516 11824
rect 195244 11772 195296 11824
rect 107568 11704 107620 11756
rect 194968 11704 195020 11756
rect 99932 11636 99984 11688
rect 199384 11636 199436 11688
rect 184388 11568 184440 11620
rect 195612 11568 195664 11620
rect 157892 11500 157944 11552
rect 199844 11500 199896 11552
rect 97448 11432 97500 11484
rect 195520 11432 195572 11484
rect 195888 11432 195940 11484
rect 199292 11432 199344 11484
rect 195060 11364 195112 11416
rect 200396 11840 200448 11892
rect 186688 11296 186740 11348
rect 199384 11296 199436 11348
rect 92848 11228 92900 11280
rect 123116 11160 123168 11212
rect 184204 11160 184256 11212
rect 195244 11160 195296 11212
rect 198464 11160 198516 11212
rect 199936 11160 199988 11212
rect 200856 11228 200908 11280
rect 201316 11228 201368 11280
rect 201960 11228 202012 11280
rect 202512 11228 202564 11280
rect 202972 11228 203024 11280
rect 203432 11228 203484 11280
rect 203984 11160 204036 11212
rect 204536 11160 204588 11212
rect 205088 11228 205140 11280
rect 205640 11568 205692 11620
rect 206192 11228 206244 11280
rect 98460 11092 98512 11144
rect 195336 11092 195388 11144
rect 199844 11092 199896 11144
rect 207480 11228 207532 11280
rect 208124 11228 208176 11280
rect 208584 11228 208636 11280
rect 209964 11228 210016 11280
rect 104072 11024 104124 11076
rect 195244 11024 195296 11076
rect 195612 11024 195664 11076
rect 97264 10888 97316 10940
rect 195520 10956 195572 11008
rect 198556 10956 198608 11008
rect 198648 10888 198700 10940
rect 199200 11024 199252 11076
rect 205456 11024 205508 11076
rect 205548 11024 205600 11076
rect 205640 11024 205692 11076
rect 207020 11024 207072 11076
rect 207296 11092 207348 11144
rect 210056 11160 210108 11212
rect 210700 11228 210752 11280
rect 211160 11228 211212 11280
rect 211804 11228 211856 11280
rect 212908 11364 212960 11416
rect 212724 11228 212776 11280
rect 213828 11228 213880 11280
rect 213920 11228 213972 11280
rect 214380 11432 214432 11484
rect 215392 11228 215444 11280
rect 215576 11228 215628 11280
rect 199936 10956 199988 11008
rect 201316 10956 201368 11008
rect 201408 10956 201460 11008
rect 207388 11024 207440 11076
rect 213644 11092 213696 11144
rect 214012 11092 214064 11144
rect 217048 11228 217100 11280
rect 217232 11228 217284 11280
rect 217600 11228 217652 11280
rect 218336 11228 218388 11280
rect 219256 11296 219308 11348
rect 219440 11228 219492 11280
rect 219900 11160 219952 11212
rect 220360 11228 220412 11280
rect 220912 11228 220964 11280
rect 221648 11228 221700 11280
rect 222200 11228 222252 11280
rect 222476 11228 222528 11280
rect 223212 11228 223264 11280
rect 223764 11228 223816 11280
rect 216772 11092 216824 11144
rect 224960 11228 225012 11280
rect 225420 11228 225472 11280
rect 225788 11228 225840 11280
rect 226432 11228 226484 11280
rect 226984 11228 227036 11280
rect 227352 11228 227404 11280
rect 228088 11228 228140 11280
rect 228456 11228 228508 11280
rect 229192 11228 229244 11280
rect 229836 11228 229888 11280
rect 230388 11228 230440 11280
rect 230848 11228 230900 11280
rect 231400 11228 231452 11280
rect 231860 11228 231912 11280
rect 232320 11228 232372 11280
rect 233424 11228 233476 11280
rect 233608 11228 233660 11280
rect 233884 11228 233936 11280
rect 234712 11228 234764 11280
rect 234988 11228 235040 11280
rect 235724 11228 235776 11280
rect 236276 11228 236328 11280
rect 236920 11228 236972 11280
rect 237380 11228 237432 11280
rect 237932 11228 237984 11280
rect 238300 11228 238352 11280
rect 238944 11228 238996 11280
rect 239496 11228 239548 11280
rect 240140 11228 240192 11280
rect 240416 11228 240468 11280
rect 241152 11228 241204 11280
rect 241612 11228 241664 11280
rect 242900 11228 242952 11280
rect 243360 11228 243412 11280
rect 244464 11228 244516 11280
rect 245016 11228 245068 11280
rect 245384 11228 245436 11280
rect 246120 11228 246172 11280
rect 246672 11228 246724 11280
rect 246948 11228 247000 11280
rect 247684 11228 247736 11280
rect 248604 11228 248656 11280
rect 249340 11228 249392 11280
rect 249984 11228 250036 11280
rect 250260 11228 250312 11280
rect 224776 11092 224828 11144
rect 226892 11092 226944 11144
rect 211068 11024 211120 11076
rect 229284 11024 229336 11076
rect 236644 11024 236696 11076
rect 239404 11024 239456 11076
rect 251548 11228 251600 11280
rect 251916 11228 251968 11280
rect 252744 11228 252796 11280
rect 253112 11228 253164 11280
rect 254216 11296 254268 11348
rect 254032 11228 254084 11280
rect 255320 11228 255372 11280
rect 255872 11228 255924 11280
rect 256424 11228 256476 11280
rect 277124 11636 277176 11688
rect 359740 11636 359792 11688
rect 248512 11092 248564 11144
rect 251272 11092 251324 11144
rect 255688 11092 255740 11144
rect 255228 11024 255280 11076
rect 359924 11568 359976 11620
rect 258724 11500 258776 11552
rect 354404 11500 354456 11552
rect 258632 11432 258684 11484
rect 358636 11432 358688 11484
rect 258540 11364 258592 11416
rect 311256 11364 311308 11416
rect 207296 10956 207348 11008
rect 212080 10956 212132 11008
rect 212172 10956 212224 11008
rect 224776 10956 224828 11008
rect 229652 10956 229704 11008
rect 239220 10956 239272 11008
rect 254952 10956 255004 11008
rect 346768 11296 346820 11348
rect 347596 11296 347648 11348
rect 355784 11296 355836 11348
rect 102876 10820 102928 10872
rect 96068 10752 96120 10804
rect 195152 10752 195204 10804
rect 195336 10820 195388 10872
rect 201224 10820 201276 10872
rect 201500 10888 201552 10940
rect 216772 10888 216824 10940
rect 220176 10820 220228 10872
rect 221372 10820 221424 10872
rect 206928 10752 206980 10804
rect 207020 10752 207072 10804
rect 101956 10684 102008 10736
rect 205640 10684 205692 10736
rect 205732 10684 205784 10736
rect 212172 10684 212224 10736
rect 212356 10752 212408 10804
rect 225052 10752 225104 10804
rect 226892 10820 226944 10872
rect 235724 10888 235776 10940
rect 236644 10888 236696 10940
rect 248696 10888 248748 10940
rect 249064 10888 249116 10940
rect 229744 10820 229796 10872
rect 239404 10820 239456 10872
rect 238852 10752 238904 10804
rect 219440 10684 219492 10736
rect 220084 10684 220136 10736
rect 258540 10820 258592 10872
rect 248696 10752 248748 10804
rect 336280 11160 336332 11212
rect 342720 11160 342772 11212
rect 355416 11160 355468 11212
rect 360752 11228 360804 11280
rect 360936 11228 360988 11280
rect 361304 11228 361356 11280
rect 362040 11228 362092 11280
rect 362408 11228 362460 11280
rect 363144 11432 363196 11484
rect 363696 11228 363748 11280
rect 364248 11228 364300 11280
rect 258816 11092 258868 11144
rect 364524 11160 364576 11212
rect 365260 11228 365312 11280
rect 365812 11228 365864 11280
rect 366364 11228 366416 11280
rect 366732 11228 366784 11280
rect 367468 11228 367520 11280
rect 368020 11228 368072 11280
rect 368664 11228 368716 11280
rect 368940 11160 368992 11212
rect 369768 11228 369820 11280
rect 370136 11228 370188 11280
rect 370688 11228 370740 11280
rect 371056 11228 371108 11280
rect 371792 11228 371844 11280
rect 372160 11228 372212 11280
rect 372896 11228 372948 11280
rect 373264 11228 373316 11280
rect 374000 11228 374052 11280
rect 374368 11228 374420 11280
rect 375104 11228 375156 11280
rect 375472 11228 375524 11280
rect 376208 11228 376260 11280
rect 377036 11228 377088 11280
rect 377312 11228 377364 11280
rect 377588 11228 377640 11280
rect 378416 11228 378468 11280
rect 378692 11228 378744 11280
rect 379428 11228 379480 11280
rect 380348 11228 380400 11280
rect 355784 11092 355836 11144
rect 251180 10684 251232 10736
rect 255320 10684 255372 10736
rect 260840 10752 260892 10804
rect 195244 10616 195296 10668
rect 198648 10616 198700 10668
rect 198740 10616 198792 10668
rect 201500 10616 201552 10668
rect 202880 10616 202932 10668
rect 205088 10616 205140 10668
rect 205180 10616 205232 10668
rect 106188 10548 106240 10600
rect 206008 10548 206060 10600
rect 206100 10548 206152 10600
rect 212724 10548 212776 10600
rect 213276 10548 213328 10600
rect 219992 10548 220044 10600
rect 109868 10480 109920 10532
rect 206836 10480 206888 10532
rect 206928 10480 206980 10532
rect 211160 10480 211212 10532
rect 211252 10480 211304 10532
rect 217876 10480 217928 10532
rect 218796 10480 218848 10532
rect 225144 10548 225196 10600
rect 238944 10548 238996 10600
rect 239404 10548 239456 10600
rect 245384 10548 245436 10600
rect 250812 10548 250864 10600
rect 258816 10548 258868 10600
rect 229744 10480 229796 10532
rect 238852 10480 238904 10532
rect 246948 10480 247000 10532
rect 247224 10480 247276 10532
rect 258724 10480 258776 10532
rect 122564 10412 122616 10464
rect 199292 10412 199344 10464
rect 199384 10412 199436 10464
rect 203432 10412 203484 10464
rect 203524 10412 203576 10464
rect 205180 10412 205232 10464
rect 205640 10412 205692 10464
rect 209964 10412 210016 10464
rect 210240 10412 210292 10464
rect 240416 10412 240468 10464
rect 241520 10412 241572 10464
rect 251916 10412 251968 10464
rect 256976 10412 257028 10464
rect 354496 11024 354548 11076
rect 262036 10956 262088 11008
rect 362408 11024 362460 11076
rect 362592 11092 362644 11144
rect 267096 10888 267148 10940
rect 361396 10956 361448 11008
rect 363420 10956 363472 11008
rect 368020 10956 368072 11008
rect 355416 10888 355468 10940
rect 362592 10888 362644 10940
rect 364984 10888 365036 10940
rect 272156 10820 272208 10872
rect 360292 10820 360344 10872
rect 363328 10820 363380 10872
rect 368940 10820 368992 10872
rect 354496 10752 354548 10804
rect 359556 10752 359608 10804
rect 361396 10752 361448 10804
rect 363696 10752 363748 10804
rect 364156 10752 364208 10804
rect 282276 10684 282328 10736
rect 360108 10684 360160 10736
rect 360660 10684 360712 10736
rect 364524 10684 364576 10736
rect 381544 11228 381596 11280
rect 382096 11228 382148 11280
rect 382464 11228 382516 11280
rect 383200 11228 383252 11280
rect 384672 11228 384724 11280
rect 385224 11228 385276 11280
rect 385960 11228 386012 11280
rect 386512 11228 386564 11280
rect 374460 10752 374512 10804
rect 380348 10752 380400 10804
rect 287428 10616 287480 10668
rect 292580 10548 292632 10600
rect 360200 10548 360252 10600
rect 360568 10616 360620 10668
rect 365812 10616 365864 10668
rect 381544 10684 381596 10736
rect 382464 10616 382516 10668
rect 363420 10548 363472 10600
rect 367100 10548 367152 10600
rect 374460 10548 374512 10600
rect 379980 10548 380032 10600
rect 383568 10956 383620 11008
rect 385868 11092 385920 11144
rect 387984 11228 388036 11280
rect 387064 11092 387116 11144
rect 385776 11024 385828 11076
rect 388996 11160 389048 11212
rect 389824 11228 389876 11280
rect 390652 11228 390704 11280
rect 391388 11228 391440 11280
rect 391940 11228 391992 11280
rect 392492 11228 392544 11280
rect 392860 11228 392912 11280
rect 393504 11228 393556 11280
rect 394056 11228 394108 11280
rect 394700 11228 394752 11280
rect 395160 11228 395212 11280
rect 395528 11228 395580 11280
rect 396264 11228 396316 11280
rect 397920 11228 397972 11280
rect 398472 11228 398524 11280
rect 390560 10956 390612 11008
rect 396080 10956 396132 11008
rect 397460 10956 397512 11008
rect 399300 11092 399352 11144
rect 399852 11092 399904 11144
rect 400680 11228 400732 11280
rect 400956 11228 401008 11280
rect 402336 11228 402388 11280
rect 403900 11228 403952 11280
rect 438860 11228 438912 11280
rect 440148 11228 440200 11280
rect 440424 11228 440476 11280
rect 440700 11228 440752 11280
rect 441804 11296 441856 11348
rect 442908 11296 442960 11348
rect 443184 11228 443236 11280
rect 443460 11228 443512 11280
rect 440332 11024 440384 11076
rect 400312 10956 400364 11008
rect 401968 10956 402020 11008
rect 403072 10956 403124 11008
rect 403624 10956 403676 11008
rect 440240 10956 440292 11008
rect 441620 10956 441672 11008
rect 442080 10956 442132 11008
rect 441712 10888 441764 10940
rect 442632 10956 442684 11008
rect 444012 11228 444064 11280
rect 444564 11228 444616 11280
rect 444748 11228 444800 11280
rect 445024 11228 445076 11280
rect 445300 11228 445352 11280
rect 445852 11364 445904 11416
rect 445852 11228 445904 11280
rect 446128 11228 446180 11280
rect 446680 11500 446732 11552
rect 446680 11296 446732 11348
rect 447784 11296 447836 11348
rect 448060 11296 448112 11348
rect 443092 10956 443144 11008
rect 447140 10956 447192 11008
rect 444380 10888 444432 10940
rect 447232 10888 447284 10940
rect 447692 10956 447744 11008
rect 448336 10888 448388 10940
rect 478880 10956 478932 11008
rect 480720 11228 480772 11280
rect 481272 11228 481324 11280
rect 481824 11296 481876 11348
rect 480352 10956 480404 11008
rect 480260 10888 480312 10940
rect 481180 11092 481232 11144
rect 482100 11228 482152 11280
rect 482284 11228 482336 11280
rect 482836 11296 482888 11348
rect 483112 11296 483164 11348
rect 483664 11364 483716 11416
rect 483664 11228 483716 11280
rect 481640 10888 481692 10940
rect 483020 10888 483072 10940
rect 484216 11228 484268 11280
rect 484492 11296 484544 11348
rect 486148 11296 486200 11348
rect 486424 11228 486476 11280
rect 486700 11296 486752 11348
rect 486976 11296 487028 11348
rect 487252 11228 487304 11280
rect 487528 11228 487580 11280
rect 487804 11228 487856 11280
rect 488080 11228 488132 11280
rect 488356 11228 488408 11280
rect 488540 11296 488592 11348
rect 488816 11296 488868 11348
rect 484124 10956 484176 11008
rect 484952 10956 485004 11008
rect 485044 10956 485096 11008
rect 484308 10888 484360 10940
rect 485780 11092 485832 11144
rect 297732 10480 297784 10532
rect 370136 10480 370188 10532
rect 302424 10412 302476 10464
rect 371056 10412 371108 10464
rect 378140 10412 378192 10464
rect 385224 10412 385276 10464
rect 145748 10344 145800 10396
rect 205824 10344 205876 10396
rect 210332 10344 210384 10396
rect 220084 10344 220136 10396
rect 220176 10344 220228 10396
rect 230848 10344 230900 10396
rect 239036 10344 239088 10396
rect 249064 10344 249116 10396
rect 307484 10344 307536 10396
rect 372160 10344 372212 10396
rect 376852 10344 376904 10396
rect 383200 10344 383252 10396
rect 56600 10276 56652 10328
rect 145840 10276 145892 10328
rect 149704 10276 149756 10328
rect 205640 10276 205692 10328
rect 210148 10276 210200 10328
rect 212356 10276 212408 10328
rect 212448 10276 212500 10328
rect 217600 10276 217652 10328
rect 217876 10276 217928 10328
rect 220912 10276 220964 10328
rect 251916 10276 251968 10328
rect 258632 10276 258684 10328
rect 312452 10276 312504 10328
rect 373264 10276 373316 10328
rect 382188 10276 382240 10328
rect 385960 10276 386012 10328
rect 95148 10208 95200 10260
rect 176660 10208 176712 10260
rect 187884 10208 187936 10260
rect 198464 10208 198516 10260
rect 198648 10208 198700 10260
rect 205364 10208 205416 10260
rect 206008 10208 206060 10260
rect 213920 10208 213972 10260
rect 214104 10208 214156 10260
rect 316316 10208 316368 10260
rect 317512 10208 317564 10260
rect 374368 10208 374420 10260
rect 382924 10208 382976 10260
rect 386512 10208 386564 10260
rect 173072 10140 173124 10192
rect 225788 10140 225840 10192
rect 322480 10140 322532 10192
rect 375472 10140 375524 10192
rect 112812 10072 112864 10124
rect 175372 10072 175424 10124
rect 176292 10072 176344 10124
rect 227352 10072 227404 10124
rect 332508 10072 332560 10124
rect 377588 10072 377640 10124
rect 93768 10004 93820 10056
rect 186228 10004 186280 10056
rect 186320 10004 186372 10056
rect 205640 10004 205692 10056
rect 92112 9936 92164 9988
rect 195060 9936 195112 9988
rect 195152 9936 195204 9988
rect 198372 9936 198424 9988
rect 198556 9936 198608 9988
rect 202880 9936 202932 9988
rect 203616 9936 203668 9988
rect 206744 10004 206796 10056
rect 206836 10004 206888 10056
rect 217232 10004 217284 10056
rect 219992 10004 220044 10056
rect 321284 10004 321336 10056
rect 337476 10004 337528 10056
rect 378692 10004 378744 10056
rect 205824 9936 205876 9988
rect 214012 9936 214064 9988
rect 218428 9936 218480 9988
rect 326344 9936 326396 9988
rect 340144 9936 340196 9988
rect 379428 9936 379480 9988
rect 178040 9868 178092 9920
rect 211252 9868 211304 9920
rect 213828 9868 213880 9920
rect 229652 9868 229704 9920
rect 262404 9868 262456 9920
rect 368572 9868 368624 9920
rect 67574 9766 67626 9818
rect 67638 9766 67690 9818
rect 67702 9766 67754 9818
rect 67766 9766 67818 9818
rect 67830 9766 67882 9818
rect 199502 9766 199554 9818
rect 199566 9766 199618 9818
rect 199630 9766 199682 9818
rect 199694 9766 199746 9818
rect 199758 9766 199810 9818
rect 331430 9766 331482 9818
rect 331494 9766 331546 9818
rect 331558 9766 331610 9818
rect 331622 9766 331674 9818
rect 331686 9766 331738 9818
rect 463358 9766 463410 9818
rect 463422 9766 463474 9818
rect 463486 9766 463538 9818
rect 463550 9766 463602 9818
rect 463614 9766 463666 9818
rect 127808 9664 127860 9716
rect 186596 9664 186648 9716
rect 198464 9664 198516 9716
rect 200856 9664 200908 9716
rect 200948 9664 201000 9716
rect 205272 9664 205324 9716
rect 205548 9664 205600 9716
rect 306380 9664 306432 9716
rect 123392 9596 123444 9648
rect 82452 9460 82504 9512
rect 74724 9392 74776 9444
rect 167092 9392 167144 9444
rect 171784 9528 171836 9580
rect 178040 9528 178092 9580
rect 184388 9571 184440 9580
rect 184388 9537 184397 9571
rect 184397 9537 184431 9571
rect 184431 9537 184440 9571
rect 184388 9528 184440 9537
rect 191472 9528 191524 9580
rect 195888 9571 195940 9580
rect 195888 9537 195897 9571
rect 195897 9537 195931 9571
rect 195931 9537 195940 9571
rect 195888 9528 195940 9537
rect 167368 9460 167420 9512
rect 194692 9503 194744 9512
rect 194692 9469 194701 9503
rect 194701 9469 194735 9503
rect 194735 9469 194744 9503
rect 194692 9460 194744 9469
rect 90180 9324 90232 9376
rect 191472 9367 191524 9376
rect 191472 9333 191481 9367
rect 191481 9333 191515 9367
rect 191515 9333 191524 9367
rect 191472 9324 191524 9333
rect 203616 9571 203668 9580
rect 203616 9537 203625 9571
rect 203625 9537 203659 9571
rect 203659 9537 203668 9571
rect 203616 9528 203668 9537
rect 206284 9571 206336 9580
rect 206284 9537 206293 9571
rect 206293 9537 206327 9571
rect 206327 9537 206336 9571
rect 206284 9528 206336 9537
rect 211068 9571 211120 9580
rect 211068 9537 211077 9571
rect 211077 9537 211111 9571
rect 211111 9537 211120 9571
rect 211068 9528 211120 9537
rect 213828 9571 213880 9580
rect 213828 9537 213837 9571
rect 213837 9537 213871 9571
rect 213871 9537 213880 9571
rect 213828 9528 213880 9537
rect 202420 9503 202472 9512
rect 202420 9469 202429 9503
rect 202429 9469 202463 9503
rect 202463 9469 202472 9503
rect 202420 9460 202472 9469
rect 205456 9503 205508 9512
rect 205456 9469 205465 9503
rect 205465 9469 205499 9503
rect 205499 9469 205508 9503
rect 205456 9460 205508 9469
rect 210240 9503 210292 9512
rect 210240 9469 210249 9503
rect 210249 9469 210283 9503
rect 210283 9469 210292 9503
rect 210240 9460 210292 9469
rect 212540 9460 212592 9512
rect 217968 9503 218020 9512
rect 217968 9469 217977 9503
rect 217977 9469 218011 9503
rect 218011 9469 218020 9503
rect 217968 9460 218020 9469
rect 218796 9639 218848 9648
rect 218796 9605 218805 9639
rect 218805 9605 218839 9639
rect 218839 9605 218848 9639
rect 218796 9596 218848 9605
rect 221372 9639 221424 9648
rect 221372 9605 221381 9639
rect 221381 9605 221415 9639
rect 221415 9605 221424 9639
rect 221372 9596 221424 9605
rect 248604 9596 248656 9648
rect 340144 9639 340196 9648
rect 229100 9528 229152 9580
rect 220360 9460 220412 9512
rect 220544 9503 220596 9512
rect 220544 9469 220553 9503
rect 220553 9469 220587 9503
rect 220587 9469 220596 9503
rect 220544 9460 220596 9469
rect 224684 9503 224736 9512
rect 224684 9469 224693 9503
rect 224693 9469 224727 9503
rect 224727 9469 224736 9503
rect 224684 9460 224736 9469
rect 228272 9503 228324 9512
rect 228272 9469 228281 9503
rect 228281 9469 228315 9503
rect 228315 9469 228324 9503
rect 228272 9460 228324 9469
rect 232044 9460 232096 9512
rect 200764 9392 200816 9444
rect 232320 9392 232372 9444
rect 234436 9528 234488 9580
rect 236000 9503 236052 9512
rect 236000 9469 236009 9503
rect 236009 9469 236043 9503
rect 236043 9469 236052 9503
rect 236000 9460 236052 9469
rect 239956 9571 240008 9580
rect 239956 9537 239965 9571
rect 239965 9537 239999 9571
rect 239999 9537 240008 9571
rect 239956 9528 240008 9537
rect 244004 9571 244056 9580
rect 244004 9537 244013 9571
rect 244013 9537 244047 9571
rect 244047 9537 244056 9571
rect 244004 9528 244056 9537
rect 340144 9605 340153 9639
rect 340153 9605 340187 9639
rect 340187 9605 340196 9639
rect 340144 9596 340196 9605
rect 342720 9639 342772 9648
rect 342720 9605 342729 9639
rect 342729 9605 342763 9639
rect 342763 9605 342772 9639
rect 342720 9596 342772 9605
rect 382096 9664 382148 9716
rect 346768 9571 346820 9580
rect 346768 9537 346777 9571
rect 346777 9537 346811 9571
rect 346811 9537 346820 9571
rect 346768 9528 346820 9537
rect 347596 9571 347648 9580
rect 347596 9537 347605 9571
rect 347605 9537 347639 9571
rect 347639 9537 347648 9571
rect 347596 9528 347648 9537
rect 350080 9528 350132 9580
rect 236828 9503 236880 9512
rect 236828 9469 236837 9503
rect 236837 9469 236871 9503
rect 236871 9469 236880 9503
rect 236828 9460 236880 9469
rect 239680 9503 239732 9512
rect 239680 9469 239689 9503
rect 239689 9469 239723 9503
rect 239723 9469 239732 9503
rect 239680 9460 239732 9469
rect 243728 9503 243780 9512
rect 243728 9469 243737 9503
rect 243737 9469 243771 9503
rect 243771 9469 243780 9503
rect 243728 9460 243780 9469
rect 338948 9503 339000 9512
rect 338948 9469 338957 9503
rect 338957 9469 338991 9503
rect 338991 9469 339000 9503
rect 338948 9460 339000 9469
rect 344100 9503 344152 9512
rect 344100 9469 344109 9503
rect 344109 9469 344143 9503
rect 344143 9469 344152 9503
rect 344100 9460 344152 9469
rect 349344 9503 349396 9512
rect 349344 9469 349353 9503
rect 349353 9469 349387 9503
rect 349387 9469 349396 9503
rect 349344 9460 349396 9469
rect 351920 9503 351972 9512
rect 351920 9469 351929 9503
rect 351929 9469 351963 9503
rect 351963 9469 351972 9503
rect 351920 9460 351972 9469
rect 354404 9596 354456 9648
rect 354588 9596 354640 9648
rect 355324 9528 355376 9580
rect 357900 9528 357952 9580
rect 358636 9571 358688 9580
rect 358636 9537 358645 9571
rect 358645 9537 358679 9571
rect 358679 9537 358688 9571
rect 358636 9528 358688 9537
rect 367284 9596 367336 9648
rect 368572 9639 368624 9648
rect 368572 9605 368581 9639
rect 368581 9605 368615 9639
rect 368615 9605 368624 9639
rect 368572 9596 368624 9605
rect 199200 9324 199252 9376
rect 229100 9367 229152 9376
rect 229100 9333 229109 9367
rect 229109 9333 229143 9367
rect 229143 9333 229152 9367
rect 229100 9324 229152 9333
rect 241520 9324 241572 9376
rect 244004 9324 244056 9376
rect 255688 9324 255740 9376
rect 260196 9324 260248 9376
rect 354588 9392 354640 9444
rect 357072 9503 357124 9512
rect 357072 9469 357081 9503
rect 357081 9469 357115 9503
rect 357115 9469 357124 9503
rect 357072 9460 357124 9469
rect 360200 9460 360252 9512
rect 362132 9503 362184 9512
rect 362132 9469 362141 9503
rect 362141 9469 362175 9503
rect 362175 9469 362184 9503
rect 362132 9460 362184 9469
rect 363696 9503 363748 9512
rect 363696 9469 363705 9503
rect 363705 9469 363739 9503
rect 363739 9469 363748 9503
rect 363696 9460 363748 9469
rect 368848 9571 368900 9580
rect 368848 9537 368857 9571
rect 368857 9537 368891 9571
rect 368891 9537 368900 9571
rect 368848 9528 368900 9537
rect 379244 9596 379296 9648
rect 371332 9571 371384 9580
rect 371332 9537 371341 9571
rect 371341 9537 371375 9571
rect 371375 9537 371384 9571
rect 371332 9528 371384 9537
rect 374276 9528 374328 9580
rect 371056 9503 371108 9512
rect 371056 9469 371065 9503
rect 371065 9469 371099 9503
rect 371099 9469 371108 9503
rect 371056 9460 371108 9469
rect 372712 9460 372764 9512
rect 373540 9460 373592 9512
rect 375932 9503 375984 9512
rect 375932 9469 375941 9503
rect 375941 9469 375975 9503
rect 375975 9469 375984 9503
rect 375932 9460 375984 9469
rect 376760 9528 376812 9580
rect 378324 9503 378376 9512
rect 378324 9469 378333 9503
rect 378333 9469 378367 9503
rect 378367 9469 378376 9503
rect 378324 9460 378376 9469
rect 379152 9528 379204 9580
rect 382188 9596 382240 9648
rect 350080 9367 350132 9376
rect 350080 9333 350089 9367
rect 350089 9333 350123 9367
rect 350123 9333 350132 9367
rect 350080 9324 350132 9333
rect 355324 9367 355376 9376
rect 355324 9333 355333 9367
rect 355333 9333 355367 9367
rect 355367 9333 355376 9367
rect 355324 9324 355376 9333
rect 357900 9367 357952 9376
rect 357900 9333 357909 9367
rect 357909 9333 357943 9367
rect 357943 9333 357952 9367
rect 357900 9324 357952 9333
rect 373632 9392 373684 9444
rect 373816 9392 373868 9444
rect 379980 9460 380032 9512
rect 380808 9503 380860 9512
rect 380808 9469 380817 9503
rect 380817 9469 380851 9503
rect 380851 9469 380860 9503
rect 380808 9460 380860 9469
rect 388996 9596 389048 9648
rect 383016 9460 383068 9512
rect 385776 9392 385828 9444
rect 367100 9324 367152 9376
rect 367284 9367 367336 9376
rect 367284 9333 367293 9367
rect 367293 9333 367327 9367
rect 367327 9333 367336 9367
rect 367284 9324 367336 9333
rect 368848 9324 368900 9376
rect 373540 9324 373592 9376
rect 374276 9367 374328 9376
rect 374276 9333 374285 9367
rect 374285 9333 374319 9367
rect 374319 9333 374328 9367
rect 374276 9324 374328 9333
rect 376760 9367 376812 9376
rect 376760 9333 376769 9367
rect 376769 9333 376803 9367
rect 376803 9333 376812 9367
rect 376760 9324 376812 9333
rect 379152 9367 379204 9376
rect 379152 9333 379161 9367
rect 379161 9333 379195 9367
rect 379195 9333 379204 9367
rect 379152 9324 379204 9333
rect 379244 9324 379296 9376
rect 384672 9324 384724 9376
rect 66914 9222 66966 9274
rect 66978 9222 67030 9274
rect 67042 9222 67094 9274
rect 67106 9222 67158 9274
rect 67170 9222 67222 9274
rect 198842 9222 198894 9274
rect 198906 9222 198958 9274
rect 198970 9222 199022 9274
rect 199034 9222 199086 9274
rect 199098 9222 199150 9274
rect 330770 9222 330822 9274
rect 330834 9222 330886 9274
rect 330898 9222 330950 9274
rect 330962 9222 331014 9274
rect 331026 9222 331078 9274
rect 462698 9222 462750 9274
rect 462762 9222 462814 9274
rect 462826 9222 462878 9274
rect 462890 9222 462942 9274
rect 462954 9222 463006 9274
rect 87604 9120 87656 9172
rect 194692 9120 194744 9172
rect 194968 9120 195020 9172
rect 215392 9120 215444 9172
rect 232872 9120 232924 9172
rect 338948 9120 339000 9172
rect 357440 9120 357492 9172
rect 375932 9120 375984 9172
rect 376760 9120 376812 9172
rect 387984 9120 388036 9172
rect 110788 9052 110840 9104
rect 217968 9052 218020 9104
rect 229100 9052 229152 9104
rect 250260 9052 250312 9104
rect 265348 9052 265400 9104
rect 371056 9052 371108 9104
rect 374276 9052 374328 9104
rect 385868 9052 385920 9104
rect 43812 8848 43864 8900
rect 168748 8984 168800 9036
rect 160100 8891 160152 8900
rect 160100 8857 160109 8891
rect 160109 8857 160143 8891
rect 160143 8857 160152 8891
rect 160100 8848 160152 8857
rect 167552 8891 167604 8900
rect 167552 8857 167561 8891
rect 167561 8857 167595 8891
rect 167595 8857 167604 8891
rect 167552 8848 167604 8857
rect 171784 8916 171836 8968
rect 173072 8959 173124 8968
rect 173072 8925 173081 8959
rect 173081 8925 173115 8959
rect 173115 8925 173124 8959
rect 173072 8916 173124 8925
rect 176292 8959 176344 8968
rect 176292 8925 176301 8959
rect 176301 8925 176335 8959
rect 176335 8925 176344 8959
rect 176292 8916 176344 8925
rect 168748 8780 168800 8832
rect 171232 8848 171284 8900
rect 175280 8891 175332 8900
rect 175280 8857 175289 8891
rect 175289 8857 175323 8891
rect 175323 8857 175332 8891
rect 175280 8848 175332 8857
rect 175464 8780 175516 8832
rect 176752 8984 176804 9036
rect 239680 8984 239732 9036
rect 239956 8984 240008 9036
rect 251180 8984 251232 9036
rect 275652 8984 275704 9036
rect 380808 8984 380860 9036
rect 187516 8916 187568 8968
rect 179420 8891 179472 8900
rect 179420 8857 179429 8891
rect 179429 8857 179463 8891
rect 179463 8857 179472 8891
rect 179420 8848 179472 8857
rect 186412 8848 186464 8900
rect 187700 8916 187752 8968
rect 229192 8916 229244 8968
rect 236828 8916 236880 8968
rect 254032 8916 254084 8968
rect 321284 8959 321336 8968
rect 321284 8925 321293 8959
rect 321293 8925 321327 8959
rect 321327 8925 321336 8959
rect 321284 8916 321336 8925
rect 322480 8959 322532 8968
rect 322480 8925 322489 8959
rect 322489 8925 322523 8959
rect 322523 8925 322532 8959
rect 322480 8916 322532 8925
rect 326344 8959 326396 8968
rect 326344 8925 326353 8959
rect 326353 8925 326387 8959
rect 326387 8925 326396 8959
rect 326344 8916 326396 8925
rect 327540 8916 327592 8968
rect 332508 8959 332560 8968
rect 332508 8925 332517 8959
rect 332517 8925 332551 8959
rect 332551 8925 332560 8959
rect 332508 8916 332560 8925
rect 336280 8959 336332 8968
rect 336280 8925 336289 8959
rect 336289 8925 336323 8959
rect 336323 8925 336332 8959
rect 336280 8916 336332 8925
rect 337476 8959 337528 8968
rect 337476 8925 337485 8959
rect 337485 8925 337519 8959
rect 337519 8925 337528 8959
rect 337476 8916 337528 8925
rect 355324 8916 355376 8968
rect 364156 8916 364208 8968
rect 365812 8916 365864 8968
rect 378324 8916 378376 8968
rect 187516 8780 187568 8832
rect 187792 8848 187844 8900
rect 212448 8848 212500 8900
rect 224132 8848 224184 8900
rect 200764 8780 200816 8832
rect 362132 8848 362184 8900
rect 383568 8848 383620 8900
rect 327540 8823 327592 8832
rect 327540 8789 327549 8823
rect 327549 8789 327583 8823
rect 327583 8789 327592 8823
rect 327540 8780 327592 8789
rect 371332 8780 371384 8832
rect 382924 8780 382976 8832
rect 67574 8678 67626 8730
rect 67638 8678 67690 8730
rect 67702 8678 67754 8730
rect 67766 8678 67818 8730
rect 67830 8678 67882 8730
rect 199502 8678 199554 8730
rect 199566 8678 199618 8730
rect 199630 8678 199682 8730
rect 199694 8678 199746 8730
rect 199758 8678 199810 8730
rect 331430 8678 331482 8730
rect 331494 8678 331546 8730
rect 331558 8678 331610 8730
rect 331622 8678 331674 8730
rect 331686 8678 331738 8730
rect 463358 8678 463410 8730
rect 463422 8678 463474 8730
rect 463486 8678 463538 8730
rect 463550 8678 463602 8730
rect 463614 8678 463666 8730
rect 135260 8576 135312 8628
rect 167552 8576 167604 8628
rect 175372 8576 175424 8628
rect 219900 8576 219952 8628
rect 302424 8619 302476 8628
rect 302424 8585 302433 8619
rect 302433 8585 302467 8619
rect 302467 8585 302476 8619
rect 302424 8576 302476 8585
rect 307484 8619 307536 8628
rect 307484 8585 307493 8619
rect 307493 8585 307527 8619
rect 307527 8585 307536 8619
rect 307484 8576 307536 8585
rect 312452 8619 312504 8628
rect 312452 8585 312461 8619
rect 312461 8585 312495 8619
rect 312495 8585 312504 8619
rect 312452 8576 312504 8585
rect 312912 8576 312964 8628
rect 351920 8576 351972 8628
rect 357900 8576 357952 8628
rect 376852 8576 376904 8628
rect 379152 8576 379204 8628
rect 387064 8576 387116 8628
rect 36084 8372 36136 8424
rect 145748 8551 145800 8560
rect 145748 8517 145757 8551
rect 145757 8517 145791 8551
rect 145791 8517 145800 8551
rect 145748 8508 145800 8517
rect 145840 8508 145892 8560
rect 195612 8508 195664 8560
rect 198648 8508 198700 8560
rect 199200 8508 199252 8560
rect 237380 8508 237432 8560
rect 242164 8508 242216 8560
rect 349344 8508 349396 8560
rect 350080 8508 350132 8560
rect 364984 8508 365036 8560
rect 367284 8508 367336 8560
rect 378140 8508 378192 8560
rect 33508 8304 33560 8356
rect 149704 8483 149756 8492
rect 149704 8449 149713 8483
rect 149713 8449 149747 8483
rect 149747 8449 149756 8483
rect 149704 8440 149756 8449
rect 157892 8483 157944 8492
rect 157892 8449 157901 8483
rect 157901 8449 157935 8483
rect 157935 8449 157944 8483
rect 157892 8440 157944 8449
rect 222476 8440 222528 8492
rect 302424 8440 302476 8492
rect 306380 8483 306432 8492
rect 306380 8449 306389 8483
rect 306389 8449 306423 8483
rect 306423 8449 306432 8483
rect 306380 8440 306432 8449
rect 307484 8440 307536 8492
rect 311256 8483 311308 8492
rect 311256 8449 311265 8483
rect 311265 8449 311299 8483
rect 311299 8449 311308 8483
rect 311256 8440 311308 8449
rect 312452 8440 312504 8492
rect 316316 8483 316368 8492
rect 316316 8449 316325 8483
rect 316325 8449 316359 8483
rect 316359 8449 316368 8483
rect 316316 8440 316368 8449
rect 317512 8483 317564 8492
rect 317512 8449 317521 8483
rect 317521 8449 317555 8483
rect 317555 8449 317564 8483
rect 317512 8440 317564 8449
rect 149060 8372 149112 8424
rect 156696 8415 156748 8424
rect 156696 8381 156705 8415
rect 156705 8381 156739 8415
rect 156739 8381 156748 8415
rect 156696 8372 156748 8381
rect 191472 8372 191524 8424
rect 233884 8372 233936 8424
rect 301228 8415 301280 8424
rect 301228 8381 301237 8415
rect 301237 8381 301271 8415
rect 301271 8381 301280 8415
rect 301228 8372 301280 8381
rect 366272 8372 366324 8424
rect 367468 8372 367520 8424
rect 85580 8236 85632 8288
rect 186320 8304 186372 8356
rect 198740 8304 198792 8356
rect 276020 8304 276072 8356
rect 160100 8236 160152 8288
rect 186504 8236 186556 8288
rect 201960 8236 202012 8288
rect 202052 8236 202104 8288
rect 207480 8236 207532 8288
rect 361488 8236 361540 8288
rect 400956 8236 401008 8288
rect 430212 8236 430264 8288
rect 448336 8304 448388 8356
rect 447048 8236 447100 8288
rect 448060 8236 448112 8288
rect 481824 8236 481876 8288
rect 483112 8236 483164 8288
rect 486148 8236 486200 8288
rect 488540 8236 488592 8288
rect 66914 8134 66966 8186
rect 66978 8134 67030 8186
rect 67042 8134 67094 8186
rect 67106 8134 67158 8186
rect 67170 8134 67222 8186
rect 198842 8134 198894 8186
rect 198906 8134 198958 8186
rect 198970 8134 199022 8186
rect 199034 8134 199086 8186
rect 199098 8134 199150 8186
rect 330770 8134 330822 8186
rect 330834 8134 330886 8186
rect 330898 8134 330950 8186
rect 330962 8134 331014 8186
rect 331026 8134 331078 8186
rect 462698 8134 462750 8186
rect 462762 8134 462814 8186
rect 462826 8134 462878 8186
rect 462890 8134 462942 8186
rect 462954 8134 463006 8186
rect 35900 8032 35952 8084
rect 101312 8032 101364 8084
rect 122564 8075 122616 8084
rect 122564 8041 122573 8075
rect 122573 8041 122607 8075
rect 122607 8041 122616 8075
rect 122564 8032 122616 8041
rect 123300 8032 123352 8084
rect 221648 8032 221700 8084
rect 277124 8075 277176 8084
rect 277124 8041 277133 8075
rect 277133 8041 277167 8075
rect 277167 8041 277176 8075
rect 277124 8032 277176 8041
rect 282276 8075 282328 8084
rect 282276 8041 282285 8075
rect 282285 8041 282319 8075
rect 282319 8041 282328 8075
rect 282276 8032 282328 8041
rect 287152 8032 287204 8084
rect 287428 8075 287480 8084
rect 287428 8041 287437 8075
rect 287437 8041 287471 8075
rect 287471 8041 287480 8075
rect 287428 8032 287480 8041
rect 292580 8075 292632 8084
rect 292580 8041 292589 8075
rect 292589 8041 292623 8075
rect 292623 8041 292632 8075
rect 292580 8032 292632 8041
rect 293868 8032 293920 8084
rect 378416 8032 378468 8084
rect 392124 8032 392176 8084
rect 394700 8032 394752 8084
rect 445576 8032 445628 8084
rect 447048 8032 447100 8084
rect 481732 8032 481784 8084
rect 484492 8032 484544 8084
rect 487528 8032 487580 8084
rect 501328 8032 501380 8084
rect 59268 7964 59320 8016
rect 135260 7964 135312 8016
rect 139032 7964 139084 8016
rect 246120 7964 246172 8016
rect 267648 7964 267700 8016
rect 364248 7964 364300 8016
rect 365720 7964 365772 8016
rect 371792 7964 371844 8016
rect 372528 7964 372580 8016
rect 376208 7964 376260 8016
rect 382280 7964 382332 8016
rect 402336 7964 402388 8016
rect 426164 7964 426216 8016
rect 447784 7964 447836 8016
rect 482008 7964 482060 8016
rect 485044 7964 485096 8016
rect 486976 7964 487028 8016
rect 496176 7964 496228 8016
rect 22468 7896 22520 7948
rect 99472 7896 99524 7948
rect 121000 7896 121052 7948
rect 228456 7896 228508 7948
rect 276020 7939 276072 7948
rect 276020 7905 276029 7939
rect 276029 7905 276063 7939
rect 276063 7905 276072 7939
rect 276020 7896 276072 7905
rect 71044 7828 71096 7880
rect 86316 7828 86368 7880
rect 42984 7760 43036 7812
rect 91376 7828 91428 7880
rect 14740 7692 14792 7744
rect 91284 7760 91336 7812
rect 86592 7692 86644 7744
rect 96712 7871 96764 7880
rect 91836 7760 91888 7812
rect 96712 7837 96721 7871
rect 96721 7837 96755 7871
rect 96755 7837 96764 7871
rect 96712 7828 96764 7837
rect 114836 7828 114888 7880
rect 122564 7828 122616 7880
rect 92848 7803 92900 7812
rect 92848 7769 92857 7803
rect 92857 7769 92891 7803
rect 92891 7769 92900 7803
rect 92848 7760 92900 7769
rect 91744 7692 91796 7744
rect 94044 7735 94096 7744
rect 94044 7701 94053 7735
rect 94053 7701 94087 7735
rect 94087 7701 94096 7735
rect 94044 7692 94096 7701
rect 95240 7735 95292 7744
rect 95240 7701 95249 7735
rect 95249 7701 95283 7735
rect 95283 7701 95292 7735
rect 95240 7692 95292 7701
rect 97632 7735 97684 7744
rect 97632 7701 97641 7735
rect 97641 7701 97675 7735
rect 97675 7701 97684 7735
rect 97632 7692 97684 7701
rect 113640 7803 113692 7812
rect 113640 7769 113649 7803
rect 113649 7769 113683 7803
rect 113683 7769 113692 7803
rect 113640 7760 113692 7769
rect 126336 7803 126388 7812
rect 126336 7769 126345 7803
rect 126345 7769 126379 7803
rect 126379 7769 126388 7803
rect 126336 7760 126388 7769
rect 131396 7803 131448 7812
rect 131396 7769 131405 7803
rect 131405 7769 131439 7803
rect 131439 7769 131448 7803
rect 131396 7760 131448 7769
rect 132040 7828 132092 7880
rect 136640 7803 136692 7812
rect 136640 7769 136649 7803
rect 136649 7769 136683 7803
rect 136683 7769 136692 7803
rect 136640 7760 136692 7769
rect 141240 7828 141292 7880
rect 149704 7828 149756 7880
rect 268384 7828 268436 7880
rect 277124 7828 277176 7880
rect 282276 7828 282328 7880
rect 287152 7828 287204 7880
rect 239496 7760 239548 7812
rect 114836 7735 114888 7744
rect 114836 7701 114845 7735
rect 114845 7701 114879 7735
rect 114879 7701 114888 7735
rect 114836 7692 114888 7701
rect 127716 7735 127768 7744
rect 127716 7701 127725 7735
rect 127725 7701 127759 7735
rect 127759 7701 127768 7735
rect 127716 7692 127768 7701
rect 132868 7735 132920 7744
rect 132868 7701 132877 7735
rect 132877 7701 132911 7735
rect 132911 7701 132920 7735
rect 132868 7692 132920 7701
rect 186596 7692 186648 7744
rect 234988 7692 235040 7744
rect 251456 7692 251508 7744
rect 252468 7735 252520 7744
rect 252468 7701 252477 7735
rect 252477 7701 252511 7735
rect 252511 7701 252520 7735
rect 252468 7692 252520 7701
rect 258356 7692 258408 7744
rect 280344 7760 280396 7812
rect 286140 7803 286192 7812
rect 286140 7769 286149 7803
rect 286149 7769 286183 7803
rect 286183 7769 286192 7803
rect 286140 7760 286192 7769
rect 291200 7803 291252 7812
rect 291200 7769 291209 7803
rect 291209 7769 291243 7803
rect 291243 7769 291252 7803
rect 291200 7760 291252 7769
rect 292580 7828 292632 7880
rect 297732 7871 297784 7880
rect 297732 7837 297741 7871
rect 297741 7837 297775 7871
rect 297775 7837 297784 7871
rect 297732 7828 297784 7837
rect 364708 7896 364760 7948
rect 366272 7828 366324 7880
rect 367100 7896 367152 7948
rect 372896 7896 372948 7948
rect 375564 7896 375616 7948
rect 400680 7896 400732 7948
rect 480444 7896 480496 7948
rect 483664 7896 483716 7948
rect 487804 7896 487856 7948
rect 503904 7896 503956 7948
rect 392860 7828 392912 7880
rect 419908 7828 419960 7880
rect 447232 7828 447284 7880
rect 487252 7828 487304 7880
rect 498752 7828 498804 7880
rect 296168 7803 296220 7812
rect 296168 7769 296177 7803
rect 296177 7769 296211 7803
rect 296211 7769 296220 7803
rect 296168 7760 296220 7769
rect 366364 7760 366416 7812
rect 368480 7760 368532 7812
rect 374000 7760 374052 7812
rect 374276 7760 374328 7812
rect 393504 7760 393556 7812
rect 393964 7760 394016 7812
rect 440148 7760 440200 7812
rect 488080 7760 488132 7812
rect 506480 7760 506532 7812
rect 349068 7692 349120 7744
rect 403900 7692 403952 7744
rect 414756 7692 414808 7744
rect 446680 7692 446732 7744
rect 488356 7692 488408 7744
rect 509056 7692 509108 7744
rect 67574 7590 67626 7642
rect 67638 7590 67690 7642
rect 67702 7590 67754 7642
rect 67766 7590 67818 7642
rect 67830 7590 67882 7642
rect 199502 7590 199554 7642
rect 199566 7590 199618 7642
rect 199630 7590 199682 7642
rect 199694 7590 199746 7642
rect 199758 7590 199810 7642
rect 331430 7590 331482 7642
rect 331494 7590 331546 7642
rect 331558 7590 331610 7642
rect 331622 7590 331674 7642
rect 331686 7590 331738 7642
rect 463358 7590 463410 7642
rect 463422 7590 463474 7642
rect 463486 7590 463538 7642
rect 463550 7590 463602 7642
rect 463614 7590 463666 7642
rect 29920 7488 29972 7540
rect 97632 7488 97684 7540
rect 63500 7420 63552 7472
rect 95240 7420 95292 7472
rect 92204 7352 92256 7404
rect 93492 7395 93544 7404
rect 93492 7361 93501 7395
rect 93501 7361 93535 7395
rect 93535 7361 93544 7395
rect 93492 7352 93544 7361
rect 96068 7463 96120 7472
rect 96068 7429 96077 7463
rect 96077 7429 96111 7463
rect 96111 7429 96120 7463
rect 96068 7420 96120 7429
rect 97264 7463 97316 7472
rect 97264 7429 97273 7463
rect 97273 7429 97307 7463
rect 97307 7429 97316 7463
rect 97264 7420 97316 7429
rect 92388 7284 92440 7336
rect 94044 7284 94096 7336
rect 96712 7395 96764 7404
rect 96712 7361 96721 7395
rect 96721 7361 96755 7395
rect 96755 7361 96764 7395
rect 96712 7352 96764 7361
rect 98460 7463 98512 7472
rect 98460 7429 98469 7463
rect 98469 7429 98503 7463
rect 98503 7429 98512 7463
rect 98460 7420 98512 7429
rect 94872 7327 94924 7336
rect 94872 7293 94881 7327
rect 94881 7293 94915 7327
rect 94915 7293 94924 7327
rect 94872 7284 94924 7293
rect 96620 7284 96672 7336
rect 126336 7488 126388 7540
rect 127716 7488 127768 7540
rect 201500 7488 201552 7540
rect 237012 7488 237064 7540
rect 101864 7463 101916 7472
rect 101864 7429 101873 7463
rect 101873 7429 101907 7463
rect 101907 7429 101916 7463
rect 101864 7420 101916 7429
rect 99472 7395 99524 7404
rect 99472 7361 99481 7395
rect 99481 7361 99515 7395
rect 99515 7361 99524 7395
rect 99472 7352 99524 7361
rect 100668 7395 100720 7404
rect 100668 7361 100677 7395
rect 100677 7361 100711 7395
rect 100711 7361 100720 7395
rect 100668 7352 100720 7361
rect 101312 7395 101364 7404
rect 101312 7361 101321 7395
rect 101321 7361 101355 7395
rect 101355 7361 101364 7395
rect 101312 7352 101364 7361
rect 131396 7420 131448 7472
rect 141240 7420 141292 7472
rect 210700 7420 210752 7472
rect 250812 7463 250864 7472
rect 250812 7429 250821 7463
rect 250821 7429 250855 7463
rect 250855 7429 250864 7463
rect 250812 7420 250864 7429
rect 256976 7531 257028 7540
rect 256976 7497 256985 7531
rect 256985 7497 257019 7531
rect 257019 7497 257028 7531
rect 256976 7488 257028 7497
rect 262036 7531 262088 7540
rect 262036 7497 262045 7531
rect 262045 7497 262079 7531
rect 262079 7497 262088 7531
rect 262036 7488 262088 7497
rect 267096 7531 267148 7540
rect 267096 7497 267105 7531
rect 267105 7497 267139 7531
rect 267139 7497 267148 7531
rect 267096 7488 267148 7497
rect 272156 7531 272208 7540
rect 272156 7497 272165 7531
rect 272165 7497 272199 7531
rect 272199 7497 272208 7531
rect 272156 7488 272208 7497
rect 358820 7488 358872 7540
rect 368664 7488 368716 7540
rect 370780 7488 370832 7540
rect 375104 7488 375156 7540
rect 375380 7488 375432 7540
rect 394056 7488 394108 7540
rect 486424 7488 486476 7540
rect 491024 7488 491076 7540
rect 344100 7420 344152 7472
rect 362316 7420 362368 7472
rect 369768 7420 369820 7472
rect 373448 7420 373500 7472
rect 377312 7420 377364 7472
rect 486700 7420 486752 7472
rect 493600 7420 493652 7472
rect 90548 7191 90600 7200
rect 90548 7157 90557 7191
rect 90557 7157 90591 7191
rect 90591 7157 90600 7191
rect 90548 7148 90600 7157
rect 92296 7191 92348 7200
rect 92296 7157 92305 7191
rect 92305 7157 92339 7191
rect 92339 7157 92348 7191
rect 92296 7148 92348 7157
rect 96712 7148 96764 7200
rect 114836 7352 114888 7404
rect 187884 7352 187936 7404
rect 189172 7352 189224 7404
rect 208584 7352 208636 7404
rect 102232 7216 102284 7268
rect 113640 7216 113692 7268
rect 123484 7216 123536 7268
rect 218336 7216 218388 7268
rect 103244 7191 103296 7200
rect 103244 7157 103253 7191
rect 103253 7157 103287 7191
rect 103287 7157 103296 7191
rect 103244 7148 103296 7157
rect 113364 7191 113416 7200
rect 113364 7157 113373 7191
rect 113373 7157 113407 7191
rect 113407 7157 113416 7191
rect 113364 7148 113416 7157
rect 118516 7148 118568 7200
rect 226432 7148 226484 7200
rect 249524 7148 249576 7200
rect 251456 7395 251508 7404
rect 251456 7361 251465 7395
rect 251465 7361 251499 7395
rect 251499 7361 251508 7395
rect 251456 7352 251508 7361
rect 252468 7352 252520 7404
rect 253940 7352 253992 7404
rect 255228 7352 255280 7404
rect 256976 7352 257028 7404
rect 260840 7395 260892 7404
rect 260840 7361 260849 7395
rect 260849 7361 260883 7395
rect 260883 7361 260892 7395
rect 260840 7352 260892 7361
rect 262036 7352 262088 7404
rect 267096 7352 267148 7404
rect 270960 7395 271012 7404
rect 270960 7361 270969 7395
rect 270969 7361 271003 7395
rect 271003 7361 271012 7395
rect 270960 7352 271012 7361
rect 272156 7352 272208 7404
rect 364984 7352 365036 7404
rect 370688 7352 370740 7404
rect 252008 7327 252060 7336
rect 252008 7293 252017 7327
rect 252017 7293 252051 7327
rect 252051 7293 252060 7327
rect 252008 7284 252060 7293
rect 255780 7327 255832 7336
rect 255780 7293 255789 7327
rect 255789 7293 255823 7327
rect 255823 7293 255832 7327
rect 255780 7284 255832 7293
rect 264980 7284 265032 7336
rect 362040 7216 362092 7268
rect 66914 7046 66966 7098
rect 66978 7046 67030 7098
rect 67042 7046 67094 7098
rect 67106 7046 67158 7098
rect 67170 7046 67222 7098
rect 198842 7046 198894 7098
rect 198906 7046 198958 7098
rect 198970 7046 199022 7098
rect 199034 7046 199086 7098
rect 199098 7046 199150 7098
rect 330770 7046 330822 7098
rect 330834 7046 330886 7098
rect 330898 7046 330950 7098
rect 330962 7046 331014 7098
rect 331026 7046 331078 7098
rect 462698 7046 462750 7098
rect 462762 7046 462814 7098
rect 462826 7046 462878 7098
rect 462890 7046 462942 7098
rect 462954 7046 463006 7098
rect 46940 6944 46992 6996
rect 90548 6944 90600 6996
rect 94872 6944 94924 6996
rect 186688 6944 186740 6996
rect 262220 6944 262272 6996
rect 365260 6944 365312 6996
rect 78680 6876 78732 6928
rect 92296 6876 92348 6928
rect 94504 6876 94556 6928
rect 102232 6876 102284 6928
rect 125140 6876 125192 6928
rect 196716 6876 196768 6928
rect 202696 6876 202748 6928
rect 252008 6876 252060 6928
rect 360936 6876 360988 6928
rect 33140 6808 33192 6860
rect 92112 6783 92164 6792
rect 92112 6749 92121 6783
rect 92121 6749 92155 6783
rect 92155 6749 92164 6783
rect 92112 6740 92164 6749
rect 93768 6783 93820 6792
rect 93768 6749 93777 6783
rect 93777 6749 93811 6783
rect 93811 6749 93820 6783
rect 93768 6740 93820 6749
rect 94320 6740 94372 6792
rect 95148 6783 95200 6792
rect 95148 6749 95157 6783
rect 95157 6749 95191 6783
rect 95191 6749 95200 6783
rect 95148 6740 95200 6749
rect 96804 6740 96856 6792
rect 97448 6783 97500 6792
rect 97448 6749 97457 6783
rect 97457 6749 97491 6783
rect 97491 6749 97500 6783
rect 97448 6740 97500 6749
rect 100668 6672 100720 6724
rect 102876 6851 102928 6860
rect 102876 6817 102885 6851
rect 102885 6817 102919 6851
rect 102919 6817 102928 6851
rect 102876 6808 102928 6817
rect 104072 6851 104124 6860
rect 104072 6817 104081 6851
rect 104081 6817 104115 6851
rect 104115 6817 104124 6851
rect 104072 6808 104124 6817
rect 103244 6740 103296 6792
rect 104440 6740 104492 6792
rect 107292 6672 107344 6724
rect 109500 6808 109552 6860
rect 90916 6647 90968 6656
rect 90916 6613 90925 6647
rect 90925 6613 90959 6647
rect 90959 6613 90968 6647
rect 90916 6604 90968 6613
rect 92756 6647 92808 6656
rect 92756 6613 92765 6647
rect 92765 6613 92799 6647
rect 92799 6613 92808 6647
rect 92756 6604 92808 6613
rect 98368 6647 98420 6656
rect 98368 6613 98377 6647
rect 98377 6613 98411 6647
rect 98411 6613 98420 6647
rect 98368 6604 98420 6613
rect 101220 6647 101272 6656
rect 101220 6613 101229 6647
rect 101229 6613 101263 6647
rect 101263 6613 101272 6647
rect 101220 6604 101272 6613
rect 103704 6604 103756 6656
rect 110880 6715 110932 6724
rect 110880 6681 110889 6715
rect 110889 6681 110923 6715
rect 110923 6681 110932 6715
rect 110880 6672 110932 6681
rect 111524 6647 111576 6656
rect 111524 6613 111533 6647
rect 111533 6613 111567 6647
rect 111567 6613 111576 6647
rect 111524 6604 111576 6613
rect 112812 6851 112864 6860
rect 112812 6817 112821 6851
rect 112821 6817 112855 6851
rect 112855 6817 112864 6851
rect 112812 6808 112864 6817
rect 112720 6740 112772 6792
rect 113364 6740 113416 6792
rect 114652 6740 114704 6792
rect 114192 6715 114244 6724
rect 114192 6681 114201 6715
rect 114201 6681 114235 6715
rect 114235 6681 114244 6715
rect 114192 6672 114244 6681
rect 118792 6808 118844 6860
rect 224960 6808 225012 6860
rect 258356 6851 258408 6860
rect 258356 6817 258365 6851
rect 258365 6817 258399 6851
rect 258399 6817 258408 6851
rect 258356 6808 258408 6817
rect 268384 6808 268436 6860
rect 327540 6808 327592 6860
rect 377036 6808 377088 6860
rect 440976 6808 441028 6860
rect 444748 6808 444800 6860
rect 223212 6740 223264 6792
rect 225420 6672 225472 6724
rect 251364 6715 251416 6724
rect 251364 6681 251373 6715
rect 251373 6681 251407 6715
rect 251407 6681 251416 6715
rect 251364 6672 251416 6681
rect 256332 6740 256384 6792
rect 257528 6740 257580 6792
rect 259000 6783 259052 6792
rect 259000 6749 259009 6783
rect 259009 6749 259043 6783
rect 259043 6749 259052 6783
rect 259000 6740 259052 6749
rect 259920 6740 259972 6792
rect 116032 6604 116084 6656
rect 116676 6647 116728 6656
rect 116676 6613 116685 6647
rect 116685 6613 116719 6647
rect 116719 6613 116728 6647
rect 116676 6604 116728 6613
rect 120448 6604 120500 6656
rect 121644 6604 121696 6656
rect 122104 6604 122156 6656
rect 123392 6604 123444 6656
rect 124036 6604 124088 6656
rect 230480 6604 230532 6656
rect 252560 6647 252612 6656
rect 252560 6613 252569 6647
rect 252569 6613 252603 6647
rect 252603 6613 252612 6647
rect 252560 6604 252612 6613
rect 253940 6647 253992 6656
rect 253940 6613 253949 6647
rect 253949 6613 253983 6647
rect 253983 6613 253992 6647
rect 253940 6604 253992 6613
rect 254584 6647 254636 6656
rect 254584 6613 254593 6647
rect 254593 6613 254627 6647
rect 254627 6613 254636 6647
rect 254584 6604 254636 6613
rect 257160 6715 257212 6724
rect 257160 6681 257169 6715
rect 257169 6681 257203 6715
rect 257203 6681 257212 6715
rect 257160 6672 257212 6681
rect 267648 6740 267700 6792
rect 372804 6740 372856 6792
rect 401968 6740 402020 6792
rect 358820 6672 358872 6724
rect 361580 6672 361632 6724
rect 396080 6672 396132 6724
rect 432052 6672 432104 6724
rect 444012 6672 444064 6724
rect 365628 6604 365680 6656
rect 400312 6604 400364 6656
rect 408500 6604 408552 6656
rect 445024 6604 445076 6656
rect 67574 6502 67626 6554
rect 67638 6502 67690 6554
rect 67702 6502 67754 6554
rect 67766 6502 67818 6554
rect 67830 6502 67882 6554
rect 199502 6502 199554 6554
rect 199566 6502 199618 6554
rect 199630 6502 199682 6554
rect 199694 6502 199746 6554
rect 199758 6502 199810 6554
rect 331430 6502 331482 6554
rect 331494 6502 331546 6554
rect 331558 6502 331610 6554
rect 331622 6502 331674 6554
rect 331686 6502 331738 6554
rect 463358 6502 463410 6554
rect 463422 6502 463474 6554
rect 463486 6502 463538 6554
rect 463550 6502 463602 6554
rect 463614 6502 463666 6554
rect 40408 6400 40460 6452
rect 90916 6400 90968 6452
rect 62120 6332 62172 6384
rect 107292 6400 107344 6452
rect 17316 6264 17368 6316
rect 29920 6264 29972 6316
rect 12900 6196 12952 6248
rect 42984 6196 43036 6248
rect 1860 6128 1912 6180
rect 46940 6128 46992 6180
rect 68928 6128 68980 6180
rect 99932 6375 99984 6384
rect 99932 6341 99941 6375
rect 99941 6341 99975 6375
rect 99975 6341 99984 6375
rect 99932 6332 99984 6341
rect 101956 6375 102008 6384
rect 101956 6341 101965 6375
rect 101965 6341 101999 6375
rect 101999 6341 102008 6375
rect 101956 6332 102008 6341
rect 106188 6375 106240 6384
rect 106188 6341 106197 6375
rect 106197 6341 106231 6375
rect 106231 6341 106240 6375
rect 106188 6332 106240 6341
rect 100576 6264 100628 6316
rect 102600 6264 102652 6316
rect 103704 6196 103756 6248
rect 103796 6239 103848 6248
rect 103796 6205 103805 6239
rect 103805 6205 103839 6239
rect 103839 6205 103848 6239
rect 103796 6196 103848 6205
rect 42892 6060 42944 6112
rect 106924 6307 106976 6316
rect 106924 6273 106933 6307
rect 106933 6273 106967 6307
rect 106967 6273 106976 6307
rect 106924 6264 106976 6273
rect 113364 6400 113416 6452
rect 122104 6400 122156 6452
rect 131396 6400 131448 6452
rect 257160 6400 257212 6452
rect 262220 6400 262272 6452
rect 109776 6264 109828 6316
rect 111984 6264 112036 6316
rect 113180 6264 113232 6316
rect 113548 6307 113600 6316
rect 113548 6273 113557 6307
rect 113557 6273 113591 6307
rect 113591 6273 113600 6307
rect 113548 6264 113600 6273
rect 109500 6196 109552 6248
rect 114100 6239 114152 6248
rect 114100 6205 114109 6239
rect 114109 6205 114143 6239
rect 114143 6205 114152 6239
rect 114100 6196 114152 6205
rect 117504 6264 117556 6316
rect 120448 6307 120500 6316
rect 120448 6273 120457 6307
rect 120457 6273 120491 6307
rect 120491 6273 120500 6307
rect 120448 6264 120500 6273
rect 121000 6307 121052 6316
rect 121000 6273 121009 6307
rect 121009 6273 121043 6307
rect 121043 6273 121052 6307
rect 121000 6264 121052 6273
rect 121644 6307 121696 6316
rect 121644 6273 121653 6307
rect 121653 6273 121687 6307
rect 121687 6273 121696 6307
rect 121644 6264 121696 6273
rect 231860 6332 231912 6384
rect 362316 6400 362368 6452
rect 367928 6400 367980 6452
rect 397920 6400 397972 6452
rect 398840 6400 398892 6452
rect 440240 6400 440292 6452
rect 368480 6332 368532 6384
rect 369952 6332 370004 6384
rect 399852 6332 399904 6384
rect 400312 6332 400364 6384
rect 441712 6332 441764 6384
rect 442908 6332 442960 6384
rect 445852 6332 445904 6384
rect 123484 6264 123536 6316
rect 117964 6196 118016 6248
rect 118516 6239 118568 6248
rect 118516 6205 118525 6239
rect 118525 6205 118559 6239
rect 118559 6205 118568 6239
rect 118516 6196 118568 6205
rect 125140 6307 125192 6316
rect 125140 6273 125149 6307
rect 125149 6273 125183 6307
rect 125183 6273 125192 6307
rect 125140 6264 125192 6273
rect 125508 6307 125560 6316
rect 125508 6273 125517 6307
rect 125517 6273 125551 6307
rect 125551 6273 125560 6307
rect 125508 6264 125560 6273
rect 126612 6264 126664 6316
rect 127808 6307 127860 6316
rect 127808 6273 127817 6307
rect 127817 6273 127851 6307
rect 127851 6273 127860 6307
rect 127808 6264 127860 6273
rect 128360 6264 128412 6316
rect 131396 6264 131448 6316
rect 229836 6264 229888 6316
rect 260840 6264 260892 6316
rect 262312 6264 262364 6316
rect 264336 6264 264388 6316
rect 265992 6264 266044 6316
rect 123116 6128 123168 6180
rect 236276 6196 236328 6248
rect 262220 6196 262272 6248
rect 262404 6196 262456 6248
rect 124680 6128 124732 6180
rect 231400 6128 231452 6180
rect 367100 6264 367152 6316
rect 378140 6264 378192 6316
rect 442632 6264 442684 6316
rect 464528 6264 464580 6316
rect 482100 6264 482152 6316
rect 364984 6196 365036 6248
rect 381544 6196 381596 6248
rect 440700 6196 440752 6248
rect 459560 6196 459612 6248
rect 480260 6196 480312 6248
rect 369860 6128 369912 6180
rect 441620 6128 441672 6180
rect 445668 6128 445720 6180
rect 481272 6128 481324 6180
rect 94320 6103 94372 6112
rect 94320 6069 94329 6103
rect 94329 6069 94363 6103
rect 94363 6069 94372 6103
rect 94320 6060 94372 6069
rect 96804 6060 96856 6112
rect 99564 6060 99616 6112
rect 100576 6060 100628 6112
rect 102600 6103 102652 6112
rect 102600 6069 102609 6103
rect 102609 6069 102643 6103
rect 102643 6069 102652 6103
rect 102600 6060 102652 6069
rect 104440 6103 104492 6112
rect 104440 6069 104449 6103
rect 104449 6069 104483 6103
rect 104483 6069 104492 6103
rect 104440 6060 104492 6069
rect 105084 6103 105136 6112
rect 105084 6069 105093 6103
rect 105093 6069 105127 6103
rect 105127 6069 105136 6103
rect 105084 6060 105136 6069
rect 109776 6103 109828 6112
rect 109776 6069 109785 6103
rect 109785 6069 109819 6103
rect 109819 6069 109828 6103
rect 109776 6060 109828 6069
rect 111984 6060 112036 6112
rect 114652 6060 114704 6112
rect 117504 6060 117556 6112
rect 123208 6103 123260 6112
rect 123208 6069 123217 6103
rect 123217 6069 123251 6103
rect 123251 6069 123260 6103
rect 123208 6060 123260 6069
rect 126612 6103 126664 6112
rect 126612 6069 126621 6103
rect 126621 6069 126655 6103
rect 126655 6069 126664 6103
rect 126612 6060 126664 6069
rect 131764 6060 131816 6112
rect 134432 6060 134484 6112
rect 241612 6060 241664 6112
rect 256332 6103 256384 6112
rect 256332 6069 256341 6103
rect 256341 6069 256375 6103
rect 256375 6069 256384 6103
rect 256332 6060 256384 6069
rect 257528 6103 257580 6112
rect 257528 6069 257537 6103
rect 257537 6069 257571 6103
rect 257571 6069 257580 6103
rect 257528 6060 257580 6069
rect 259000 6103 259052 6112
rect 259000 6069 259009 6103
rect 259009 6069 259043 6103
rect 259043 6069 259052 6103
rect 259000 6060 259052 6069
rect 259920 6103 259972 6112
rect 259920 6069 259929 6103
rect 259929 6069 259963 6103
rect 259963 6069 259972 6103
rect 259920 6060 259972 6069
rect 260840 6103 260892 6112
rect 260840 6069 260849 6103
rect 260849 6069 260883 6103
rect 260883 6069 260892 6103
rect 260840 6060 260892 6069
rect 264336 6103 264388 6112
rect 264336 6069 264345 6103
rect 264345 6069 264379 6103
rect 264379 6069 264388 6103
rect 264336 6060 264388 6069
rect 66914 5958 66966 6010
rect 66978 5958 67030 6010
rect 67042 5958 67094 6010
rect 67106 5958 67158 6010
rect 67170 5958 67222 6010
rect 198842 5958 198894 6010
rect 198906 5958 198958 6010
rect 198970 5958 199022 6010
rect 199034 5958 199086 6010
rect 199098 5958 199150 6010
rect 330770 5958 330822 6010
rect 330834 5958 330886 6010
rect 330898 5958 330950 6010
rect 330962 5958 331014 6010
rect 331026 5958 331078 6010
rect 462698 5958 462750 6010
rect 462762 5958 462814 6010
rect 462826 5958 462878 6010
rect 462890 5958 462942 6010
rect 462954 5958 463006 6010
rect 48780 5856 48832 5908
rect 102600 5856 102652 5908
rect 75920 5788 75972 5840
rect 111524 5856 111576 5908
rect 114100 5856 114152 5908
rect 123300 5856 123352 5908
rect 127348 5856 127400 5908
rect 103796 5788 103848 5840
rect 19892 5720 19944 5772
rect 98368 5720 98420 5772
rect 107568 5763 107620 5772
rect 107568 5729 107577 5763
rect 107577 5729 107611 5763
rect 107611 5729 107620 5763
rect 107568 5720 107620 5729
rect 110880 5788 110932 5840
rect 120172 5788 120224 5840
rect 115388 5720 115440 5772
rect 98644 5652 98696 5704
rect 47400 5584 47452 5636
rect 106924 5584 106976 5636
rect 56508 5516 56560 5568
rect 105084 5516 105136 5568
rect 107660 5516 107712 5568
rect 109868 5695 109920 5704
rect 109868 5661 109877 5695
rect 109877 5661 109911 5695
rect 109911 5661 109920 5695
rect 109868 5652 109920 5661
rect 117136 5652 117188 5704
rect 118792 5652 118844 5704
rect 108764 5516 108816 5568
rect 113548 5516 113600 5568
rect 115480 5559 115532 5568
rect 115480 5525 115489 5559
rect 115489 5525 115523 5559
rect 115523 5525 115532 5559
rect 115480 5516 115532 5525
rect 118884 5559 118936 5568
rect 118884 5525 118893 5559
rect 118893 5525 118927 5559
rect 118927 5525 118936 5559
rect 118884 5516 118936 5525
rect 120724 5695 120776 5704
rect 120724 5661 120733 5695
rect 120733 5661 120767 5695
rect 120767 5661 120776 5695
rect 120724 5652 120776 5661
rect 122840 5652 122892 5704
rect 124036 5652 124088 5704
rect 124128 5695 124180 5704
rect 124128 5661 124137 5695
rect 124137 5661 124171 5695
rect 124171 5661 124180 5695
rect 124128 5652 124180 5661
rect 124680 5763 124732 5772
rect 124680 5729 124689 5763
rect 124689 5729 124723 5763
rect 124723 5729 124732 5763
rect 124680 5720 124732 5729
rect 127348 5652 127400 5704
rect 130660 5695 130712 5704
rect 130660 5661 130669 5695
rect 130669 5661 130703 5695
rect 130703 5661 130712 5695
rect 130660 5652 130712 5661
rect 130936 5695 130988 5704
rect 130936 5661 130945 5695
rect 130945 5661 130979 5695
rect 130979 5661 130988 5695
rect 130936 5652 130988 5661
rect 131764 5695 131816 5704
rect 131764 5661 131773 5695
rect 131773 5661 131807 5695
rect 131807 5661 131816 5695
rect 131764 5652 131816 5661
rect 132040 5695 132092 5704
rect 132040 5661 132049 5695
rect 132049 5661 132083 5695
rect 132083 5661 132092 5695
rect 132040 5652 132092 5661
rect 134432 5695 134484 5704
rect 134432 5661 134441 5695
rect 134441 5661 134475 5695
rect 134475 5661 134484 5695
rect 134432 5652 134484 5661
rect 135352 5652 135404 5704
rect 135536 5763 135588 5772
rect 135536 5729 135545 5763
rect 135545 5729 135579 5763
rect 135579 5729 135588 5763
rect 135536 5720 135588 5729
rect 149704 5856 149756 5908
rect 228088 5788 228140 5840
rect 149704 5720 149756 5772
rect 226984 5720 227036 5772
rect 372528 5856 372580 5908
rect 138296 5652 138348 5704
rect 139032 5627 139084 5636
rect 139032 5593 139041 5627
rect 139041 5593 139075 5627
rect 139075 5593 139084 5627
rect 139032 5584 139084 5593
rect 263140 5652 263192 5704
rect 223764 5584 223816 5636
rect 252652 5584 252704 5636
rect 268384 5652 268436 5704
rect 365720 5788 365772 5840
rect 269672 5652 269724 5704
rect 370780 5720 370832 5772
rect 373448 5584 373500 5636
rect 128176 5559 128228 5568
rect 128176 5525 128185 5559
rect 128185 5525 128219 5559
rect 128219 5525 128228 5559
rect 128176 5516 128228 5525
rect 130108 5559 130160 5568
rect 130108 5525 130117 5559
rect 130117 5525 130151 5559
rect 130151 5525 130160 5559
rect 130108 5516 130160 5525
rect 130660 5516 130712 5568
rect 133604 5559 133656 5568
rect 133604 5525 133613 5559
rect 133613 5525 133647 5559
rect 133647 5525 133656 5559
rect 133604 5516 133656 5525
rect 138204 5559 138256 5568
rect 138204 5525 138213 5559
rect 138213 5525 138247 5559
rect 138247 5525 138256 5559
rect 138204 5516 138256 5525
rect 141700 5516 141752 5568
rect 262312 5559 262364 5568
rect 262312 5525 262321 5559
rect 262321 5525 262355 5559
rect 262355 5525 262364 5559
rect 262312 5516 262364 5525
rect 263140 5559 263192 5568
rect 263140 5525 263149 5559
rect 263149 5525 263183 5559
rect 263183 5525 263192 5559
rect 263140 5516 263192 5525
rect 265992 5559 266044 5568
rect 265992 5525 266001 5559
rect 266001 5525 266035 5559
rect 266035 5525 266044 5559
rect 265992 5516 266044 5525
rect 67574 5414 67626 5466
rect 67638 5414 67690 5466
rect 67702 5414 67754 5466
rect 67766 5414 67818 5466
rect 67830 5414 67882 5466
rect 199502 5414 199554 5466
rect 199566 5414 199618 5466
rect 199630 5414 199682 5466
rect 199694 5414 199746 5466
rect 199758 5414 199810 5466
rect 331430 5414 331482 5466
rect 331494 5414 331546 5466
rect 331558 5414 331610 5466
rect 331622 5414 331674 5466
rect 331686 5414 331738 5466
rect 463358 5414 463410 5466
rect 463422 5414 463474 5466
rect 463486 5414 463538 5466
rect 463550 5414 463602 5466
rect 463614 5414 463666 5466
rect 18052 5312 18104 5364
rect 96620 5312 96672 5364
rect 9588 5244 9640 5296
rect 92388 5244 92440 5296
rect 5172 5176 5224 5228
rect 94504 5176 94556 5228
rect 115112 5176 115164 5228
rect 125692 5176 125744 5228
rect 127624 5176 127676 5228
rect 6828 5108 6880 5160
rect 78680 5108 78732 5160
rect 82820 5108 82872 5160
rect 117136 5151 117188 5160
rect 117136 5117 117145 5151
rect 117145 5117 117179 5151
rect 117179 5117 117188 5151
rect 117136 5108 117188 5117
rect 128084 5151 128136 5160
rect 128084 5117 128093 5151
rect 128093 5117 128127 5151
rect 128127 5117 128136 5151
rect 128084 5108 128136 5117
rect 68836 5040 68888 5092
rect 45652 4972 45704 5024
rect 68928 4972 68980 5024
rect 76564 5040 76616 5092
rect 124128 5040 124180 5092
rect 131212 5176 131264 5228
rect 132684 5176 132736 5228
rect 130844 5151 130896 5160
rect 130844 5117 130853 5151
rect 130853 5117 130887 5151
rect 130887 5117 130896 5151
rect 130844 5108 130896 5117
rect 133512 5151 133564 5160
rect 133512 5117 133521 5151
rect 133521 5117 133555 5151
rect 133555 5117 133564 5151
rect 133512 5108 133564 5117
rect 134340 5219 134392 5228
rect 134340 5185 134349 5219
rect 134349 5185 134383 5219
rect 134383 5185 134392 5219
rect 134340 5176 134392 5185
rect 241152 5312 241204 5364
rect 252560 5312 252612 5364
rect 360752 5312 360804 5364
rect 389180 5312 389232 5364
rect 403624 5312 403676 5364
rect 426992 5312 427044 5364
rect 443092 5312 443144 5364
rect 443736 5312 443788 5364
rect 446128 5312 446180 5364
rect 477500 5312 477552 5364
rect 481640 5312 481692 5364
rect 137008 5244 137060 5296
rect 137100 5176 137152 5228
rect 140504 5176 140556 5228
rect 141332 5219 141384 5228
rect 141332 5185 141341 5219
rect 141341 5185 141375 5219
rect 141375 5185 141384 5219
rect 141332 5176 141384 5185
rect 141700 5176 141752 5228
rect 144552 5219 144604 5228
rect 144552 5185 144561 5219
rect 144561 5185 144595 5219
rect 144595 5185 144604 5219
rect 144552 5176 144604 5185
rect 137836 5151 137888 5160
rect 137836 5117 137845 5151
rect 137845 5117 137879 5151
rect 137879 5117 137888 5151
rect 137836 5108 137888 5117
rect 142436 5151 142488 5160
rect 142436 5117 142445 5151
rect 142445 5117 142479 5151
rect 142479 5117 142488 5151
rect 142436 5108 142488 5117
rect 144828 5151 144880 5160
rect 144828 5117 144837 5151
rect 144837 5117 144871 5151
rect 144871 5117 144880 5151
rect 144828 5108 144880 5117
rect 145840 5244 145892 5296
rect 236920 5244 236972 5296
rect 291108 5244 291160 5296
rect 391940 5244 391992 5296
rect 417056 5244 417108 5296
rect 443184 5244 443236 5296
rect 145472 5176 145524 5228
rect 145932 5219 145984 5228
rect 145932 5185 145941 5219
rect 145941 5185 145975 5219
rect 145975 5185 145984 5219
rect 145932 5176 145984 5185
rect 148048 5219 148100 5228
rect 148048 5185 148057 5219
rect 148057 5185 148091 5219
rect 148091 5185 148100 5219
rect 148048 5176 148100 5185
rect 148968 5108 149020 5160
rect 270592 5176 270644 5228
rect 285956 5176 286008 5228
rect 390560 5176 390612 5228
rect 403992 5176 404044 5228
rect 443000 5176 443052 5228
rect 233608 5108 233660 5160
rect 271696 5151 271748 5160
rect 271696 5117 271705 5151
rect 271705 5117 271739 5151
rect 271739 5117 271748 5151
rect 271696 5108 271748 5117
rect 288532 5108 288584 5160
rect 391388 5108 391440 5160
rect 400404 5108 400456 5160
rect 441804 5108 441856 5160
rect 475292 5108 475344 5160
rect 480720 5108 480772 5160
rect 481732 5108 481784 5160
rect 482008 5108 482060 5160
rect 237932 5040 237984 5092
rect 283380 5040 283432 5092
rect 390652 5040 390704 5092
rect 404360 5040 404412 5092
rect 439136 5040 439188 5092
rect 120724 4972 120776 5024
rect 122840 4972 122892 5024
rect 125692 5015 125744 5024
rect 125692 4981 125701 5015
rect 125701 4981 125735 5015
rect 125735 4981 125744 5015
rect 125692 4972 125744 4981
rect 129556 5015 129608 5024
rect 129556 4981 129565 5015
rect 129565 4981 129599 5015
rect 129599 4981 129608 5015
rect 129556 4972 129608 4981
rect 132684 5015 132736 5024
rect 132684 4981 132693 5015
rect 132693 4981 132727 5015
rect 132727 4981 132736 5015
rect 132684 4972 132736 4981
rect 135352 5015 135404 5024
rect 135352 4981 135361 5015
rect 135361 4981 135395 5015
rect 135395 4981 135404 5015
rect 135352 4972 135404 4981
rect 137008 5015 137060 5024
rect 137008 4981 137017 5015
rect 137017 4981 137051 5015
rect 137051 4981 137060 5015
rect 137008 4972 137060 4981
rect 137100 4972 137152 5024
rect 140504 5015 140556 5024
rect 140504 4981 140513 5015
rect 140513 4981 140547 5015
rect 140547 4981 140556 5015
rect 140504 4972 140556 4981
rect 140688 4972 140740 5024
rect 144552 4972 144604 5024
rect 144644 4972 144696 5024
rect 148048 4972 148100 5024
rect 268384 5015 268436 5024
rect 268384 4981 268393 5015
rect 268393 4981 268427 5015
rect 268427 4981 268436 5015
rect 268384 4972 268436 4981
rect 269672 5015 269724 5024
rect 269672 4981 269681 5015
rect 269681 4981 269715 5015
rect 269715 4981 269724 5015
rect 269672 4972 269724 4981
rect 270592 5015 270644 5024
rect 270592 4981 270601 5015
rect 270601 4981 270635 5015
rect 270635 4981 270644 5015
rect 270592 4972 270644 4981
rect 360660 4972 360712 5024
rect 440332 5040 440384 5092
rect 440148 4972 440200 5024
rect 444564 4972 444616 5024
rect 456800 4972 456852 5024
rect 478880 4972 478932 5024
rect 66914 4870 66966 4922
rect 66978 4870 67030 4922
rect 67042 4870 67094 4922
rect 67106 4870 67158 4922
rect 67170 4870 67222 4922
rect 198842 4870 198894 4922
rect 198906 4870 198958 4922
rect 198970 4870 199022 4922
rect 199034 4870 199086 4922
rect 199098 4870 199150 4922
rect 330770 4870 330822 4922
rect 330834 4870 330886 4922
rect 330898 4870 330950 4922
rect 330962 4870 331014 4922
rect 331026 4870 331078 4922
rect 462698 4870 462750 4922
rect 462762 4870 462814 4922
rect 462826 4870 462878 4922
rect 462890 4870 462942 4922
rect 462954 4870 463006 4922
rect 12164 4768 12216 4820
rect 63500 4768 63552 4820
rect 73988 4768 74040 4820
rect 122840 4768 122892 4820
rect 123392 4768 123444 4820
rect 128176 4768 128228 4820
rect 130844 4768 130896 4820
rect 59176 4700 59228 4752
rect 94320 4700 94372 4752
rect 97172 4700 97224 4752
rect 132684 4700 132736 4752
rect 79232 4632 79284 4684
rect 92756 4632 92808 4684
rect 94136 4632 94188 4684
rect 129556 4632 129608 4684
rect 130384 4632 130436 4684
rect 135352 4700 135404 4752
rect 138112 4768 138164 4820
rect 243360 4768 243412 4820
rect 280804 4768 280856 4820
rect 389824 4768 389876 4820
rect 390560 4768 390612 4820
rect 438860 4768 438912 4820
rect 439136 4768 439188 4820
rect 445760 4768 445812 4820
rect 450820 4768 450872 4820
rect 481916 4768 481968 4820
rect 488448 4768 488500 4820
rect 511632 4768 511684 4820
rect 23204 4564 23256 4616
rect 96712 4564 96764 4616
rect 112628 4564 112680 4616
rect 130844 4564 130896 4616
rect 131028 4564 131080 4616
rect 91560 4496 91612 4548
rect 123392 4496 123444 4548
rect 102324 4428 102376 4480
rect 130384 4496 130436 4548
rect 131212 4539 131264 4548
rect 131212 4505 131221 4539
rect 131221 4505 131255 4539
rect 131255 4505 131264 4539
rect 131212 4496 131264 4505
rect 138112 4632 138164 4684
rect 141608 4700 141660 4752
rect 247684 4700 247736 4752
rect 293684 4700 293736 4752
rect 392492 4700 392544 4752
rect 137928 4607 137980 4616
rect 137928 4573 137937 4607
rect 137937 4573 137971 4607
rect 137971 4573 137980 4607
rect 137928 4564 137980 4573
rect 127624 4471 127676 4480
rect 127624 4437 127633 4471
rect 127633 4437 127667 4471
rect 127667 4437 127676 4471
rect 127624 4428 127676 4437
rect 127716 4428 127768 4480
rect 134340 4428 134392 4480
rect 136180 4471 136232 4480
rect 136180 4437 136189 4471
rect 136189 4437 136223 4471
rect 136223 4437 136232 4471
rect 136180 4428 136232 4437
rect 145840 4632 145892 4684
rect 141056 4564 141108 4616
rect 246672 4632 246724 4684
rect 271696 4632 271748 4684
rect 293868 4632 293920 4684
rect 309140 4632 309192 4684
rect 395528 4632 395580 4684
rect 149152 4607 149204 4616
rect 149152 4573 149161 4607
rect 149161 4573 149195 4607
rect 149195 4573 149204 4607
rect 149152 4564 149204 4573
rect 255872 4564 255924 4616
rect 322020 4564 322072 4616
rect 398472 4564 398524 4616
rect 141608 4539 141660 4548
rect 141608 4505 141617 4539
rect 141617 4505 141651 4539
rect 141651 4505 141660 4539
rect 141608 4496 141660 4505
rect 244464 4496 244516 4548
rect 244832 4496 244884 4548
rect 312912 4496 312964 4548
rect 334900 4496 334952 4548
rect 361488 4496 361540 4548
rect 145472 4471 145524 4480
rect 145472 4437 145481 4471
rect 145481 4437 145515 4471
rect 145515 4437 145524 4471
rect 145472 4428 145524 4437
rect 249892 4428 249944 4480
rect 357072 4428 357124 4480
rect 67574 4326 67626 4378
rect 67638 4326 67690 4378
rect 67702 4326 67754 4378
rect 67766 4326 67818 4378
rect 67830 4326 67882 4378
rect 199502 4326 199554 4378
rect 199566 4326 199618 4378
rect 199630 4326 199682 4378
rect 199694 4326 199746 4378
rect 199758 4326 199810 4378
rect 331430 4326 331482 4378
rect 331494 4326 331546 4378
rect 331558 4326 331610 4378
rect 331622 4326 331674 4378
rect 331686 4326 331738 4378
rect 463358 4326 463410 4378
rect 463422 4326 463474 4378
rect 463486 4326 463538 4378
rect 463550 4326 463602 4378
rect 463614 4326 463666 4378
rect 109960 4224 110012 4276
rect 138204 4224 138256 4276
rect 142436 4224 142488 4276
rect 249340 4224 249392 4276
rect 128084 4156 128136 4208
rect 234712 4156 234764 4208
rect 84292 4088 84344 4140
rect 126612 4088 126664 4140
rect 126888 4088 126940 4140
rect 137928 4088 137980 4140
rect 48228 4020 48280 4072
rect 75920 4020 75972 4072
rect 79048 4020 79100 4072
rect 125140 4020 125192 4072
rect 133052 4020 133104 4072
rect 141700 4088 141752 4140
rect 144000 4063 144052 4072
rect 144000 4029 144009 4063
rect 144009 4029 144043 4063
rect 144043 4029 144052 4063
rect 144000 4020 144052 4029
rect 4436 3952 4488 4004
rect 71044 3952 71096 4004
rect 76472 3952 76524 4004
rect 123208 3952 123260 4004
rect 130844 3952 130896 4004
rect 71412 3884 71464 3936
rect 121644 3884 121696 3936
rect 122932 3884 122984 3936
rect 133144 3884 133196 3936
rect 143172 3995 143224 4004
rect 143172 3961 143181 3995
rect 143181 3961 143215 3995
rect 143215 3961 143224 3995
rect 143172 3952 143224 3961
rect 140964 3884 141016 3936
rect 141056 3884 141108 3936
rect 141700 3884 141752 3936
rect 144736 3952 144788 4004
rect 148140 4088 148192 4140
rect 148692 4063 148744 4072
rect 148692 4029 148701 4063
rect 148701 4029 148735 4063
rect 148735 4029 148744 4063
rect 148692 4020 148744 4029
rect 150808 4131 150860 4140
rect 150808 4097 150817 4131
rect 150817 4097 150851 4131
rect 150851 4097 150860 4131
rect 150808 4088 150860 4097
rect 150900 4020 150952 4072
rect 205364 4088 205416 4140
rect 210424 4088 210476 4140
rect 301412 4088 301464 4140
rect 375380 4088 375432 4140
rect 440240 4088 440292 4140
rect 445300 4088 445352 4140
rect 251272 4020 251324 4072
rect 298836 4020 298888 4072
rect 374276 4020 374328 4072
rect 378692 4020 378744 4072
rect 403072 4020 403124 4072
rect 151176 3952 151228 4004
rect 253112 3952 253164 4004
rect 319260 3952 319312 4004
rect 397460 3952 397512 4004
rect 256424 3884 256476 3936
rect 355508 3884 355560 3936
rect 440424 3884 440476 3936
rect 66914 3782 66966 3834
rect 66978 3782 67030 3834
rect 67042 3782 67094 3834
rect 67106 3782 67158 3834
rect 67170 3782 67222 3834
rect 198842 3782 198894 3834
rect 198906 3782 198958 3834
rect 198970 3782 199022 3834
rect 199034 3782 199086 3834
rect 199098 3782 199150 3834
rect 330770 3782 330822 3834
rect 330834 3782 330886 3834
rect 330898 3782 330950 3834
rect 330962 3782 331014 3834
rect 331026 3782 331078 3834
rect 462698 3782 462750 3834
rect 462762 3782 462814 3834
rect 462826 3782 462878 3834
rect 462890 3782 462942 3834
rect 462954 3782 463006 3834
rect 1860 3723 1912 3732
rect 1860 3689 1869 3723
rect 1869 3689 1903 3723
rect 1903 3689 1912 3723
rect 1860 3680 1912 3689
rect 4436 3723 4488 3732
rect 4436 3689 4445 3723
rect 4445 3689 4479 3723
rect 4479 3689 4488 3723
rect 4436 3680 4488 3689
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 9588 3723 9640 3732
rect 9588 3689 9597 3723
rect 9597 3689 9631 3723
rect 9631 3689 9640 3723
rect 9588 3680 9640 3689
rect 12164 3723 12216 3732
rect 12164 3689 12173 3723
rect 12173 3689 12207 3723
rect 12207 3689 12216 3723
rect 12164 3680 12216 3689
rect 14740 3723 14792 3732
rect 14740 3689 14749 3723
rect 14749 3689 14783 3723
rect 14783 3689 14792 3723
rect 14740 3680 14792 3689
rect 17316 3723 17368 3732
rect 17316 3689 17325 3723
rect 17325 3689 17359 3723
rect 17359 3689 17368 3723
rect 17316 3680 17368 3689
rect 19892 3723 19944 3732
rect 19892 3689 19901 3723
rect 19901 3689 19935 3723
rect 19935 3689 19944 3723
rect 19892 3680 19944 3689
rect 22468 3723 22520 3732
rect 22468 3689 22477 3723
rect 22477 3689 22511 3723
rect 22511 3689 22520 3723
rect 22468 3680 22520 3689
rect 33140 3680 33192 3732
rect 36084 3723 36136 3732
rect 36084 3689 36093 3723
rect 36093 3689 36127 3723
rect 36127 3689 36136 3723
rect 36084 3680 36136 3689
rect 43812 3723 43864 3732
rect 43812 3689 43821 3723
rect 43821 3689 43855 3723
rect 43855 3689 43864 3723
rect 43812 3680 43864 3689
rect 45652 3723 45704 3732
rect 45652 3689 45661 3723
rect 45661 3689 45695 3723
rect 45695 3689 45704 3723
rect 45652 3680 45704 3689
rect 48228 3723 48280 3732
rect 48228 3689 48237 3723
rect 48237 3689 48271 3723
rect 48271 3689 48280 3723
rect 48228 3680 48280 3689
rect 59268 3723 59320 3732
rect 59268 3689 59277 3723
rect 59277 3689 59311 3723
rect 59311 3689 59320 3723
rect 59268 3680 59320 3689
rect 31852 3612 31904 3664
rect 62120 3680 62172 3732
rect 63500 3680 63552 3732
rect 67272 3680 67324 3732
rect 120448 3680 120500 3732
rect 122932 3723 122984 3732
rect 122932 3689 122941 3723
rect 122941 3689 122975 3723
rect 122975 3689 122984 3723
rect 122932 3680 122984 3689
rect 130844 3723 130896 3732
rect 130844 3689 130853 3723
rect 130853 3689 130887 3723
rect 130887 3689 130896 3723
rect 130844 3680 130896 3689
rect 133144 3680 133196 3732
rect 140688 3680 140740 3732
rect 140964 3680 141016 3732
rect 144644 3680 144696 3732
rect 148692 3680 148744 3732
rect 194692 3680 194744 3732
rect 194784 3680 194836 3732
rect 35900 3544 35952 3596
rect 47400 3544 47452 3596
rect 109684 3544 109736 3596
rect 109960 3655 110012 3664
rect 109960 3621 109969 3655
rect 109969 3621 110003 3655
rect 110003 3621 110012 3655
rect 109960 3612 110012 3621
rect 115112 3655 115164 3664
rect 115112 3621 115121 3655
rect 115121 3621 115155 3655
rect 115155 3621 115164 3655
rect 115112 3612 115164 3621
rect 111064 3544 111116 3596
rect 29368 3476 29420 3528
rect 36084 3476 36136 3528
rect 40684 3519 40736 3528
rect 40684 3485 40693 3519
rect 40693 3485 40727 3519
rect 40727 3485 40736 3519
rect 40684 3476 40736 3485
rect 43812 3476 43864 3528
rect 45836 3519 45888 3528
rect 45836 3485 45845 3519
rect 45845 3485 45879 3519
rect 45879 3485 45888 3519
rect 45836 3476 45888 3485
rect 1308 3408 1360 3460
rect 3976 3408 4028 3460
rect 6184 3383 6236 3392
rect 6184 3349 6193 3383
rect 6193 3349 6227 3383
rect 6227 3349 6236 3383
rect 9128 3408 9180 3460
rect 6184 3340 6236 3349
rect 11336 3383 11388 3392
rect 11336 3349 11345 3383
rect 11345 3349 11379 3383
rect 11379 3349 11388 3383
rect 14280 3408 14332 3460
rect 19248 3408 19300 3460
rect 11336 3340 11388 3349
rect 16580 3383 16632 3392
rect 16580 3349 16589 3383
rect 16589 3349 16623 3383
rect 16623 3349 16632 3383
rect 16580 3340 16632 3349
rect 21640 3383 21692 3392
rect 21640 3349 21649 3383
rect 21649 3349 21683 3383
rect 21683 3349 21692 3383
rect 24584 3408 24636 3460
rect 21640 3340 21692 3349
rect 24860 3340 24912 3392
rect 28908 3408 28960 3460
rect 33140 3408 33192 3460
rect 27620 3383 27672 3392
rect 27620 3349 27629 3383
rect 27629 3349 27663 3383
rect 27663 3349 27672 3383
rect 27620 3340 27672 3349
rect 32772 3383 32824 3392
rect 32772 3349 32781 3383
rect 32781 3349 32815 3383
rect 32815 3349 32824 3383
rect 32772 3340 32824 3349
rect 39120 3340 39172 3392
rect 43168 3340 43220 3392
rect 55128 3476 55180 3528
rect 59268 3476 59320 3528
rect 60648 3476 60700 3528
rect 49700 3340 49752 3392
rect 51540 3383 51592 3392
rect 51540 3349 51549 3383
rect 51549 3349 51583 3383
rect 51583 3349 51592 3383
rect 51540 3340 51592 3349
rect 52736 3383 52788 3392
rect 52736 3349 52745 3383
rect 52745 3349 52779 3383
rect 52779 3349 52788 3383
rect 52736 3340 52788 3349
rect 62948 3408 63000 3460
rect 55956 3383 56008 3392
rect 55956 3349 55965 3383
rect 55965 3349 55999 3383
rect 55999 3349 56008 3383
rect 55956 3340 56008 3349
rect 56692 3340 56744 3392
rect 60740 3340 60792 3392
rect 67272 3476 67324 3528
rect 69020 3519 69072 3528
rect 69020 3485 69029 3519
rect 69029 3485 69063 3519
rect 69063 3485 69072 3519
rect 69020 3476 69072 3485
rect 71228 3476 71280 3528
rect 74724 3519 74776 3528
rect 74724 3485 74733 3519
rect 74733 3485 74767 3519
rect 74767 3485 74776 3519
rect 74724 3476 74776 3485
rect 63132 3408 63184 3460
rect 76472 3451 76524 3460
rect 76472 3417 76481 3451
rect 76481 3417 76515 3451
rect 76515 3417 76524 3451
rect 76472 3408 76524 3417
rect 76656 3451 76708 3460
rect 76656 3417 76665 3451
rect 76665 3417 76699 3451
rect 76699 3417 76708 3451
rect 76656 3408 76708 3417
rect 79048 3451 79100 3460
rect 79048 3417 79057 3451
rect 79057 3417 79091 3451
rect 79091 3417 79100 3451
rect 79048 3408 79100 3417
rect 81900 3519 81952 3528
rect 81900 3485 81909 3519
rect 81909 3485 81943 3519
rect 81943 3485 81952 3519
rect 81900 3476 81952 3485
rect 64880 3340 64932 3392
rect 69020 3340 69072 3392
rect 71412 3383 71464 3392
rect 71412 3349 71421 3383
rect 71421 3349 71455 3383
rect 71455 3349 71464 3383
rect 71412 3340 71464 3349
rect 71504 3340 71556 3392
rect 78496 3383 78548 3392
rect 78496 3349 78505 3383
rect 78505 3349 78539 3383
rect 78539 3349 78548 3383
rect 82452 3451 82504 3460
rect 82452 3417 82461 3451
rect 82461 3417 82495 3451
rect 82495 3417 82504 3451
rect 82452 3408 82504 3417
rect 78496 3340 78548 3349
rect 81532 3340 81584 3392
rect 81900 3340 81952 3392
rect 83648 3383 83700 3392
rect 83648 3349 83657 3383
rect 83657 3349 83691 3383
rect 83691 3349 83700 3383
rect 86960 3451 87012 3460
rect 86960 3417 86969 3451
rect 86969 3417 87003 3451
rect 87003 3417 87012 3451
rect 86960 3408 87012 3417
rect 89628 3519 89680 3528
rect 89628 3485 89637 3519
rect 89637 3485 89671 3519
rect 89671 3485 89680 3519
rect 89628 3476 89680 3485
rect 89720 3476 89772 3528
rect 90180 3519 90232 3528
rect 90180 3485 90189 3519
rect 90189 3485 90223 3519
rect 90223 3485 90232 3519
rect 90180 3476 90232 3485
rect 92112 3451 92164 3460
rect 92112 3417 92121 3451
rect 92121 3417 92155 3451
rect 92155 3417 92164 3451
rect 92112 3408 92164 3417
rect 83648 3340 83700 3349
rect 84292 3383 84344 3392
rect 84292 3349 84301 3383
rect 84301 3349 84335 3383
rect 84335 3349 84344 3383
rect 84292 3340 84344 3349
rect 86868 3383 86920 3392
rect 86868 3349 86877 3383
rect 86877 3349 86911 3383
rect 86911 3349 86920 3383
rect 86868 3340 86920 3349
rect 87420 3340 87472 3392
rect 92020 3383 92072 3392
rect 92020 3349 92029 3383
rect 92029 3349 92063 3383
rect 92063 3349 92072 3383
rect 92020 3340 92072 3349
rect 92572 3340 92624 3392
rect 97908 3476 97960 3528
rect 94596 3383 94648 3392
rect 94596 3349 94605 3383
rect 94605 3349 94639 3383
rect 94639 3349 94648 3383
rect 94596 3340 94648 3349
rect 94780 3340 94832 3392
rect 97908 3383 97960 3392
rect 97908 3349 97917 3383
rect 97917 3349 97951 3383
rect 97951 3349 97960 3383
rect 97908 3340 97960 3349
rect 99104 3383 99156 3392
rect 99104 3349 99113 3383
rect 99113 3349 99147 3383
rect 99147 3349 99156 3383
rect 102140 3408 102192 3460
rect 105084 3519 105136 3528
rect 105084 3485 105093 3519
rect 105093 3485 105127 3519
rect 105127 3485 105136 3519
rect 105084 3476 105136 3485
rect 112720 3476 112772 3528
rect 105636 3451 105688 3460
rect 105636 3417 105645 3451
rect 105645 3417 105679 3451
rect 105679 3417 105688 3451
rect 105636 3408 105688 3417
rect 107568 3451 107620 3460
rect 107568 3417 107577 3451
rect 107577 3417 107611 3451
rect 107611 3417 107620 3451
rect 107568 3408 107620 3417
rect 99104 3340 99156 3349
rect 99748 3383 99800 3392
rect 99748 3349 99757 3383
rect 99757 3349 99791 3383
rect 99791 3349 99800 3383
rect 99748 3340 99800 3349
rect 102324 3383 102376 3392
rect 102324 3349 102333 3383
rect 102333 3349 102367 3383
rect 102367 3349 102376 3383
rect 102324 3340 102376 3349
rect 102508 3340 102560 3392
rect 107476 3383 107528 3392
rect 107476 3349 107485 3383
rect 107485 3349 107519 3383
rect 107519 3349 107528 3383
rect 107476 3340 107528 3349
rect 109132 3340 109184 3392
rect 111064 3408 111116 3460
rect 117504 3476 117556 3528
rect 133052 3544 133104 3596
rect 134340 3612 134392 3664
rect 135260 3612 135312 3664
rect 188068 3612 188120 3664
rect 195152 3612 195204 3664
rect 145472 3544 145524 3596
rect 148140 3544 148192 3596
rect 158720 3544 158772 3596
rect 179420 3544 179472 3596
rect 180800 3544 180852 3596
rect 196164 3612 196216 3664
rect 210424 3680 210476 3732
rect 265992 3680 266044 3732
rect 270500 3680 270552 3732
rect 357440 3680 357492 3732
rect 372620 3680 372672 3732
rect 399300 3680 399352 3732
rect 301228 3612 301280 3664
rect 306564 3612 306616 3664
rect 395160 3612 395212 3664
rect 420920 3612 420972 3664
rect 444380 3612 444432 3664
rect 195336 3544 195388 3596
rect 296168 3544 296220 3596
rect 303988 3544 304040 3596
rect 392124 3544 392176 3596
rect 435364 3544 435416 3596
rect 480352 3544 480404 3596
rect 117596 3408 117648 3460
rect 122656 3408 122708 3460
rect 111892 3340 111944 3392
rect 114560 3383 114612 3392
rect 114560 3349 114569 3383
rect 114569 3349 114603 3383
rect 114603 3349 114612 3383
rect 114560 3340 114612 3349
rect 119344 3340 119396 3392
rect 121092 3383 121144 3392
rect 121092 3349 121101 3383
rect 121101 3349 121135 3383
rect 121135 3349 121144 3383
rect 121092 3340 121144 3349
rect 124220 3340 124272 3392
rect 125692 3340 125744 3392
rect 130476 3476 130528 3528
rect 132500 3476 132552 3528
rect 243728 3476 243780 3528
rect 273076 3476 273128 3528
rect 365812 3476 365864 3528
rect 395436 3476 395488 3528
rect 442080 3476 442132 3528
rect 128360 3340 128412 3392
rect 136088 3408 136140 3460
rect 220544 3408 220596 3460
rect 257620 3408 257672 3460
rect 363696 3408 363748 3460
rect 397368 3408 397420 3460
rect 443460 3408 443512 3460
rect 455972 3408 456024 3460
rect 482284 3408 482336 3460
rect 236000 3340 236052 3392
rect 296260 3340 296312 3392
rect 364708 3340 364760 3392
rect 67574 3238 67626 3290
rect 67638 3238 67690 3290
rect 67702 3238 67754 3290
rect 67766 3238 67818 3290
rect 67830 3238 67882 3290
rect 199502 3238 199554 3290
rect 199566 3238 199618 3290
rect 199630 3238 199682 3290
rect 199694 3238 199746 3290
rect 199758 3238 199810 3290
rect 331430 3238 331482 3290
rect 331494 3238 331546 3290
rect 331558 3238 331610 3290
rect 331622 3238 331674 3290
rect 331686 3238 331738 3290
rect 463358 3238 463410 3290
rect 463422 3238 463474 3290
rect 463486 3238 463538 3290
rect 463550 3238 463602 3290
rect 463614 3238 463666 3290
rect 61108 3136 61160 3188
rect 82820 3136 82872 3188
rect 94596 3136 94648 3188
rect 131764 3136 131816 3188
rect 132868 3136 132920 3188
rect 189172 3136 189224 3188
rect 194692 3136 194744 3188
rect 254216 3136 254268 3188
rect 351920 3136 351972 3188
rect 396264 3136 396316 3188
rect 485780 3136 485832 3188
rect 488540 3179 488592 3188
rect 488540 3145 488549 3179
rect 488549 3145 488583 3179
rect 488583 3145 488592 3179
rect 488540 3136 488592 3145
rect 491024 3179 491076 3188
rect 491024 3145 491033 3179
rect 491033 3145 491067 3179
rect 491067 3145 491076 3179
rect 491024 3136 491076 3145
rect 493600 3179 493652 3188
rect 493600 3145 493609 3179
rect 493609 3145 493643 3179
rect 493643 3145 493652 3179
rect 493600 3136 493652 3145
rect 496176 3179 496228 3188
rect 496176 3145 496185 3179
rect 496185 3145 496219 3179
rect 496219 3145 496228 3179
rect 496176 3136 496228 3145
rect 498752 3179 498804 3188
rect 498752 3145 498761 3179
rect 498761 3145 498795 3179
rect 498795 3145 498804 3179
rect 498752 3136 498804 3145
rect 501328 3179 501380 3188
rect 501328 3145 501337 3179
rect 501337 3145 501371 3179
rect 501371 3145 501380 3179
rect 501328 3136 501380 3145
rect 503904 3179 503956 3188
rect 503904 3145 503913 3179
rect 503913 3145 503947 3179
rect 503947 3145 503956 3179
rect 503904 3136 503956 3145
rect 506480 3179 506532 3188
rect 506480 3145 506489 3179
rect 506489 3145 506523 3179
rect 506523 3145 506532 3179
rect 506480 3136 506532 3145
rect 509056 3179 509108 3188
rect 509056 3145 509065 3179
rect 509065 3145 509099 3179
rect 509099 3145 509108 3179
rect 509056 3136 509108 3145
rect 511632 3179 511684 3188
rect 511632 3145 511641 3179
rect 511641 3145 511675 3179
rect 511675 3145 511684 3179
rect 511632 3136 511684 3145
rect 71228 3111 71280 3120
rect 71228 3077 71237 3111
rect 71237 3077 71271 3111
rect 71271 3077 71280 3111
rect 71228 3068 71280 3077
rect 74540 3068 74592 3120
rect 78496 3068 78548 3120
rect 78680 3068 78732 3120
rect 83648 3068 83700 3120
rect 86868 3068 86920 3120
rect 91560 3068 91612 3120
rect 96712 3068 96764 3120
rect 99104 3068 99156 3120
rect 99748 3068 99800 3120
rect 133604 3068 133656 3120
rect 27620 3000 27672 3052
rect 51540 2932 51592 2984
rect 85580 2932 85632 2984
rect 100852 3000 100904 3052
rect 107568 3000 107620 3052
rect 109684 3000 109736 3052
rect 116676 3000 116728 3052
rect 117596 3043 117648 3052
rect 117596 3009 117605 3043
rect 117605 3009 117639 3043
rect 117639 3009 117648 3043
rect 117596 3000 117648 3009
rect 128360 3000 128412 3052
rect 136088 3068 136140 3120
rect 181076 3068 181128 3120
rect 205456 3068 205508 3120
rect 210516 3068 210568 3120
rect 252652 3068 252704 3120
rect 134340 3000 134392 3052
rect 149152 3000 149204 3052
rect 184204 3000 184256 3052
rect 192852 3000 192904 3052
rect 195980 3000 196032 3052
rect 212540 3000 212592 3052
rect 101220 2932 101272 2984
rect 107476 2932 107528 2984
rect 137008 2932 137060 2984
rect 144000 2932 144052 2984
rect 249984 2932 250036 2984
rect 36820 2864 36872 2916
rect 40684 2864 40736 2916
rect 41328 2864 41380 2916
rect 45836 2864 45888 2916
rect 67916 2864 67968 2916
rect 71228 2864 71280 2916
rect 71780 2864 71832 2916
rect 76656 2864 76708 2916
rect 80060 2864 80112 2916
rect 86960 2864 87012 2916
rect 92020 2864 92072 2916
rect 130108 2864 130160 2916
rect 166908 2864 166960 2916
rect 195152 2864 195204 2916
rect 1308 2796 1360 2848
rect 3976 2839 4028 2848
rect 3976 2805 3985 2839
rect 3985 2805 4019 2839
rect 4019 2805 4028 2839
rect 3976 2796 4028 2805
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 8484 2796 8536 2848
rect 9128 2839 9180 2848
rect 9128 2805 9137 2839
rect 9137 2805 9171 2839
rect 9171 2805 9180 2839
rect 9128 2796 9180 2805
rect 14280 2839 14332 2848
rect 14280 2805 14289 2839
rect 14289 2805 14323 2839
rect 14323 2805 14332 2839
rect 14280 2796 14332 2805
rect 19248 2796 19300 2848
rect 23848 2796 23900 2848
rect 24584 2839 24636 2848
rect 24584 2805 24593 2839
rect 24593 2805 24627 2839
rect 24627 2805 24636 2839
rect 24584 2796 24636 2805
rect 28908 2796 28960 2848
rect 34888 2839 34940 2848
rect 34888 2805 34897 2839
rect 34897 2805 34931 2839
rect 34931 2805 34940 2839
rect 34888 2796 34940 2805
rect 37464 2839 37516 2848
rect 37464 2805 37473 2839
rect 37473 2805 37507 2839
rect 37507 2805 37516 2839
rect 37464 2796 37516 2805
rect 42800 2839 42852 2848
rect 42800 2805 42809 2839
rect 42809 2805 42843 2839
rect 42843 2805 42852 2839
rect 42800 2796 42852 2805
rect 50528 2839 50580 2848
rect 50528 2805 50537 2839
rect 50537 2805 50571 2839
rect 50571 2805 50580 2839
rect 50528 2796 50580 2805
rect 53104 2839 53156 2848
rect 53104 2805 53113 2839
rect 53113 2805 53147 2839
rect 53147 2805 53156 2839
rect 53104 2796 53156 2805
rect 53840 2796 53892 2848
rect 55128 2796 55180 2848
rect 58256 2839 58308 2848
rect 58256 2805 58265 2839
rect 58265 2805 58299 2839
rect 58299 2805 58308 2839
rect 58256 2796 58308 2805
rect 59360 2796 59412 2848
rect 60648 2796 60700 2848
rect 65248 2796 65300 2848
rect 68560 2839 68612 2848
rect 68560 2805 68569 2839
rect 68569 2805 68603 2839
rect 68603 2805 68612 2839
rect 68560 2796 68612 2805
rect 70400 2796 70452 2848
rect 71504 2796 71556 2848
rect 73160 2796 73212 2848
rect 81440 2839 81492 2848
rect 81440 2805 81449 2839
rect 81449 2805 81483 2839
rect 81483 2805 81492 2839
rect 81440 2796 81492 2805
rect 84016 2839 84068 2848
rect 84016 2805 84025 2839
rect 84025 2805 84059 2839
rect 84059 2805 84068 2839
rect 84016 2796 84068 2805
rect 89536 2796 89588 2848
rect 89720 2796 89772 2848
rect 92112 2796 92164 2848
rect 96620 2796 96672 2848
rect 99472 2839 99524 2848
rect 99472 2805 99481 2839
rect 99481 2805 99515 2839
rect 99515 2805 99524 2839
rect 99472 2796 99524 2805
rect 102140 2839 102192 2848
rect 102140 2805 102149 2839
rect 102149 2805 102183 2839
rect 102183 2805 102192 2839
rect 102140 2796 102192 2805
rect 104624 2839 104676 2848
rect 104624 2805 104633 2839
rect 104633 2805 104667 2839
rect 104667 2805 104676 2839
rect 104624 2796 104676 2805
rect 107384 2796 107436 2848
rect 111708 2796 111760 2848
rect 112352 2839 112404 2848
rect 112352 2805 112361 2839
rect 112361 2805 112395 2839
rect 112395 2805 112404 2839
rect 112352 2796 112404 2805
rect 112996 2796 113048 2848
rect 114652 2796 114704 2848
rect 115296 2796 115348 2848
rect 120080 2839 120132 2848
rect 120080 2805 120089 2839
rect 120089 2805 120123 2839
rect 120123 2805 120132 2839
rect 120080 2796 120132 2805
rect 121460 2796 121512 2848
rect 122656 2839 122708 2848
rect 122656 2805 122665 2839
rect 122665 2805 122699 2839
rect 122699 2805 122708 2839
rect 122656 2796 122708 2805
rect 128176 2796 128228 2848
rect 138020 2839 138072 2848
rect 138020 2805 138029 2839
rect 138029 2805 138063 2839
rect 138063 2805 138072 2839
rect 138020 2796 138072 2805
rect 143080 2839 143132 2848
rect 143080 2805 143089 2839
rect 143089 2805 143123 2839
rect 143123 2805 143132 2839
rect 143080 2796 143132 2805
rect 148232 2839 148284 2848
rect 148232 2805 148241 2839
rect 148241 2805 148275 2839
rect 148275 2805 148284 2839
rect 148232 2796 148284 2805
rect 153384 2839 153436 2848
rect 153384 2805 153393 2839
rect 153393 2805 153427 2839
rect 153427 2805 153436 2839
rect 153384 2796 153436 2805
rect 158536 2839 158588 2848
rect 158536 2805 158545 2839
rect 158545 2805 158579 2839
rect 158579 2805 158588 2839
rect 158536 2796 158588 2805
rect 163688 2839 163740 2848
rect 163688 2805 163697 2839
rect 163697 2805 163731 2839
rect 163731 2805 163740 2839
rect 163688 2796 163740 2805
rect 168380 2796 168432 2848
rect 173992 2839 174044 2848
rect 173992 2805 174001 2839
rect 174001 2805 174035 2839
rect 174035 2805 174044 2839
rect 173992 2796 174044 2805
rect 178040 2796 178092 2848
rect 179144 2839 179196 2848
rect 179144 2805 179153 2839
rect 179153 2805 179187 2839
rect 179187 2805 179196 2839
rect 179144 2796 179196 2805
rect 183560 2796 183612 2848
rect 189080 2796 189132 2848
rect 190460 2796 190512 2848
rect 202420 2864 202472 2916
rect 200028 2839 200080 2848
rect 200028 2805 200037 2839
rect 200037 2805 200071 2839
rect 200071 2805 200080 2839
rect 200028 2796 200080 2805
rect 205088 2839 205140 2848
rect 205088 2805 205097 2839
rect 205097 2805 205131 2839
rect 205131 2805 205140 2839
rect 205088 2796 205140 2805
rect 210240 2839 210292 2848
rect 210240 2805 210249 2839
rect 210249 2805 210283 2839
rect 210283 2805 210292 2839
rect 210240 2796 210292 2805
rect 215392 2839 215444 2848
rect 215392 2805 215401 2839
rect 215401 2805 215435 2839
rect 215435 2805 215444 2839
rect 215392 2796 215444 2805
rect 220544 2839 220596 2848
rect 220544 2805 220553 2839
rect 220553 2805 220587 2839
rect 220587 2805 220596 2839
rect 220544 2796 220596 2805
rect 226064 2796 226116 2848
rect 514208 2839 514260 2848
rect 514208 2805 514217 2839
rect 514217 2805 514251 2839
rect 514251 2805 514260 2839
rect 514208 2796 514260 2805
rect 66914 2694 66966 2746
rect 66978 2694 67030 2746
rect 67042 2694 67094 2746
rect 67106 2694 67158 2746
rect 67170 2694 67222 2746
rect 198842 2694 198894 2746
rect 198906 2694 198958 2746
rect 198970 2694 199022 2746
rect 199034 2694 199086 2746
rect 199098 2694 199150 2746
rect 330770 2694 330822 2746
rect 330834 2694 330886 2746
rect 330898 2694 330950 2746
rect 330962 2694 331014 2746
rect 331026 2694 331078 2746
rect 462698 2694 462750 2746
rect 462762 2694 462814 2746
rect 462826 2694 462878 2746
rect 462890 2694 462942 2746
rect 462954 2694 463006 2746
rect 5172 2635 5224 2644
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 59176 2592 59228 2644
rect 61108 2635 61160 2644
rect 61108 2601 61117 2635
rect 61117 2601 61151 2635
rect 61151 2601 61160 2635
rect 61108 2592 61160 2601
rect 68836 2635 68888 2644
rect 68836 2601 68845 2635
rect 68845 2601 68879 2635
rect 68879 2601 68888 2635
rect 68836 2592 68888 2601
rect 73988 2635 74040 2644
rect 73988 2601 73997 2635
rect 73997 2601 74031 2635
rect 74031 2601 74040 2635
rect 73988 2592 74040 2601
rect 76564 2635 76616 2644
rect 76564 2601 76573 2635
rect 76573 2601 76607 2635
rect 76607 2601 76616 2635
rect 76564 2592 76616 2601
rect 81716 2635 81768 2644
rect 81716 2601 81725 2635
rect 81725 2601 81759 2635
rect 81759 2601 81768 2635
rect 81716 2592 81768 2601
rect 87604 2635 87656 2644
rect 87604 2601 87613 2635
rect 87613 2601 87647 2635
rect 87647 2601 87656 2635
rect 87604 2592 87656 2601
rect 92388 2592 92440 2644
rect 97172 2635 97224 2644
rect 97172 2601 97181 2635
rect 97181 2601 97215 2635
rect 97215 2601 97224 2635
rect 97172 2592 97224 2601
rect 99104 2592 99156 2644
rect 103060 2635 103112 2644
rect 103060 2601 103069 2635
rect 103069 2601 103103 2635
rect 103103 2601 103112 2635
rect 103060 2592 103112 2601
rect 103428 2592 103480 2644
rect 107844 2592 107896 2644
rect 107936 2592 107988 2644
rect 109040 2592 109092 2644
rect 110052 2635 110104 2644
rect 110052 2601 110061 2635
rect 110061 2601 110095 2635
rect 110095 2601 110104 2635
rect 110052 2592 110104 2601
rect 110788 2635 110840 2644
rect 110788 2601 110797 2635
rect 110797 2601 110831 2635
rect 110831 2601 110840 2635
rect 110788 2592 110840 2601
rect 112628 2635 112680 2644
rect 112628 2601 112637 2635
rect 112637 2601 112671 2635
rect 112671 2601 112680 2635
rect 112628 2592 112680 2601
rect 12900 2567 12952 2576
rect 12900 2533 12909 2567
rect 12909 2533 12943 2567
rect 12943 2533 12952 2567
rect 12900 2524 12952 2533
rect 18052 2567 18104 2576
rect 18052 2533 18061 2567
rect 18061 2533 18095 2567
rect 18095 2533 18104 2567
rect 18052 2524 18104 2533
rect 42892 2524 42944 2576
rect 5172 2388 5224 2440
rect 6736 2388 6788 2440
rect 12900 2388 12952 2440
rect 18052 2388 18104 2440
rect 848 2320 900 2372
rect 6000 2320 6052 2372
rect 6552 2320 6604 2372
rect 10784 2320 10836 2372
rect 15936 2320 15988 2372
rect 23204 2363 23256 2372
rect 23204 2329 23213 2363
rect 23213 2329 23247 2363
rect 23247 2329 23256 2363
rect 23204 2320 23256 2329
rect 28356 2363 28408 2372
rect 28356 2329 28365 2363
rect 28365 2329 28399 2363
rect 28399 2329 28408 2363
rect 28356 2320 28408 2329
rect 4160 2252 4212 2304
rect 7012 2295 7064 2304
rect 7012 2261 7021 2295
rect 7021 2261 7055 2295
rect 7055 2261 7064 2295
rect 7012 2252 7064 2261
rect 9588 2252 9640 2304
rect 14740 2295 14792 2304
rect 14740 2261 14749 2295
rect 14749 2261 14783 2295
rect 14783 2261 14792 2295
rect 14740 2252 14792 2261
rect 17316 2295 17368 2304
rect 17316 2261 17325 2295
rect 17325 2261 17359 2295
rect 17359 2261 17368 2295
rect 17316 2252 17368 2261
rect 20720 2252 20772 2304
rect 23940 2295 23992 2304
rect 23940 2261 23949 2295
rect 23949 2261 23983 2295
rect 23983 2261 23992 2295
rect 23940 2252 23992 2261
rect 25044 2295 25096 2304
rect 25044 2261 25053 2295
rect 25053 2261 25087 2295
rect 25087 2261 25096 2295
rect 25044 2252 25096 2261
rect 27620 2295 27672 2304
rect 27620 2261 27629 2295
rect 27629 2261 27663 2295
rect 27663 2261 27672 2295
rect 27620 2252 27672 2261
rect 28264 2252 28316 2304
rect 33508 2499 33560 2508
rect 33508 2465 33517 2499
rect 33517 2465 33551 2499
rect 33551 2465 33560 2499
rect 33508 2456 33560 2465
rect 41236 2499 41288 2508
rect 40408 2388 40460 2440
rect 41236 2465 41245 2499
rect 41245 2465 41279 2499
rect 41279 2465 41288 2499
rect 41236 2456 41288 2465
rect 103980 2456 104032 2508
rect 42800 2388 42852 2440
rect 34888 2320 34940 2372
rect 37464 2320 37516 2372
rect 30196 2295 30248 2304
rect 30196 2261 30205 2295
rect 30205 2261 30239 2295
rect 30239 2261 30248 2295
rect 30196 2252 30248 2261
rect 32772 2295 32824 2304
rect 32772 2261 32781 2295
rect 32781 2261 32815 2295
rect 32815 2261 32824 2295
rect 32772 2252 32824 2261
rect 35348 2295 35400 2304
rect 35348 2261 35357 2295
rect 35357 2261 35391 2295
rect 35391 2261 35400 2295
rect 35348 2252 35400 2261
rect 37924 2295 37976 2304
rect 37924 2261 37933 2295
rect 37933 2261 37967 2295
rect 37967 2261 37976 2295
rect 37924 2252 37976 2261
rect 38660 2252 38712 2304
rect 44088 2252 44140 2304
rect 48964 2431 49016 2440
rect 48964 2397 48973 2431
rect 48973 2397 49007 2431
rect 49007 2397 49016 2431
rect 48964 2388 49016 2397
rect 50528 2388 50580 2440
rect 53104 2388 53156 2440
rect 53564 2431 53616 2440
rect 53564 2397 53573 2431
rect 53573 2397 53607 2431
rect 53607 2397 53616 2431
rect 53564 2388 53616 2397
rect 56600 2431 56652 2440
rect 56600 2397 56609 2431
rect 56609 2397 56643 2431
rect 56643 2397 56652 2431
rect 56600 2388 56652 2397
rect 57980 2388 58032 2440
rect 58256 2388 58308 2440
rect 52644 2320 52696 2372
rect 46020 2252 46072 2304
rect 50804 2295 50856 2304
rect 50804 2261 50813 2295
rect 50813 2261 50847 2295
rect 50847 2261 50856 2295
rect 50804 2252 50856 2261
rect 53380 2295 53432 2304
rect 53380 2261 53389 2295
rect 53389 2261 53423 2295
rect 53423 2261 53432 2295
rect 53380 2252 53432 2261
rect 57888 2320 57940 2372
rect 65248 2388 65300 2440
rect 68560 2388 68612 2440
rect 73160 2388 73212 2440
rect 75552 2388 75604 2440
rect 79232 2388 79284 2440
rect 87604 2388 87656 2440
rect 94136 2388 94188 2440
rect 95332 2431 95384 2440
rect 95332 2397 95341 2431
rect 95341 2397 95375 2431
rect 95375 2397 95384 2431
rect 95332 2388 95384 2397
rect 99196 2388 99248 2440
rect 81440 2320 81492 2372
rect 84108 2320 84160 2372
rect 86776 2320 86828 2372
rect 89536 2363 89588 2372
rect 89536 2329 89545 2363
rect 89545 2329 89579 2363
rect 89579 2329 89588 2363
rect 89536 2320 89588 2329
rect 58532 2295 58584 2304
rect 58532 2261 58541 2295
rect 58541 2261 58575 2295
rect 58575 2261 58584 2295
rect 58532 2252 58584 2261
rect 63684 2295 63736 2304
rect 63684 2261 63693 2295
rect 63693 2261 63727 2295
rect 63727 2261 63736 2295
rect 63684 2252 63736 2261
rect 64420 2295 64472 2304
rect 64420 2261 64429 2295
rect 64429 2261 64463 2295
rect 64463 2261 64472 2295
rect 64420 2252 64472 2261
rect 66260 2295 66312 2304
rect 66260 2261 66269 2295
rect 66269 2261 66303 2295
rect 66303 2261 66312 2295
rect 66260 2252 66312 2261
rect 71412 2295 71464 2304
rect 71412 2261 71421 2295
rect 71421 2261 71455 2295
rect 71455 2261 71464 2295
rect 71412 2252 71464 2261
rect 72148 2295 72200 2304
rect 72148 2261 72157 2295
rect 72157 2261 72191 2295
rect 72191 2261 72200 2295
rect 72148 2252 72200 2261
rect 75460 2295 75512 2304
rect 75460 2261 75469 2295
rect 75469 2261 75503 2295
rect 75503 2261 75512 2295
rect 75460 2252 75512 2261
rect 77300 2252 77352 2304
rect 79876 2295 79928 2304
rect 79876 2261 79885 2295
rect 79885 2261 79919 2295
rect 79919 2261 79928 2295
rect 79876 2252 79928 2261
rect 84292 2295 84344 2304
rect 84292 2261 84301 2295
rect 84301 2261 84335 2295
rect 84335 2261 84344 2295
rect 84292 2252 84344 2261
rect 84476 2252 84528 2304
rect 86960 2252 87012 2304
rect 91284 2252 91336 2304
rect 92296 2252 92348 2304
rect 96620 2320 96672 2372
rect 99472 2320 99524 2372
rect 103060 2388 103112 2440
rect 104164 2524 104216 2576
rect 107384 2567 107436 2576
rect 107384 2533 107393 2567
rect 107393 2533 107427 2567
rect 107427 2533 107436 2567
rect 107384 2524 107436 2533
rect 111708 2524 111760 2576
rect 126888 2592 126940 2644
rect 141148 2592 141200 2644
rect 187332 2592 187384 2644
rect 187424 2592 187476 2644
rect 193220 2635 193272 2644
rect 193220 2601 193229 2635
rect 193229 2601 193263 2635
rect 193263 2601 193272 2635
rect 193220 2592 193272 2601
rect 194508 2592 194560 2644
rect 205364 2635 205416 2644
rect 205364 2601 205373 2635
rect 205373 2601 205407 2635
rect 205407 2601 205416 2635
rect 205364 2592 205416 2601
rect 208584 2635 208636 2644
rect 208584 2601 208593 2635
rect 208593 2601 208627 2635
rect 208627 2601 208636 2635
rect 208584 2592 208636 2601
rect 210516 2635 210568 2644
rect 210516 2601 210525 2635
rect 210525 2601 210559 2635
rect 210559 2601 210568 2635
rect 210516 2592 210568 2601
rect 224132 2635 224184 2644
rect 224132 2601 224141 2635
rect 224141 2601 224175 2635
rect 224175 2601 224184 2635
rect 224132 2592 224184 2601
rect 229192 2635 229244 2644
rect 229192 2601 229201 2635
rect 229201 2601 229235 2635
rect 229235 2601 229244 2635
rect 229192 2592 229244 2601
rect 231860 2635 231912 2644
rect 231860 2601 231869 2635
rect 231869 2601 231903 2635
rect 231903 2601 231912 2635
rect 231860 2592 231912 2601
rect 232872 2592 232924 2644
rect 234436 2635 234488 2644
rect 234436 2601 234445 2635
rect 234445 2601 234479 2635
rect 234479 2601 234488 2635
rect 234436 2592 234488 2601
rect 237012 2635 237064 2644
rect 237012 2601 237021 2635
rect 237021 2601 237055 2635
rect 237055 2601 237064 2635
rect 237012 2592 237064 2601
rect 242164 2635 242216 2644
rect 242164 2601 242173 2635
rect 242173 2601 242207 2635
rect 242207 2601 242216 2635
rect 242164 2592 242216 2601
rect 244832 2592 244884 2644
rect 247224 2635 247276 2644
rect 247224 2601 247233 2635
rect 247233 2601 247267 2635
rect 247267 2601 247276 2635
rect 247224 2592 247276 2601
rect 249892 2635 249944 2644
rect 249892 2601 249901 2635
rect 249901 2601 249935 2635
rect 249935 2601 249944 2635
rect 249892 2592 249944 2601
rect 257620 2635 257672 2644
rect 257620 2601 257629 2635
rect 257629 2601 257663 2635
rect 257663 2601 257672 2635
rect 257620 2592 257672 2601
rect 260196 2635 260248 2644
rect 260196 2601 260205 2635
rect 260205 2601 260239 2635
rect 260239 2601 260248 2635
rect 260196 2592 260248 2601
rect 265348 2635 265400 2644
rect 265348 2601 265357 2635
rect 265357 2601 265391 2635
rect 265391 2601 265400 2635
rect 265348 2592 265400 2601
rect 270500 2635 270552 2644
rect 270500 2601 270509 2635
rect 270509 2601 270543 2635
rect 270543 2601 270552 2635
rect 270500 2592 270552 2601
rect 273076 2635 273128 2644
rect 273076 2601 273085 2635
rect 273085 2601 273119 2635
rect 273119 2601 273128 2635
rect 273076 2592 273128 2601
rect 275652 2635 275704 2644
rect 275652 2601 275661 2635
rect 275661 2601 275695 2635
rect 275695 2601 275704 2635
rect 275652 2592 275704 2601
rect 280804 2635 280856 2644
rect 280804 2601 280813 2635
rect 280813 2601 280847 2635
rect 280847 2601 280856 2635
rect 280804 2592 280856 2601
rect 283380 2635 283432 2644
rect 283380 2601 283389 2635
rect 283389 2601 283423 2635
rect 283423 2601 283432 2635
rect 283380 2592 283432 2601
rect 285956 2635 286008 2644
rect 285956 2601 285965 2635
rect 285965 2601 285999 2635
rect 285999 2601 286008 2635
rect 285956 2592 286008 2601
rect 288532 2635 288584 2644
rect 288532 2601 288541 2635
rect 288541 2601 288575 2635
rect 288575 2601 288584 2635
rect 288532 2592 288584 2601
rect 291108 2635 291160 2644
rect 291108 2601 291117 2635
rect 291117 2601 291151 2635
rect 291151 2601 291160 2635
rect 291108 2592 291160 2601
rect 293684 2635 293736 2644
rect 293684 2601 293693 2635
rect 293693 2601 293727 2635
rect 293727 2601 293736 2635
rect 293684 2592 293736 2601
rect 296260 2635 296312 2644
rect 296260 2601 296269 2635
rect 296269 2601 296303 2635
rect 296303 2601 296312 2635
rect 296260 2592 296312 2601
rect 298836 2635 298888 2644
rect 298836 2601 298845 2635
rect 298845 2601 298879 2635
rect 298879 2601 298888 2635
rect 298836 2592 298888 2601
rect 301412 2635 301464 2644
rect 301412 2601 301421 2635
rect 301421 2601 301455 2635
rect 301455 2601 301464 2635
rect 301412 2592 301464 2601
rect 107660 2456 107712 2508
rect 107844 2456 107896 2508
rect 110052 2456 110104 2508
rect 110328 2456 110380 2508
rect 109776 2388 109828 2440
rect 110788 2388 110840 2440
rect 172520 2524 172572 2576
rect 172612 2524 172664 2576
rect 176752 2524 176804 2576
rect 177212 2524 177264 2576
rect 180800 2524 180852 2576
rect 182916 2567 182968 2576
rect 182916 2533 182925 2567
rect 182925 2533 182959 2567
rect 182959 2533 182968 2567
rect 182916 2524 182968 2533
rect 260840 2524 260892 2576
rect 282460 2524 282512 2576
rect 291200 2524 291252 2576
rect 126428 2456 126480 2508
rect 130476 2456 130528 2508
rect 119436 2388 119488 2440
rect 104624 2320 104676 2372
rect 99748 2295 99800 2304
rect 99748 2261 99757 2295
rect 99757 2261 99791 2295
rect 99791 2261 99800 2295
rect 99748 2252 99800 2261
rect 104900 2295 104952 2304
rect 104900 2261 104909 2295
rect 104909 2261 104943 2295
rect 104943 2261 104952 2295
rect 104900 2252 104952 2261
rect 106372 2295 106424 2304
rect 106372 2261 106381 2295
rect 106381 2261 106415 2295
rect 106415 2261 106424 2295
rect 112352 2320 112404 2372
rect 115296 2363 115348 2372
rect 115296 2329 115305 2363
rect 115305 2329 115339 2363
rect 115339 2329 115348 2363
rect 115296 2320 115348 2329
rect 120080 2320 120132 2372
rect 128268 2388 128320 2440
rect 130660 2431 130712 2440
rect 130660 2397 130669 2431
rect 130669 2397 130703 2431
rect 130703 2397 130712 2431
rect 130660 2388 130712 2397
rect 127072 2320 127124 2372
rect 128176 2363 128228 2372
rect 128176 2329 128185 2363
rect 128185 2329 128219 2363
rect 128219 2329 128228 2363
rect 128176 2320 128228 2329
rect 128360 2320 128412 2372
rect 106372 2252 106424 2261
rect 107752 2252 107804 2304
rect 109224 2252 109276 2304
rect 115204 2295 115256 2304
rect 115204 2261 115213 2295
rect 115213 2261 115247 2295
rect 115247 2261 115256 2295
rect 115204 2252 115256 2261
rect 120356 2295 120408 2304
rect 120356 2261 120365 2295
rect 120365 2261 120399 2295
rect 120399 2261 120408 2295
rect 120356 2252 120408 2261
rect 122932 2295 122984 2304
rect 122932 2261 122941 2295
rect 122941 2261 122975 2295
rect 122975 2261 122984 2295
rect 122932 2252 122984 2261
rect 125508 2295 125560 2304
rect 125508 2261 125517 2295
rect 125517 2261 125551 2295
rect 125551 2261 125560 2295
rect 125508 2252 125560 2261
rect 126244 2295 126296 2304
rect 126244 2261 126253 2295
rect 126253 2261 126287 2295
rect 126287 2261 126296 2295
rect 126244 2252 126296 2261
rect 128084 2295 128136 2304
rect 128084 2261 128093 2295
rect 128093 2261 128127 2295
rect 128127 2261 128136 2295
rect 128084 2252 128136 2261
rect 130844 2295 130896 2304
rect 130844 2261 130853 2295
rect 130853 2261 130887 2295
rect 130887 2261 130896 2295
rect 130844 2252 130896 2261
rect 150808 2456 150860 2508
rect 253940 2456 253992 2508
rect 263416 2456 263468 2508
rect 133972 2295 134024 2304
rect 133972 2261 133981 2295
rect 133981 2261 134015 2295
rect 134015 2261 134024 2295
rect 133972 2252 134024 2261
rect 138112 2388 138164 2440
rect 141148 2431 141200 2440
rect 141148 2397 141157 2431
rect 141157 2397 141191 2431
rect 141191 2397 141200 2431
rect 141148 2388 141200 2397
rect 143080 2388 143132 2440
rect 136456 2252 136508 2304
rect 143448 2363 143500 2372
rect 143448 2329 143457 2363
rect 143457 2329 143491 2363
rect 143491 2329 143500 2363
rect 143448 2320 143500 2329
rect 148232 2388 148284 2440
rect 146852 2363 146904 2372
rect 144920 2252 144972 2304
rect 146852 2329 146861 2363
rect 146861 2329 146895 2363
rect 146895 2329 146904 2363
rect 146852 2320 146904 2329
rect 148600 2363 148652 2372
rect 148600 2329 148609 2363
rect 148609 2329 148643 2363
rect 148643 2329 148652 2363
rect 148600 2320 148652 2329
rect 153384 2388 153436 2440
rect 158904 2431 158956 2440
rect 158904 2397 158913 2431
rect 158913 2397 158947 2431
rect 158947 2397 158956 2431
rect 158904 2388 158956 2397
rect 158536 2320 158588 2372
rect 161940 2388 161992 2440
rect 163688 2320 163740 2372
rect 146668 2252 146720 2304
rect 151268 2295 151320 2304
rect 151268 2261 151277 2295
rect 151277 2261 151311 2295
rect 151311 2261 151320 2295
rect 151268 2252 151320 2261
rect 152004 2295 152056 2304
rect 152004 2261 152013 2295
rect 152013 2261 152047 2295
rect 152047 2261 152056 2295
rect 152004 2252 152056 2261
rect 156420 2295 156472 2304
rect 156420 2261 156429 2295
rect 156429 2261 156463 2295
rect 156463 2261 156472 2295
rect 156420 2252 156472 2261
rect 157156 2295 157208 2304
rect 157156 2261 157165 2295
rect 157165 2261 157199 2295
rect 157199 2261 157208 2295
rect 157156 2252 157208 2261
rect 161572 2295 161624 2304
rect 161572 2261 161581 2295
rect 161581 2261 161615 2295
rect 161615 2261 161624 2295
rect 161572 2252 161624 2261
rect 162308 2295 162360 2304
rect 162308 2261 162317 2295
rect 162317 2261 162351 2295
rect 162351 2261 162360 2295
rect 162308 2252 162360 2261
rect 164148 2295 164200 2304
rect 164148 2261 164157 2295
rect 164157 2261 164191 2295
rect 164191 2261 164200 2295
rect 164148 2252 164200 2261
rect 168380 2320 168432 2372
rect 177212 2431 177264 2440
rect 177212 2397 177221 2431
rect 177221 2397 177255 2431
rect 177255 2397 177264 2431
rect 177212 2388 177264 2397
rect 179144 2388 179196 2440
rect 182916 2388 182968 2440
rect 184296 2388 184348 2440
rect 187424 2388 187476 2440
rect 188068 2431 188120 2440
rect 188068 2397 188077 2431
rect 188077 2397 188111 2431
rect 188111 2397 188120 2431
rect 188068 2388 188120 2397
rect 173992 2320 174044 2372
rect 175004 2320 175056 2372
rect 183560 2320 183612 2372
rect 185492 2320 185544 2372
rect 186780 2320 186832 2372
rect 186872 2320 186924 2372
rect 191748 2388 191800 2440
rect 193220 2388 193272 2440
rect 195152 2431 195204 2440
rect 195152 2397 195161 2431
rect 195161 2397 195195 2431
rect 195195 2397 195204 2431
rect 195152 2388 195204 2397
rect 197820 2431 197872 2440
rect 197820 2397 197829 2431
rect 197829 2397 197863 2431
rect 197863 2397 197872 2431
rect 197820 2388 197872 2397
rect 200028 2388 200080 2440
rect 203064 2388 203116 2440
rect 205088 2388 205140 2440
rect 208584 2388 208636 2440
rect 210240 2388 210292 2440
rect 213276 2431 213328 2440
rect 213276 2397 213285 2431
rect 213285 2397 213319 2431
rect 213319 2397 213328 2431
rect 213276 2388 213328 2397
rect 215392 2388 215444 2440
rect 218428 2431 218480 2440
rect 218428 2397 218437 2431
rect 218437 2397 218471 2431
rect 218471 2397 218480 2431
rect 218428 2388 218480 2397
rect 220544 2388 220596 2440
rect 224132 2388 224184 2440
rect 229192 2388 229244 2440
rect 231860 2388 231912 2440
rect 234436 2388 234488 2440
rect 237012 2388 237064 2440
rect 239036 2431 239088 2440
rect 239036 2397 239045 2431
rect 239045 2397 239079 2431
rect 239079 2397 239088 2431
rect 239036 2388 239088 2397
rect 242164 2388 242216 2440
rect 244832 2388 244884 2440
rect 247224 2388 247276 2440
rect 249892 2388 249944 2440
rect 251916 2431 251968 2440
rect 251916 2397 251925 2431
rect 251925 2397 251959 2431
rect 251959 2397 251968 2431
rect 251916 2388 251968 2397
rect 189080 2320 189132 2372
rect 167460 2295 167512 2304
rect 167460 2261 167469 2295
rect 167469 2261 167503 2295
rect 167503 2261 167512 2295
rect 167460 2252 167512 2261
rect 169300 2295 169352 2304
rect 169300 2261 169309 2295
rect 169309 2261 169343 2295
rect 169343 2261 169352 2295
rect 169300 2252 169352 2261
rect 171140 2252 171192 2304
rect 172612 2295 172664 2304
rect 172612 2261 172621 2295
rect 172621 2261 172655 2295
rect 172655 2261 172664 2295
rect 172612 2252 172664 2261
rect 174452 2295 174504 2304
rect 174452 2261 174461 2295
rect 174461 2261 174495 2295
rect 174495 2261 174504 2295
rect 174452 2252 174504 2261
rect 174636 2252 174688 2304
rect 179604 2295 179656 2304
rect 179604 2261 179613 2295
rect 179613 2261 179647 2295
rect 179647 2261 179656 2295
rect 179604 2252 179656 2261
rect 182180 2295 182232 2304
rect 182180 2261 182189 2295
rect 182189 2261 182223 2295
rect 182223 2261 182232 2295
rect 182180 2252 182232 2261
rect 183652 2252 183704 2304
rect 195336 2320 195388 2372
rect 195060 2295 195112 2304
rect 195060 2261 195069 2295
rect 195069 2261 195103 2295
rect 195103 2261 195112 2295
rect 195060 2252 195112 2261
rect 195152 2252 195204 2304
rect 226064 2363 226116 2372
rect 226064 2329 226073 2363
rect 226073 2329 226107 2363
rect 226107 2329 226116 2363
rect 226064 2320 226116 2329
rect 233240 2320 233292 2372
rect 195980 2252 196032 2304
rect 200212 2295 200264 2304
rect 200212 2261 200221 2295
rect 200221 2261 200255 2295
rect 200255 2261 200264 2295
rect 200212 2252 200264 2261
rect 202788 2295 202840 2304
rect 202788 2261 202797 2295
rect 202797 2261 202831 2295
rect 202831 2261 202840 2295
rect 202788 2252 202840 2261
rect 207940 2295 207992 2304
rect 207940 2261 207949 2295
rect 207949 2261 207983 2295
rect 207983 2261 207992 2295
rect 207940 2252 207992 2261
rect 213092 2295 213144 2304
rect 213092 2261 213101 2295
rect 213101 2261 213135 2295
rect 213135 2261 213144 2295
rect 213092 2252 213144 2261
rect 215668 2295 215720 2304
rect 215668 2261 215677 2295
rect 215677 2261 215711 2295
rect 215711 2261 215720 2295
rect 215668 2252 215720 2261
rect 218244 2295 218296 2304
rect 218244 2261 218253 2295
rect 218253 2261 218287 2295
rect 218287 2261 218296 2295
rect 218244 2252 218296 2261
rect 220820 2295 220872 2304
rect 220820 2261 220829 2295
rect 220829 2261 220863 2295
rect 220863 2261 220872 2295
rect 220820 2252 220872 2261
rect 223396 2295 223448 2304
rect 223396 2261 223405 2295
rect 223405 2261 223439 2295
rect 223439 2261 223448 2295
rect 223396 2252 223448 2261
rect 225972 2295 226024 2304
rect 225972 2261 225981 2295
rect 225981 2261 226015 2295
rect 226015 2261 226024 2295
rect 225972 2252 226024 2261
rect 228548 2295 228600 2304
rect 228548 2261 228557 2295
rect 228557 2261 228591 2295
rect 228591 2261 228600 2295
rect 228548 2252 228600 2261
rect 229100 2252 229152 2304
rect 233700 2295 233752 2304
rect 233700 2261 233709 2295
rect 233709 2261 233743 2295
rect 233743 2261 233752 2295
rect 233700 2252 233752 2261
rect 236276 2295 236328 2304
rect 236276 2261 236285 2295
rect 236285 2261 236319 2295
rect 236319 2261 236328 2295
rect 236276 2252 236328 2261
rect 243912 2320 243964 2372
rect 241428 2295 241480 2304
rect 241428 2261 241437 2295
rect 241437 2261 241471 2295
rect 241471 2261 241480 2295
rect 241428 2252 241480 2261
rect 242900 2252 242952 2304
rect 244096 2252 244148 2304
rect 247040 2252 247092 2304
rect 257620 2388 257672 2440
rect 260196 2388 260248 2440
rect 262220 2431 262272 2440
rect 262220 2397 262229 2431
rect 262229 2397 262263 2431
rect 262263 2397 262272 2431
rect 262220 2388 262272 2397
rect 265348 2388 265400 2440
rect 291752 2456 291804 2508
rect 298192 2456 298244 2508
rect 303988 2635 304040 2644
rect 303988 2601 303997 2635
rect 303997 2601 304031 2635
rect 304031 2601 304040 2635
rect 303988 2592 304040 2601
rect 306564 2635 306616 2644
rect 306564 2601 306573 2635
rect 306573 2601 306607 2635
rect 306607 2601 306616 2635
rect 306564 2592 306616 2601
rect 309140 2635 309192 2644
rect 309140 2601 309149 2635
rect 309149 2601 309183 2635
rect 309183 2601 309192 2635
rect 309140 2592 309192 2601
rect 303528 2524 303580 2576
rect 306380 2456 306432 2508
rect 319260 2592 319312 2644
rect 322020 2635 322072 2644
rect 322020 2601 322029 2635
rect 322029 2601 322063 2635
rect 322063 2601 322072 2635
rect 322020 2592 322072 2601
rect 270500 2388 270552 2440
rect 273076 2388 273128 2440
rect 275652 2388 275704 2440
rect 253848 2252 253900 2304
rect 255044 2295 255096 2304
rect 255044 2261 255053 2295
rect 255053 2261 255087 2295
rect 255087 2261 255096 2295
rect 255044 2252 255096 2261
rect 255412 2252 255464 2304
rect 258080 2252 258132 2304
rect 260840 2252 260892 2304
rect 263600 2252 263652 2304
rect 267188 2295 267240 2304
rect 267188 2261 267197 2295
rect 267197 2261 267231 2295
rect 267231 2261 267240 2295
rect 267188 2252 267240 2261
rect 267924 2295 267976 2304
rect 267924 2261 267933 2295
rect 267933 2261 267967 2295
rect 267967 2261 267976 2295
rect 267924 2252 267976 2261
rect 268016 2252 268068 2304
rect 269856 2252 269908 2304
rect 280804 2388 280856 2440
rect 283380 2388 283432 2440
rect 285956 2388 286008 2440
rect 288532 2388 288584 2440
rect 291108 2388 291160 2440
rect 293684 2388 293736 2440
rect 296260 2388 296312 2440
rect 298836 2388 298888 2440
rect 301412 2388 301464 2440
rect 303988 2388 304040 2440
rect 306564 2388 306616 2440
rect 309140 2388 309192 2440
rect 314292 2388 314344 2440
rect 302700 2320 302752 2372
rect 276020 2252 276072 2304
rect 278228 2295 278280 2304
rect 278228 2261 278237 2295
rect 278237 2261 278271 2295
rect 278271 2261 278280 2295
rect 278228 2252 278280 2261
rect 278780 2252 278832 2304
rect 282644 2295 282696 2304
rect 282644 2261 282653 2295
rect 282653 2261 282687 2295
rect 282687 2261 282696 2295
rect 282644 2252 282696 2261
rect 282736 2252 282788 2304
rect 285680 2252 285732 2304
rect 289912 2252 289964 2304
rect 295248 2252 295300 2304
rect 300860 2252 300912 2304
rect 309232 2320 309284 2372
rect 319444 2388 319496 2440
rect 322020 2388 322072 2440
rect 314292 2295 314344 2304
rect 314292 2261 314301 2295
rect 314301 2261 314335 2295
rect 314335 2261 314344 2295
rect 314292 2252 314344 2261
rect 316684 2320 316736 2372
rect 318708 2295 318760 2304
rect 318708 2261 318717 2295
rect 318717 2261 318751 2295
rect 318751 2261 318760 2295
rect 318708 2252 318760 2261
rect 319444 2295 319496 2304
rect 319444 2261 319453 2295
rect 319453 2261 319487 2295
rect 319487 2261 319496 2295
rect 319444 2252 319496 2261
rect 321284 2295 321336 2304
rect 321284 2261 321293 2295
rect 321293 2261 321327 2295
rect 321327 2261 321336 2295
rect 321284 2252 321336 2261
rect 334900 2567 334952 2576
rect 334900 2533 334909 2567
rect 334909 2533 334943 2567
rect 334943 2533 334952 2567
rect 334900 2524 334952 2533
rect 329748 2388 329800 2440
rect 332324 2388 332376 2440
rect 337476 2388 337528 2440
rect 340052 2388 340104 2440
rect 342628 2388 342680 2440
rect 345204 2388 345256 2440
rect 349068 2524 349120 2576
rect 355416 2524 355468 2576
rect 355508 2567 355560 2576
rect 355508 2533 355517 2567
rect 355517 2533 355551 2567
rect 355551 2533 355560 2567
rect 355508 2524 355560 2533
rect 351920 2456 351972 2508
rect 352932 2499 352984 2508
rect 352932 2465 352941 2499
rect 352941 2465 352975 2499
rect 352975 2465 352984 2499
rect 352932 2456 352984 2465
rect 360660 2635 360712 2644
rect 360660 2601 360669 2635
rect 360669 2601 360703 2635
rect 360703 2601 360712 2635
rect 360660 2592 360712 2601
rect 365076 2635 365128 2644
rect 365076 2601 365085 2635
rect 365085 2601 365119 2635
rect 365119 2601 365128 2635
rect 365076 2592 365128 2601
rect 365260 2592 365312 2644
rect 369860 2592 369912 2644
rect 373540 2592 373592 2644
rect 376116 2635 376168 2644
rect 376116 2601 376125 2635
rect 376125 2601 376159 2635
rect 376159 2601 376168 2635
rect 376116 2592 376168 2601
rect 378048 2592 378100 2644
rect 378140 2592 378192 2644
rect 383200 2592 383252 2644
rect 383292 2592 383344 2644
rect 383844 2592 383896 2644
rect 390652 2592 390704 2644
rect 394056 2592 394108 2644
rect 398748 2592 398800 2644
rect 408500 2592 408552 2644
rect 373448 2524 373500 2576
rect 380900 2524 380952 2576
rect 381084 2524 381136 2576
rect 385040 2524 385092 2576
rect 391940 2524 391992 2576
rect 392032 2524 392084 2576
rect 393320 2524 393372 2576
rect 395252 2524 395304 2576
rect 397644 2524 397696 2576
rect 400220 2524 400272 2576
rect 404360 2567 404412 2576
rect 404360 2533 404369 2567
rect 404369 2533 404403 2567
rect 404403 2533 404412 2567
rect 404360 2524 404412 2533
rect 369952 2456 370004 2508
rect 350356 2363 350408 2372
rect 350356 2329 350365 2363
rect 350365 2329 350399 2363
rect 350399 2329 350408 2363
rect 350356 2320 350408 2329
rect 324596 2295 324648 2304
rect 324596 2261 324605 2295
rect 324605 2261 324639 2295
rect 324639 2261 324648 2295
rect 324596 2252 324648 2261
rect 326436 2295 326488 2304
rect 326436 2261 326445 2295
rect 326445 2261 326479 2295
rect 326479 2261 326488 2295
rect 326436 2252 326488 2261
rect 329012 2295 329064 2304
rect 329012 2261 329021 2295
rect 329021 2261 329055 2295
rect 329055 2261 329064 2295
rect 329012 2252 329064 2261
rect 329748 2295 329800 2304
rect 329748 2261 329757 2295
rect 329757 2261 329791 2295
rect 329791 2261 329800 2295
rect 329748 2252 329800 2261
rect 331220 2252 331272 2304
rect 332324 2295 332376 2304
rect 332324 2261 332333 2295
rect 332333 2261 332367 2295
rect 332367 2261 332376 2295
rect 332324 2252 332376 2261
rect 334164 2295 334216 2304
rect 334164 2261 334173 2295
rect 334173 2261 334207 2295
rect 334207 2261 334216 2295
rect 334164 2252 334216 2261
rect 336740 2295 336792 2304
rect 336740 2261 336749 2295
rect 336749 2261 336783 2295
rect 336783 2261 336792 2295
rect 336740 2252 336792 2261
rect 337476 2295 337528 2304
rect 337476 2261 337485 2295
rect 337485 2261 337519 2295
rect 337519 2261 337528 2295
rect 337476 2252 337528 2261
rect 339316 2295 339368 2304
rect 339316 2261 339325 2295
rect 339325 2261 339359 2295
rect 339359 2261 339368 2295
rect 339316 2252 339368 2261
rect 340052 2295 340104 2304
rect 340052 2261 340061 2295
rect 340061 2261 340095 2295
rect 340095 2261 340104 2295
rect 340052 2252 340104 2261
rect 341892 2295 341944 2304
rect 341892 2261 341901 2295
rect 341901 2261 341935 2295
rect 341935 2261 341944 2295
rect 341892 2252 341944 2261
rect 342628 2295 342680 2304
rect 342628 2261 342637 2295
rect 342637 2261 342671 2295
rect 342671 2261 342680 2295
rect 342628 2252 342680 2261
rect 344468 2295 344520 2304
rect 344468 2261 344477 2295
rect 344477 2261 344511 2295
rect 344511 2261 344520 2295
rect 344468 2252 344520 2261
rect 345204 2295 345256 2304
rect 345204 2261 345213 2295
rect 345213 2261 345247 2295
rect 345247 2261 345256 2295
rect 345204 2252 345256 2261
rect 347044 2295 347096 2304
rect 347044 2261 347053 2295
rect 347053 2261 347087 2295
rect 347087 2261 347096 2295
rect 347044 2252 347096 2261
rect 352196 2295 352248 2304
rect 352196 2261 352205 2295
rect 352205 2261 352239 2295
rect 352239 2261 352248 2295
rect 352196 2252 352248 2261
rect 357992 2320 358044 2372
rect 360660 2388 360712 2440
rect 365260 2431 365312 2440
rect 365260 2397 365269 2431
rect 365269 2397 365303 2431
rect 365303 2397 365312 2431
rect 365260 2388 365312 2397
rect 368388 2388 368440 2440
rect 370964 2388 371016 2440
rect 376116 2388 376168 2440
rect 378140 2431 378192 2440
rect 378140 2397 378149 2431
rect 378149 2397 378183 2431
rect 378183 2397 378192 2431
rect 378140 2388 378192 2397
rect 381268 2388 381320 2440
rect 383936 2388 383988 2440
rect 386420 2388 386472 2440
rect 388996 2388 389048 2440
rect 391572 2388 391624 2440
rect 393320 2388 393372 2440
rect 394148 2431 394200 2440
rect 394148 2397 394157 2431
rect 394157 2397 394191 2431
rect 394191 2397 394200 2431
rect 394148 2388 394200 2397
rect 396724 2431 396776 2440
rect 396724 2397 396733 2431
rect 396733 2397 396767 2431
rect 396767 2397 396776 2431
rect 396724 2388 396776 2397
rect 400312 2456 400364 2508
rect 398748 2431 398800 2440
rect 398748 2397 398757 2431
rect 398757 2397 398791 2431
rect 398791 2397 398800 2431
rect 398748 2388 398800 2397
rect 404360 2388 404412 2440
rect 357348 2295 357400 2304
rect 357348 2261 357357 2295
rect 357357 2261 357391 2295
rect 357391 2261 357400 2295
rect 357348 2252 357400 2261
rect 358084 2295 358136 2304
rect 358084 2261 358093 2295
rect 358093 2261 358127 2295
rect 358127 2261 358136 2295
rect 358084 2252 358136 2261
rect 359924 2295 359976 2304
rect 359924 2261 359933 2295
rect 359933 2261 359967 2295
rect 359967 2261 359976 2295
rect 359924 2252 359976 2261
rect 367100 2252 367152 2304
rect 368388 2295 368440 2304
rect 368388 2261 368397 2295
rect 368397 2261 368431 2295
rect 368431 2261 368440 2295
rect 368388 2252 368440 2261
rect 370964 2295 371016 2304
rect 370964 2261 370973 2295
rect 370973 2261 371007 2295
rect 371007 2261 371016 2295
rect 370964 2252 371016 2261
rect 376392 2252 376444 2304
rect 377956 2295 378008 2304
rect 377956 2261 377965 2295
rect 377965 2261 377999 2295
rect 377999 2261 378008 2295
rect 377956 2252 378008 2261
rect 381084 2252 381136 2304
rect 381268 2295 381320 2304
rect 381268 2261 381277 2295
rect 381277 2261 381311 2295
rect 381311 2261 381320 2295
rect 381268 2252 381320 2261
rect 383108 2295 383160 2304
rect 383108 2261 383117 2295
rect 383117 2261 383151 2295
rect 383151 2261 383160 2295
rect 383108 2252 383160 2261
rect 383200 2252 383252 2304
rect 383752 2252 383804 2304
rect 383936 2252 383988 2304
rect 386420 2295 386472 2304
rect 386420 2261 386429 2295
rect 386429 2261 386463 2295
rect 386463 2261 386472 2295
rect 386420 2252 386472 2261
rect 388996 2295 389048 2304
rect 388996 2261 389005 2295
rect 389005 2261 389039 2295
rect 389039 2261 389048 2295
rect 388996 2252 389048 2261
rect 391572 2295 391624 2304
rect 391572 2261 391581 2295
rect 391581 2261 391615 2295
rect 391615 2261 391624 2295
rect 391572 2252 391624 2261
rect 403992 2320 404044 2372
rect 446588 2592 446640 2644
rect 450820 2635 450872 2644
rect 450820 2601 450829 2635
rect 450829 2601 450863 2635
rect 450863 2601 450872 2635
rect 450820 2592 450872 2601
rect 414756 2567 414808 2576
rect 414756 2533 414765 2567
rect 414765 2533 414799 2567
rect 414799 2533 414808 2567
rect 414756 2524 414808 2533
rect 419908 2567 419960 2576
rect 419908 2533 419917 2567
rect 419917 2533 419951 2567
rect 419951 2533 419960 2567
rect 419908 2524 419960 2533
rect 417332 2388 417384 2440
rect 422484 2388 422536 2440
rect 426164 2524 426216 2576
rect 430212 2567 430264 2576
rect 430212 2533 430221 2567
rect 430221 2533 430255 2567
rect 430255 2533 430264 2567
rect 430212 2524 430264 2533
rect 431776 2524 431828 2576
rect 435364 2567 435416 2576
rect 435364 2533 435373 2567
rect 435373 2533 435407 2567
rect 435407 2533 435416 2567
rect 435364 2524 435416 2533
rect 436836 2524 436888 2576
rect 427636 2388 427688 2440
rect 432788 2388 432840 2440
rect 445668 2499 445720 2508
rect 445668 2465 445677 2499
rect 445677 2465 445711 2499
rect 445711 2465 445720 2499
rect 445668 2456 445720 2465
rect 440240 2320 440292 2372
rect 450820 2388 450872 2440
rect 464528 2592 464580 2644
rect 455420 2524 455472 2576
rect 459560 2456 459612 2508
rect 455972 2431 456024 2440
rect 455972 2397 455981 2431
rect 455981 2397 456015 2431
rect 456015 2397 456024 2431
rect 455972 2388 456024 2397
rect 466092 2524 466144 2576
rect 463700 2388 463752 2440
rect 483572 2592 483624 2644
rect 484308 2635 484360 2644
rect 484308 2601 484317 2635
rect 484317 2601 484351 2635
rect 484351 2601 484360 2635
rect 484308 2592 484360 2601
rect 466368 2524 466420 2576
rect 483020 2524 483072 2576
rect 468852 2388 468904 2440
rect 471428 2388 471480 2440
rect 473912 2388 473964 2440
rect 481640 2456 481692 2508
rect 481732 2499 481784 2508
rect 481732 2465 481741 2499
rect 481741 2465 481775 2499
rect 481775 2465 481784 2499
rect 481732 2456 481784 2465
rect 488540 2456 488592 2508
rect 475384 2320 475436 2372
rect 484308 2388 484360 2440
rect 485780 2388 485832 2440
rect 488724 2388 488776 2440
rect 491024 2388 491076 2440
rect 493600 2388 493652 2440
rect 496176 2388 496228 2440
rect 498752 2388 498804 2440
rect 501328 2388 501380 2440
rect 503904 2388 503956 2440
rect 506480 2388 506532 2440
rect 509056 2388 509108 2440
rect 511632 2388 511684 2440
rect 514208 2388 514260 2440
rect 484952 2320 485004 2372
rect 398840 2252 398892 2304
rect 402428 2252 402480 2304
rect 405924 2252 405976 2304
rect 406292 2295 406344 2304
rect 406292 2261 406301 2295
rect 406301 2261 406335 2295
rect 406335 2261 406344 2295
rect 406292 2252 406344 2261
rect 407028 2295 407080 2304
rect 407028 2261 407037 2295
rect 407037 2261 407071 2295
rect 407071 2261 407080 2295
rect 407028 2252 407080 2261
rect 408868 2295 408920 2304
rect 408868 2261 408877 2295
rect 408877 2261 408911 2295
rect 408911 2261 408920 2295
rect 408868 2252 408920 2261
rect 409604 2295 409656 2304
rect 409604 2261 409613 2295
rect 409613 2261 409647 2295
rect 409647 2261 409656 2295
rect 409604 2252 409656 2261
rect 411444 2295 411496 2304
rect 411444 2261 411453 2295
rect 411453 2261 411487 2295
rect 411487 2261 411496 2295
rect 411444 2252 411496 2261
rect 414020 2295 414072 2304
rect 414020 2261 414029 2295
rect 414029 2261 414063 2295
rect 414063 2261 414072 2295
rect 414020 2252 414072 2261
rect 416504 2252 416556 2304
rect 417332 2295 417384 2304
rect 417332 2261 417341 2295
rect 417341 2261 417375 2295
rect 417375 2261 417384 2295
rect 417332 2252 417384 2261
rect 419172 2295 419224 2304
rect 419172 2261 419181 2295
rect 419181 2261 419215 2295
rect 419215 2261 419224 2295
rect 419172 2252 419224 2261
rect 421748 2295 421800 2304
rect 421748 2261 421757 2295
rect 421757 2261 421791 2295
rect 421791 2261 421800 2295
rect 421748 2252 421800 2261
rect 422484 2295 422536 2304
rect 422484 2261 422493 2295
rect 422493 2261 422527 2295
rect 422527 2261 422536 2295
rect 422484 2252 422536 2261
rect 423588 2252 423640 2304
rect 426072 2252 426124 2304
rect 427636 2295 427688 2304
rect 427636 2261 427645 2295
rect 427645 2261 427679 2295
rect 427679 2261 427688 2295
rect 427636 2252 427688 2261
rect 427728 2252 427780 2304
rect 430488 2252 430540 2304
rect 432788 2295 432840 2304
rect 432788 2261 432797 2295
rect 432797 2261 432831 2295
rect 432831 2261 432840 2295
rect 432788 2252 432840 2261
rect 434628 2252 434680 2304
rect 440516 2295 440568 2304
rect 440516 2261 440525 2295
rect 440525 2261 440559 2295
rect 440559 2261 440568 2295
rect 440516 2252 440568 2261
rect 442356 2295 442408 2304
rect 442356 2261 442365 2295
rect 442365 2261 442399 2295
rect 442399 2261 442408 2295
rect 442356 2252 442408 2261
rect 443092 2295 443144 2304
rect 443092 2261 443101 2295
rect 443101 2261 443135 2295
rect 443135 2261 443144 2295
rect 443092 2252 443144 2261
rect 444380 2252 444432 2304
rect 445760 2252 445812 2304
rect 448244 2295 448296 2304
rect 448244 2261 448253 2295
rect 448253 2261 448287 2295
rect 448287 2261 448296 2295
rect 448244 2252 448296 2261
rect 448520 2252 448572 2304
rect 451372 2252 451424 2304
rect 453396 2252 453448 2304
rect 460388 2295 460440 2304
rect 460388 2261 460397 2295
rect 460397 2261 460431 2295
rect 460431 2261 460440 2295
rect 460388 2252 460440 2261
rect 462320 2252 462372 2304
rect 463700 2295 463752 2304
rect 463700 2261 463709 2295
rect 463709 2261 463743 2295
rect 463743 2261 463752 2295
rect 463700 2252 463752 2261
rect 463792 2252 463844 2304
rect 466460 2252 466512 2304
rect 468852 2295 468904 2304
rect 468852 2261 468861 2295
rect 468861 2261 468895 2295
rect 468895 2261 468904 2295
rect 468852 2252 468904 2261
rect 469220 2252 469272 2304
rect 471428 2295 471480 2304
rect 471428 2261 471437 2295
rect 471437 2261 471471 2295
rect 471471 2261 471480 2295
rect 471428 2252 471480 2261
rect 471888 2252 471940 2304
rect 473912 2295 473964 2304
rect 473912 2261 473921 2295
rect 473921 2261 473955 2295
rect 473955 2261 473964 2295
rect 473912 2252 473964 2261
rect 474004 2252 474056 2304
rect 475936 2252 475988 2304
rect 478512 2252 478564 2304
rect 483572 2295 483624 2304
rect 483572 2261 483581 2295
rect 483581 2261 483615 2295
rect 483615 2261 483624 2295
rect 483572 2252 483624 2261
rect 486148 2295 486200 2304
rect 486148 2261 486157 2295
rect 486157 2261 486191 2295
rect 486191 2261 486200 2295
rect 486148 2252 486200 2261
rect 488724 2295 488776 2304
rect 488724 2261 488733 2295
rect 488733 2261 488767 2295
rect 488767 2261 488776 2295
rect 488724 2252 488776 2261
rect 491300 2295 491352 2304
rect 491300 2261 491309 2295
rect 491309 2261 491343 2295
rect 491343 2261 491352 2295
rect 491300 2252 491352 2261
rect 493876 2295 493928 2304
rect 493876 2261 493885 2295
rect 493885 2261 493919 2295
rect 493919 2261 493928 2295
rect 493876 2252 493928 2261
rect 496452 2295 496504 2304
rect 496452 2261 496461 2295
rect 496461 2261 496495 2295
rect 496495 2261 496504 2295
rect 496452 2252 496504 2261
rect 498200 2252 498252 2304
rect 500316 2252 500368 2304
rect 502340 2252 502392 2304
rect 505100 2252 505152 2304
rect 509332 2295 509384 2304
rect 509332 2261 509341 2295
rect 509341 2261 509375 2295
rect 509375 2261 509384 2295
rect 509332 2252 509384 2261
rect 510528 2252 510580 2304
rect 67574 2150 67626 2202
rect 67638 2150 67690 2202
rect 67702 2150 67754 2202
rect 67766 2150 67818 2202
rect 67830 2150 67882 2202
rect 199502 2150 199554 2202
rect 199566 2150 199618 2202
rect 199630 2150 199682 2202
rect 199694 2150 199746 2202
rect 199758 2150 199810 2202
rect 331430 2150 331482 2202
rect 331494 2150 331546 2202
rect 331558 2150 331610 2202
rect 331622 2150 331674 2202
rect 331686 2150 331738 2202
rect 463358 2150 463410 2202
rect 463422 2150 463474 2202
rect 463486 2150 463538 2202
rect 463550 2150 463602 2202
rect 463614 2150 463666 2202
rect 37924 2048 37976 2100
rect 98644 2048 98696 2100
rect 99748 2048 99800 2100
rect 127716 2048 127768 2100
rect 127992 2048 128044 2100
rect 136456 2048 136508 2100
rect 143448 2048 143500 2100
rect 191104 2048 191156 2100
rect 195060 2048 195112 2100
rect 263140 2048 263192 2100
rect 340052 2048 340104 2100
rect 30196 1980 30248 2032
rect 48780 1980 48832 2032
rect 53380 1980 53432 2032
rect 108672 1980 108724 2032
rect 108764 1980 108816 2032
rect 130660 1980 130712 2032
rect 139124 1980 139176 2032
rect 143080 1980 143132 2032
rect 152004 1980 152056 2032
rect 195612 1980 195664 2032
rect 200212 1980 200264 2032
rect 264336 1980 264388 2032
rect 342628 1980 342680 2032
rect 377956 2048 378008 2100
rect 383292 2048 383344 2100
rect 383936 2048 383988 2100
rect 397368 2048 397420 2100
rect 409604 2048 409656 2100
rect 443736 2048 443788 2100
rect 475384 2048 475436 2100
rect 482744 2048 482796 2100
rect 35348 1912 35400 1964
rect 56508 1912 56560 1964
rect 58532 1912 58584 1964
rect 115480 1912 115532 1964
rect 122932 1912 122984 1964
rect 141700 1912 141752 1964
rect 157156 1912 157208 1964
rect 196072 1912 196124 1964
rect 215668 1912 215720 1964
rect 268384 1912 268436 1964
rect 302332 1912 302384 1964
rect 321284 1912 321336 1964
rect 329748 1912 329800 1964
rect 365628 1912 365680 1964
rect 66720 1844 66772 1896
rect 70400 1844 70452 1896
rect 74908 1844 74960 1896
rect 78680 1844 78732 1896
rect 80244 1844 80296 1896
rect 89812 1844 89864 1896
rect 91836 1844 91888 1896
rect 102140 1844 102192 1896
rect 102232 1844 102284 1896
rect 107936 1844 107988 1896
rect 14740 1776 14792 1828
rect 96804 1776 96856 1828
rect 97448 1776 97500 1828
rect 115296 1844 115348 1896
rect 120356 1844 120408 1896
rect 143172 1844 143224 1896
rect 148968 1844 149020 1896
rect 157248 1844 157300 1896
rect 158996 1844 159048 1896
rect 109224 1776 109276 1828
rect 125508 1776 125560 1828
rect 130844 1776 130896 1828
rect 148140 1776 148192 1828
rect 7012 1708 7064 1760
rect 75552 1708 75604 1760
rect 75644 1708 75696 1760
rect 80152 1708 80204 1760
rect 80336 1708 80388 1760
rect 86960 1708 87012 1760
rect 87052 1708 87104 1760
rect 92296 1708 92348 1760
rect 25044 1640 25096 1692
rect 99564 1708 99616 1760
rect 94596 1640 94648 1692
rect 103428 1708 103480 1760
rect 107476 1708 107528 1760
rect 114928 1708 114980 1760
rect 118700 1708 118752 1760
rect 127624 1708 127676 1760
rect 128176 1708 128228 1760
rect 132592 1708 132644 1760
rect 50804 1572 50856 1624
rect 111984 1640 112036 1692
rect 112812 1640 112864 1692
rect 121460 1640 121512 1692
rect 121736 1640 121788 1692
rect 132500 1640 132552 1692
rect 104900 1572 104952 1624
rect 110788 1572 110840 1624
rect 115204 1572 115256 1624
rect 141056 1708 141108 1760
rect 145840 1708 145892 1760
rect 161940 1776 161992 1828
rect 162308 1844 162360 1896
rect 196716 1844 196768 1896
rect 220820 1844 220872 1896
rect 269672 1844 269724 1896
rect 358084 1844 358136 1896
rect 163688 1776 163740 1828
rect 148508 1708 148560 1760
rect 158536 1708 158588 1760
rect 161204 1708 161256 1760
rect 163964 1776 164016 1828
rect 167460 1776 167512 1828
rect 198740 1776 198792 1828
rect 225972 1776 226024 1828
rect 270592 1776 270644 1828
rect 352196 1776 352248 1828
rect 359832 1776 359884 1828
rect 383108 1980 383160 2032
rect 387800 1980 387852 2032
rect 391572 1980 391624 2032
rect 420920 1980 420972 2032
rect 422484 1980 422536 2032
rect 447692 1980 447744 2032
rect 463700 1980 463752 2032
rect 481824 1980 481876 2032
rect 382280 1912 382332 1964
rect 383752 1912 383804 1964
rect 392032 1912 392084 1964
rect 417332 1912 417384 1964
rect 447140 1912 447192 1964
rect 471428 1912 471480 1964
rect 484124 1912 484176 1964
rect 443092 1844 443144 1896
rect 481180 1844 481232 1896
rect 133972 1640 134024 1692
rect 172520 1708 172572 1760
rect 172612 1708 172664 1760
rect 186872 1708 186924 1760
rect 188344 1708 188396 1760
rect 192944 1708 192996 1760
rect 163964 1640 164016 1692
rect 168104 1640 168156 1692
rect 168288 1640 168340 1692
rect 185492 1640 185544 1692
rect 185860 1640 185912 1692
rect 195980 1708 196032 1760
rect 337476 1708 337528 1760
rect 372804 1708 372856 1760
rect 378692 1776 378744 1828
rect 388996 1776 389048 1828
rect 432052 1776 432104 1828
rect 468852 1776 468904 1828
rect 480260 1776 480312 1828
rect 381544 1708 381596 1760
rect 394148 1708 394200 1760
rect 440148 1708 440200 1760
rect 440516 1708 440568 1760
rect 475292 1708 475344 1760
rect 282368 1640 282420 1692
rect 291200 1640 291252 1692
rect 314292 1640 314344 1692
rect 361580 1640 361632 1692
rect 368388 1640 368440 1692
rect 400404 1640 400456 1692
rect 427636 1640 427688 1692
rect 445576 1640 445628 1692
rect 448244 1640 448296 1692
rect 477500 1640 477552 1692
rect 137008 1572 137060 1624
rect 138112 1572 138164 1624
rect 848 756 900 808
rect 1308 756 1360 808
rect 4160 824 4212 876
rect 3976 756 4028 808
rect 6000 824 6052 876
rect 6184 756 6236 808
rect 6736 756 6788 808
rect 8484 756 8536 808
rect 9588 756 9640 808
rect 11336 824 11388 876
rect 14280 1096 14332 1148
rect 10784 688 10836 740
rect 17316 960 17368 1012
rect 16580 892 16632 944
rect 19248 1300 19300 1352
rect 29092 1300 29144 1352
rect 20720 1232 20772 1284
rect 24768 1232 24820 1284
rect 28264 1232 28316 1284
rect 33508 1300 33560 1352
rect 38660 1300 38712 1352
rect 34796 1232 34848 1284
rect 35716 1232 35768 1284
rect 42800 1368 42852 1420
rect 42156 1300 42208 1352
rect 50528 1436 50580 1488
rect 51908 1436 51960 1488
rect 57888 1436 57940 1488
rect 43260 1232 43312 1284
rect 49700 1368 49752 1420
rect 49056 1300 49108 1352
rect 53840 1368 53892 1420
rect 60556 1368 60608 1420
rect 63684 1504 63736 1556
rect 69480 1504 69532 1556
rect 74540 1504 74592 1556
rect 75736 1504 75788 1556
rect 81532 1504 81584 1556
rect 84292 1504 84344 1556
rect 118700 1504 118752 1556
rect 118792 1504 118844 1556
rect 124220 1504 124272 1556
rect 62764 1436 62816 1488
rect 64880 1436 64932 1488
rect 66260 1436 66312 1488
rect 118884 1436 118936 1488
rect 119620 1436 119672 1488
rect 125692 1436 125744 1488
rect 126152 1436 126204 1488
rect 126980 1436 127032 1488
rect 128084 1436 128136 1488
rect 132224 1436 132276 1488
rect 56140 1300 56192 1352
rect 60648 1300 60700 1352
rect 60740 1300 60792 1352
rect 67916 1368 67968 1420
rect 66168 1300 66220 1352
rect 71504 1300 71556 1352
rect 73344 1300 73396 1352
rect 49792 1232 49844 1284
rect 53748 1232 53800 1284
rect 15936 756 15988 808
rect 21640 1164 21692 1216
rect 23940 1096 23992 1148
rect 23848 1028 23900 1080
rect 27620 1164 27672 1216
rect 28908 1164 28960 1216
rect 24860 824 24912 876
rect 32772 1096 32824 1148
rect 37832 1096 37884 1148
rect 44088 1096 44140 1148
rect 24768 756 24820 808
rect 29368 892 29420 944
rect 31852 960 31904 1012
rect 37464 1028 37516 1080
rect 29092 756 29144 808
rect 33140 892 33192 944
rect 36820 892 36872 944
rect 39120 1028 39172 1080
rect 40868 1028 40920 1080
rect 43168 1028 43220 1080
rect 33508 688 33560 740
rect 35716 756 35768 808
rect 37832 756 37884 808
rect 41328 960 41380 1012
rect 46020 960 46072 1012
rect 53564 1164 53616 1216
rect 56232 1232 56284 1284
rect 58992 1232 59044 1284
rect 59636 1232 59688 1284
rect 63224 1232 63276 1284
rect 47676 1096 47728 1148
rect 48964 1096 49016 1148
rect 49056 1096 49108 1148
rect 57980 1164 58032 1216
rect 58532 1164 58584 1216
rect 62764 1164 62816 1216
rect 54024 1096 54076 1148
rect 56692 1096 56744 1148
rect 57428 1096 57480 1148
rect 68560 1232 68612 1284
rect 63592 1164 63644 1216
rect 66720 1164 66772 1216
rect 66812 1164 66864 1216
rect 69480 1164 69532 1216
rect 63960 1096 64012 1148
rect 73436 1232 73488 1284
rect 69664 1164 69716 1216
rect 73620 1368 73672 1420
rect 74908 1300 74960 1352
rect 75000 1300 75052 1352
rect 86776 1368 86828 1420
rect 94136 1368 94188 1420
rect 78036 1300 78088 1352
rect 89720 1300 89772 1352
rect 89812 1300 89864 1352
rect 92572 1300 92624 1352
rect 95516 1300 95568 1352
rect 99012 1300 99064 1352
rect 73620 1232 73672 1284
rect 75460 1232 75512 1284
rect 77208 1232 77260 1284
rect 79140 1232 79192 1284
rect 80152 1232 80204 1284
rect 84108 1232 84160 1284
rect 85764 1232 85816 1284
rect 70492 1096 70544 1148
rect 87052 1164 87104 1216
rect 89904 1232 89956 1284
rect 99104 1232 99156 1284
rect 105268 1368 105320 1420
rect 107752 1368 107804 1420
rect 101128 1300 101180 1352
rect 110328 1368 110380 1420
rect 110788 1368 110840 1420
rect 136180 1504 136232 1556
rect 132500 1436 132552 1488
rect 144736 1572 144788 1624
rect 146208 1572 146260 1624
rect 148508 1572 148560 1624
rect 148600 1572 148652 1624
rect 252468 1572 252520 1624
rect 262404 1572 262456 1624
rect 264980 1572 265032 1624
rect 278228 1572 278280 1624
rect 283104 1572 283156 1624
rect 345204 1572 345256 1624
rect 389180 1572 389232 1624
rect 396724 1572 396776 1624
rect 440976 1572 441028 1624
rect 473912 1572 473964 1624
rect 484216 1572 484268 1624
rect 141424 1504 141476 1556
rect 148232 1504 148284 1556
rect 150348 1504 150400 1556
rect 161572 1504 161624 1556
rect 161756 1504 161808 1556
rect 166816 1504 166868 1556
rect 167460 1504 167512 1556
rect 174636 1504 174688 1556
rect 174820 1504 174872 1556
rect 179512 1504 179564 1556
rect 179604 1504 179656 1556
rect 259920 1504 259972 1556
rect 273996 1504 274048 1556
rect 282276 1504 282328 1556
rect 282552 1504 282604 1556
rect 285680 1504 285732 1556
rect 293500 1504 293552 1556
rect 300860 1504 300912 1556
rect 324596 1504 324648 1556
rect 372620 1504 372672 1556
rect 381268 1504 381320 1556
rect 417056 1504 417108 1556
rect 432788 1504 432840 1556
rect 456800 1504 456852 1556
rect 143724 1436 143776 1488
rect 147772 1436 147824 1488
rect 147864 1436 147916 1488
rect 153384 1436 153436 1488
rect 154580 1436 154632 1488
rect 156420 1436 156472 1488
rect 132592 1368 132644 1420
rect 144920 1368 144972 1420
rect 146668 1368 146720 1420
rect 157432 1368 157484 1420
rect 166724 1368 166776 1420
rect 166816 1368 166868 1420
rect 167000 1368 167052 1420
rect 168656 1436 168708 1488
rect 176752 1436 176804 1488
rect 176936 1436 176988 1488
rect 181076 1436 181128 1488
rect 181352 1436 181404 1488
rect 182180 1436 182232 1488
rect 109040 1300 109092 1352
rect 113180 1300 113232 1352
rect 113640 1300 113692 1352
rect 183652 1368 183704 1420
rect 186688 1436 186740 1488
rect 188344 1436 188396 1488
rect 190184 1436 190236 1488
rect 195244 1436 195296 1488
rect 195336 1436 195388 1488
rect 262312 1436 262364 1488
rect 271604 1436 271656 1488
rect 273352 1436 273404 1488
rect 282920 1436 282972 1488
rect 295248 1436 295300 1488
rect 302516 1436 302568 1488
rect 306380 1436 306432 1488
rect 313372 1436 313424 1488
rect 316684 1436 316736 1488
rect 319444 1436 319496 1488
rect 367928 1436 367980 1488
rect 370964 1436 371016 1488
rect 395436 1436 395488 1488
rect 407028 1436 407080 1488
rect 442908 1436 442960 1488
rect 249524 1368 249576 1420
rect 183812 1300 183864 1352
rect 184020 1300 184072 1352
rect 208216 1300 208268 1352
rect 219624 1300 219676 1352
rect 226064 1300 226116 1352
rect 228456 1300 228508 1352
rect 233240 1300 233292 1352
rect 234988 1300 235040 1352
rect 244004 1300 244056 1352
rect 254952 1368 255004 1420
rect 261208 1368 261260 1420
rect 106372 1232 106424 1284
rect 106556 1232 106608 1284
rect 118700 1232 118752 1284
rect 89812 1164 89864 1216
rect 47860 1028 47912 1080
rect 48044 960 48096 1012
rect 52736 960 52788 1012
rect 52644 892 52696 944
rect 40868 756 40920 808
rect 42156 756 42208 808
rect 43260 756 43312 808
rect 47676 756 47728 808
rect 48872 824 48924 876
rect 49792 756 49844 808
rect 51908 824 51960 876
rect 59360 1028 59412 1080
rect 61844 1028 61896 1080
rect 60556 960 60608 1012
rect 63224 960 63276 1012
rect 56140 892 56192 944
rect 56232 824 56284 876
rect 63500 892 63552 944
rect 65064 960 65116 1012
rect 68100 960 68152 1012
rect 68284 1028 68336 1080
rect 73160 1028 73212 1080
rect 75736 1096 75788 1148
rect 75828 1096 75880 1148
rect 81348 1096 81400 1148
rect 75644 1028 75696 1080
rect 68468 960 68520 1012
rect 69848 960 69900 1012
rect 71780 960 71832 1012
rect 72884 960 72936 1012
rect 80060 1028 80112 1080
rect 84476 1096 84528 1148
rect 84660 1096 84712 1148
rect 82452 1028 82504 1080
rect 86868 1028 86920 1080
rect 71412 892 71464 944
rect 58992 824 59044 876
rect 65248 824 65300 876
rect 68744 824 68796 876
rect 57428 688 57480 740
rect 58532 756 58584 808
rect 59636 688 59688 740
rect 60740 756 60792 808
rect 61844 756 61896 808
rect 62856 688 62908 740
rect 63960 756 64012 808
rect 65064 756 65116 808
rect 66168 756 66220 808
rect 66812 756 66864 808
rect 68284 756 68336 808
rect 69388 688 69440 740
rect 70492 688 70544 740
rect 71504 756 71556 808
rect 72884 824 72936 876
rect 73068 892 73120 944
rect 73160 824 73212 876
rect 75828 824 75880 876
rect 75000 8 75052 60
rect 75736 756 75788 808
rect 80336 892 80388 944
rect 76564 824 76616 876
rect 81440 892 81492 944
rect 86960 960 87012 1012
rect 87880 1028 87932 1080
rect 99196 1164 99248 1216
rect 100024 1164 100076 1216
rect 110696 1164 110748 1216
rect 110788 1164 110840 1216
rect 112812 1164 112864 1216
rect 113088 1164 113140 1216
rect 93308 1096 93360 1148
rect 108856 1096 108908 1148
rect 108948 1096 109000 1148
rect 113640 1096 113692 1148
rect 113824 1164 113876 1216
rect 115020 1164 115072 1216
rect 115112 1164 115164 1216
rect 126888 1232 126940 1284
rect 126980 1232 127032 1284
rect 133144 1232 133196 1284
rect 133236 1232 133288 1284
rect 123576 1164 123628 1216
rect 126152 1164 126204 1216
rect 126244 1164 126296 1216
rect 137744 1164 137796 1216
rect 141424 1232 141476 1284
rect 141516 1232 141568 1284
rect 146484 1232 146536 1284
rect 147772 1232 147824 1284
rect 151268 1232 151320 1284
rect 139308 1164 139360 1216
rect 147864 1164 147916 1216
rect 148140 1164 148192 1216
rect 151360 1164 151412 1216
rect 92204 1028 92256 1080
rect 94320 1028 94372 1080
rect 94688 1028 94740 1080
rect 90180 960 90232 1012
rect 90272 960 90324 1012
rect 94136 960 94188 1012
rect 78036 756 78088 808
rect 79140 756 79192 808
rect 80244 756 80296 808
rect 82452 756 82504 808
rect 91284 892 91336 944
rect 91376 892 91428 944
rect 94320 892 94372 944
rect 84016 824 84068 876
rect 86914 824 86966 876
rect 84660 688 84712 740
rect 85764 756 85816 808
rect 86868 552 86920 604
rect 87880 756 87932 808
rect 87236 688 87288 740
rect 91836 824 91888 876
rect 89168 484 89220 536
rect 90088 756 90140 808
rect 91376 756 91428 808
rect 92204 756 92256 808
rect 93308 756 93360 808
rect 99380 960 99432 1012
rect 102508 1028 102560 1080
rect 104164 1028 104216 1080
rect 110788 1028 110840 1080
rect 110880 1028 110932 1080
rect 113824 1028 113876 1080
rect 113916 1028 113968 1080
rect 114560 1028 114612 1080
rect 100944 960 100996 1012
rect 113364 960 113416 1012
rect 115204 1096 115256 1148
rect 121736 1096 121788 1148
rect 122104 1096 122156 1148
rect 130752 1096 130804 1148
rect 132960 1096 133012 1148
rect 139216 1096 139268 1148
rect 139400 1096 139452 1148
rect 146392 1096 146444 1148
rect 148048 1096 148100 1148
rect 150348 1096 150400 1148
rect 150440 1096 150492 1148
rect 157156 1232 157208 1284
rect 157248 1232 157300 1284
rect 183514 1232 183566 1284
rect 186136 1232 186188 1284
rect 186412 1232 186464 1284
rect 244096 1232 244148 1284
rect 244372 1232 244424 1284
rect 247592 1232 247644 1284
rect 258080 1300 258132 1352
rect 258908 1300 258960 1352
rect 263416 1300 263468 1352
rect 267832 1368 267884 1420
rect 269856 1368 269908 1420
rect 274272 1368 274324 1420
rect 282644 1368 282696 1420
rect 283196 1368 283248 1420
rect 289912 1368 289964 1420
rect 295800 1368 295852 1420
rect 298192 1368 298244 1420
rect 300216 1368 300268 1420
rect 303528 1368 303580 1420
rect 306564 1368 306616 1420
rect 318708 1368 318760 1420
rect 332324 1368 332376 1420
rect 375564 1368 375616 1420
rect 386420 1368 386472 1420
rect 426992 1368 427044 1420
rect 360200 1300 360252 1352
rect 151544 1164 151596 1216
rect 156880 1164 156932 1216
rect 156972 1164 157024 1216
rect 167000 1164 167052 1216
rect 167092 1164 167144 1216
rect 176384 1164 176436 1216
rect 176568 1164 176620 1216
rect 152372 1096 152424 1148
rect 156788 1096 156840 1148
rect 158904 1096 158956 1148
rect 166724 1096 166776 1148
rect 166816 1096 166868 1148
rect 167184 1096 167236 1148
rect 168104 1096 168156 1148
rect 170864 1096 170916 1148
rect 170956 1096 171008 1148
rect 173256 1096 173308 1148
rect 173348 1096 173400 1148
rect 181628 1164 181680 1216
rect 183652 1164 183704 1216
rect 183836 1164 183888 1216
rect 115020 1028 115072 1080
rect 118608 1028 118660 1080
rect 118792 1028 118844 1080
rect 142712 1028 142764 1080
rect 115204 960 115256 1012
rect 116492 960 116544 1012
rect 94596 892 94648 944
rect 97540 892 97592 944
rect 95516 756 95568 808
rect 97448 824 97500 876
rect 113916 892 113968 944
rect 114008 892 114060 944
rect 128268 892 128320 944
rect 97908 416 97960 468
rect 98828 756 98880 808
rect 99748 756 99800 808
rect 100944 688 100996 740
rect 102048 756 102100 808
rect 103612 824 103664 876
rect 108304 824 108356 876
rect 104164 756 104216 808
rect 105268 756 105320 808
rect 106556 756 106608 808
rect 107476 756 107528 808
rect 108764 756 108816 808
rect 110880 756 110932 808
rect 111892 756 111944 808
rect 113088 756 113140 808
rect 119620 824 119672 876
rect 114008 620 114060 672
rect 113364 552 113416 604
rect 114192 552 114244 604
rect 116492 756 116544 808
rect 114744 688 114796 740
rect 123576 824 123628 876
rect 115388 620 115440 672
rect 118516 620 118568 672
rect 118608 620 118660 672
rect 119528 620 119580 672
rect 114468 552 114520 604
rect 119712 552 119764 604
rect 114928 484 114980 536
rect 118608 484 118660 536
rect 114744 416 114796 468
rect 117504 416 117556 468
rect 114560 212 114612 264
rect 119436 212 119488 264
rect 122104 756 122156 808
rect 127992 824 128044 876
rect 130476 824 130528 876
rect 126244 756 126296 808
rect 124496 212 124548 264
rect 126428 212 126480 264
rect 128176 756 128228 808
rect 133052 960 133104 1012
rect 133144 960 133196 1012
rect 131028 892 131080 944
rect 134892 960 134944 1012
rect 139308 960 139360 1012
rect 156696 1028 156748 1080
rect 157524 1028 157576 1080
rect 142896 960 142948 1012
rect 156972 960 157024 1012
rect 139492 892 139544 944
rect 146208 892 146260 944
rect 146484 892 146536 944
rect 148048 892 148100 944
rect 137008 824 137060 876
rect 126888 620 126940 672
rect 128360 620 128412 672
rect 132960 756 133012 808
rect 134892 756 134944 808
rect 137836 824 137888 876
rect 139124 824 139176 876
rect 139216 824 139268 876
rect 143724 824 143776 876
rect 139400 688 139452 740
rect 139308 552 139360 604
rect 141516 756 141568 808
rect 146300 824 146352 876
rect 150440 892 150492 944
rect 150532 892 150584 944
rect 154580 892 154632 944
rect 157340 960 157392 1012
rect 157432 960 157484 1012
rect 145840 620 145892 672
rect 146392 8 146444 60
rect 147956 8 148008 60
rect 152372 688 152424 740
rect 154580 756 154632 808
rect 159088 824 159140 876
rect 157156 552 157208 604
rect 158996 552 159048 604
rect 157248 484 157300 536
rect 158904 484 158956 536
rect 158996 416 159048 468
rect 161204 688 161256 740
rect 161756 756 161808 808
rect 164056 620 164108 672
rect 164332 620 164384 672
rect 166264 620 166316 672
rect 166264 484 166316 536
rect 167184 960 167236 1012
rect 171140 960 171192 1012
rect 172244 1028 172296 1080
rect 172336 1028 172388 1080
rect 176476 1028 176528 1080
rect 176752 1028 176804 1080
rect 181352 1028 181404 1080
rect 183928 1096 183980 1148
rect 184020 1096 184072 1148
rect 185860 1096 185912 1148
rect 168104 892 168156 944
rect 170956 892 171008 944
rect 168288 824 168340 876
rect 177488 960 177540 1012
rect 172244 892 172296 944
rect 176936 892 176988 944
rect 183514 960 183566 1012
rect 184112 1028 184164 1080
rect 185952 1028 186004 1080
rect 186228 1164 186280 1216
rect 213092 1164 213144 1216
rect 224316 1164 224368 1216
rect 186780 1096 186832 1148
rect 195060 1096 195112 1148
rect 186688 1028 186740 1080
rect 186872 1028 186924 1080
rect 215392 1096 215444 1148
rect 219716 1096 219768 1148
rect 223396 1096 223448 1148
rect 226432 1164 226484 1216
rect 236276 1164 236328 1216
rect 238484 1164 238536 1216
rect 243912 1164 243964 1216
rect 244648 1164 244700 1216
rect 255412 1232 255464 1284
rect 256884 1232 256936 1284
rect 267832 1232 267884 1284
rect 267924 1232 267976 1284
rect 282828 1232 282880 1284
rect 283012 1232 283064 1284
rect 372712 1300 372764 1352
rect 254768 1164 254820 1216
rect 268016 1164 268068 1216
rect 268660 1164 268712 1216
rect 273260 1164 273312 1216
rect 273352 1164 273404 1216
rect 276020 1164 276072 1216
rect 278044 1164 278096 1216
rect 282552 1164 282604 1216
rect 195244 1028 195296 1080
rect 220544 1028 220596 1080
rect 222108 1028 222160 1080
rect 229100 1028 229152 1080
rect 230572 1096 230624 1148
rect 233700 1028 233752 1080
rect 237288 1096 237340 1148
rect 241428 1028 241480 1080
rect 241520 1028 241572 1080
rect 242900 1028 242952 1080
rect 242992 1028 243044 1080
rect 244372 1028 244424 1080
rect 245752 1096 245804 1148
rect 253848 1096 253900 1148
rect 253940 1096 253992 1148
rect 267188 1096 267240 1148
rect 267740 1096 267792 1148
rect 282736 1096 282788 1148
rect 247040 1028 247092 1080
rect 248052 1028 248104 1080
rect 254952 1028 255004 1080
rect 255044 1028 255096 1080
rect 261208 1028 261260 1080
rect 261300 1028 261352 1080
rect 271604 1028 271656 1080
rect 271696 1028 271748 1080
rect 282460 1028 282512 1080
rect 283104 1028 283156 1080
rect 383016 1164 383068 1216
rect 287244 1096 287296 1148
rect 292212 1096 292264 1148
rect 292304 1096 292356 1148
rect 293500 1096 293552 1148
rect 287796 1028 287848 1080
rect 291016 1028 291068 1080
rect 291108 1028 291160 1080
rect 302516 1096 302568 1148
rect 304816 1096 304868 1148
rect 311900 1096 311952 1148
rect 311992 1096 312044 1148
rect 336740 1096 336792 1148
rect 365076 1096 365128 1148
rect 177948 892 178000 944
rect 181536 892 181588 944
rect 168196 756 168248 808
rect 166724 688 166776 740
rect 168288 688 168340 740
rect 166632 620 166684 672
rect 168472 552 168524 604
rect 166540 484 166592 536
rect 168104 484 168156 536
rect 171048 756 171100 808
rect 177672 824 177724 876
rect 178684 824 178736 876
rect 183652 892 183704 944
rect 185676 892 185728 944
rect 186872 892 186924 944
rect 187884 960 187936 1012
rect 218244 960 218296 1012
rect 166908 348 166960 400
rect 170404 484 170456 536
rect 172336 688 172388 740
rect 170864 620 170916 672
rect 172796 620 172848 672
rect 173348 756 173400 808
rect 173164 688 173216 740
rect 175004 688 175056 740
rect 173072 552 173124 604
rect 173992 552 174044 604
rect 173256 8 173308 60
rect 174820 8 174872 60
rect 177028 756 177080 808
rect 183928 824 183980 876
rect 198740 892 198792 944
rect 228548 960 228600 1012
rect 231676 960 231728 1012
rect 219532 892 219584 944
rect 239128 892 239180 944
rect 239404 960 239456 1012
rect 262404 960 262456 1012
rect 262496 960 262548 1012
rect 239956 892 240008 944
rect 181260 552 181312 604
rect 179788 144 179840 196
rect 181260 144 181312 196
rect 183514 756 183566 808
rect 181904 552 181956 604
rect 183560 552 183612 604
rect 181904 144 181956 196
rect 183652 144 183704 196
rect 185676 756 185728 808
rect 187884 688 187936 740
rect 190184 756 190236 808
rect 192208 280 192260 332
rect 194600 620 194652 672
rect 192852 484 192904 536
rect 194324 484 194376 536
rect 195244 824 195296 876
rect 198004 824 198056 876
rect 219624 824 219676 876
rect 241612 892 241664 944
rect 241704 892 241756 944
rect 245752 892 245804 944
rect 246028 892 246080 944
rect 247592 892 247644 944
rect 194968 756 195020 808
rect 196348 756 196400 808
rect 212080 756 212132 808
rect 241980 824 242032 876
rect 250812 892 250864 944
rect 253756 892 253808 944
rect 274088 960 274140 1012
rect 276480 960 276532 1012
rect 282368 960 282420 1012
rect 282828 960 282880 1012
rect 254124 824 254176 876
rect 265440 892 265492 944
rect 267832 892 267884 944
rect 195152 620 195204 672
rect 194968 552 195020 604
rect 195980 552 196032 604
rect 196072 552 196124 604
rect 219532 620 219584 672
rect 195060 484 195112 536
rect 196348 484 196400 536
rect 194876 416 194928 468
rect 198004 416 198056 468
rect 192944 76 192996 128
rect 194600 76 194652 128
rect 192852 8 192904 60
rect 194508 8 194560 60
rect 198740 348 198792 400
rect 195244 280 195296 332
rect 202788 280 202840 332
rect 194968 212 195020 264
rect 210240 212 210292 264
rect 195980 144 196032 196
rect 207940 144 207992 196
rect 194784 76 194836 128
rect 205088 76 205140 128
rect 194876 8 194928 60
rect 219716 8 219768 60
rect 222108 756 222160 808
rect 224316 756 224368 808
rect 226432 756 226484 808
rect 228456 756 228508 808
rect 230572 756 230624 808
rect 231676 756 231728 808
rect 234988 756 235040 808
rect 237288 756 237340 808
rect 238484 756 238536 808
rect 241704 756 241756 808
rect 239956 688 240008 740
rect 241520 688 241572 740
rect 242992 756 243044 808
rect 246028 620 246080 672
rect 248052 756 248104 808
rect 250352 144 250404 196
rect 250812 620 250864 672
rect 250628 212 250680 264
rect 252560 212 252612 264
rect 254768 620 254820 672
rect 256884 756 256936 808
rect 258908 756 258960 808
rect 261300 756 261352 808
rect 259368 416 259420 468
rect 260840 416 260892 468
rect 262496 756 262548 808
rect 265624 824 265676 876
rect 265900 824 265952 876
rect 273168 892 273220 944
rect 273352 892 273404 944
rect 268200 824 268252 876
rect 274272 824 274324 876
rect 278044 892 278096 944
rect 274824 824 274876 876
rect 278596 892 278648 944
rect 278688 892 278740 944
rect 278964 824 279016 876
rect 280344 824 280396 876
rect 280896 892 280948 944
rect 283012 892 283064 944
rect 283196 892 283248 944
rect 282920 824 282972 876
rect 263416 756 263468 808
rect 265440 620 265492 672
rect 267740 688 267792 740
rect 268660 688 268712 740
rect 271696 756 271748 808
rect 273996 688 274048 740
rect 276480 756 276532 808
rect 278596 756 278648 808
rect 280896 552 280948 604
rect 282828 756 282880 808
rect 287796 824 287848 876
rect 287244 756 287296 808
rect 289544 824 289596 876
rect 289728 892 289780 944
rect 293868 960 293920 1012
rect 302700 1028 302752 1080
rect 306932 1028 306984 1080
rect 297548 960 297600 1012
rect 300216 960 300268 1012
rect 300400 960 300452 1012
rect 291752 824 291804 876
rect 291108 756 291160 808
rect 295800 892 295852 944
rect 302792 960 302844 1012
rect 315304 960 315356 1012
rect 316500 960 316552 1012
rect 293868 756 293920 808
rect 302332 824 302384 876
rect 306564 824 306616 876
rect 308128 892 308180 944
rect 334164 1028 334216 1080
rect 357992 1028 358044 1080
rect 362592 1028 362644 1080
rect 316868 960 316920 1012
rect 331220 960 331272 1012
rect 359924 960 359976 1012
rect 367100 1028 367152 1080
rect 316960 892 317012 944
rect 341892 892 341944 944
rect 357348 892 357400 944
rect 307208 824 307260 876
rect 307392 824 307444 876
rect 313372 824 313424 876
rect 293868 484 293920 536
rect 300400 756 300452 808
rect 298560 76 298612 128
rect 300400 76 300452 128
rect 302608 756 302660 808
rect 304816 756 304868 808
rect 306932 756 306984 808
rect 308128 756 308180 808
rect 311072 756 311124 808
rect 315672 756 315724 808
rect 315948 756 316000 808
rect 316960 756 317012 808
rect 339316 824 339368 876
rect 359832 824 359884 876
rect 376392 1096 376444 1148
rect 373540 1028 373592 1080
rect 355416 756 355468 808
rect 318064 212 318116 264
rect 329012 212 329064 264
rect 318248 144 318300 196
rect 326436 144 326488 196
rect 317880 8 317932 60
rect 347044 76 347096 128
rect 318064 8 318116 60
rect 344468 8 344520 60
rect 362592 756 362644 808
rect 442356 1028 442408 1080
rect 373448 756 373500 808
rect 380900 756 380952 808
rect 383844 756 383896 808
rect 385040 756 385092 808
rect 387800 756 387852 808
rect 390652 756 390704 808
rect 391940 756 391992 808
rect 394056 756 394108 808
rect 395252 756 395304 808
rect 397644 756 397696 808
rect 400220 756 400272 808
rect 402428 756 402480 808
rect 406292 756 406344 808
rect 405924 688 405976 740
rect 408868 756 408920 808
rect 411444 756 411496 808
rect 414020 756 414072 808
rect 416504 756 416556 808
rect 419172 756 419224 808
rect 421748 756 421800 808
rect 423588 756 423640 808
rect 426072 756 426124 808
rect 427728 756 427780 808
rect 430488 756 430540 808
rect 431776 756 431828 808
rect 434628 756 434680 808
rect 436836 756 436888 808
rect 444380 892 444432 944
rect 445760 824 445812 876
rect 448520 1232 448572 1284
rect 451372 1164 451424 1216
rect 460388 1300 460440 1352
rect 481548 1300 481600 1352
rect 491300 1300 491352 1352
rect 453396 1096 453448 1148
rect 455420 824 455472 876
rect 462320 1232 462372 1284
rect 470600 1232 470652 1284
rect 474004 1232 474056 1284
rect 485964 1232 486016 1284
rect 496452 1232 496504 1284
rect 463792 1164 463844 1216
rect 472900 1164 472952 1216
rect 478512 1164 478564 1216
rect 483756 1164 483808 1216
rect 493876 1164 493928 1216
rect 464252 1096 464304 1148
rect 469220 1096 469272 1148
rect 466460 1028 466512 1080
rect 471888 960 471940 1012
rect 464252 756 464304 808
rect 470600 824 470652 876
rect 475936 892 475988 944
rect 478880 1096 478932 1148
rect 488724 1096 488776 1148
rect 483572 960 483624 1012
rect 491116 1096 491168 1148
rect 499212 1232 499264 1284
rect 498292 1164 498344 1216
rect 510528 1164 510580 1216
rect 499120 1096 499172 1148
rect 505100 1096 505152 1148
rect 498200 1028 498252 1080
rect 499212 1028 499264 1080
rect 502340 1028 502392 1080
rect 500316 960 500368 1012
rect 472900 756 472952 808
rect 486148 824 486200 876
rect 478880 756 478932 808
rect 481548 756 481600 808
rect 483756 756 483808 808
rect 485964 756 486016 808
rect 499120 892 499172 944
rect 491116 688 491168 740
rect 509332 824 509384 876
rect 498292 756 498344 808
rect 514208 8 514260 60
<< metal2 >>
rect -1076 11960 -756 11972
rect -1076 11904 -1064 11960
rect -1008 11904 -984 11960
rect -928 11904 -904 11960
rect -848 11904 -824 11960
rect -768 11904 -756 11960
rect -1076 11880 -756 11904
rect -1076 11824 -1064 11880
rect -1008 11824 -984 11880
rect -928 11824 -904 11880
rect -848 11824 -824 11880
rect -768 11824 -756 11880
rect -1076 11800 -756 11824
rect -1076 11744 -1064 11800
rect -1008 11744 -984 11800
rect -928 11744 -904 11800
rect -848 11744 -824 11800
rect -768 11744 -756 11800
rect -1076 11720 -756 11744
rect -1076 11664 -1064 11720
rect -1008 11664 -984 11720
rect -928 11664 -904 11720
rect -848 11664 -824 11720
rect -768 11664 -756 11720
rect -1076 9648 -756 11664
rect -1076 9592 -1064 9648
rect -1008 9592 -984 9648
rect -928 9592 -904 9648
rect -848 9592 -824 9648
rect -768 9592 -756 9648
rect -1076 9568 -756 9592
rect -1076 9512 -1064 9568
rect -1008 9512 -984 9568
rect -928 9512 -904 9568
rect -848 9512 -824 9568
rect -768 9512 -756 9568
rect -1076 9488 -756 9512
rect -1076 9432 -1064 9488
rect -1008 9432 -984 9488
rect -928 9432 -904 9488
rect -848 9432 -824 9488
rect -768 9432 -756 9488
rect -1076 9408 -756 9432
rect -1076 9352 -1064 9408
rect -1008 9352 -984 9408
rect -928 9352 -904 9408
rect -848 9352 -824 9408
rect -768 9352 -756 9408
rect -1076 7744 -756 9352
rect -1076 7688 -1064 7744
rect -1008 7688 -984 7744
rect -928 7688 -904 7744
rect -848 7688 -824 7744
rect -768 7688 -756 7744
rect -1076 7664 -756 7688
rect -1076 7608 -1064 7664
rect -1008 7608 -984 7664
rect -928 7608 -904 7664
rect -848 7608 -824 7664
rect -768 7608 -756 7664
rect -1076 7584 -756 7608
rect -1076 7528 -1064 7584
rect -1008 7528 -984 7584
rect -928 7528 -904 7584
rect -848 7528 -824 7584
rect -768 7528 -756 7584
rect -1076 7504 -756 7528
rect -1076 7448 -1064 7504
rect -1008 7448 -984 7504
rect -928 7448 -904 7504
rect -848 7448 -824 7504
rect -768 7448 -756 7504
rect -1076 5840 -756 7448
rect -1076 5784 -1064 5840
rect -1008 5784 -984 5840
rect -928 5784 -904 5840
rect -848 5784 -824 5840
rect -768 5784 -756 5840
rect -1076 5760 -756 5784
rect -1076 5704 -1064 5760
rect -1008 5704 -984 5760
rect -928 5704 -904 5760
rect -848 5704 -824 5760
rect -768 5704 -756 5760
rect -1076 5680 -756 5704
rect -1076 5624 -1064 5680
rect -1008 5624 -984 5680
rect -928 5624 -904 5680
rect -848 5624 -824 5680
rect -768 5624 -756 5680
rect -1076 5600 -756 5624
rect -1076 5544 -1064 5600
rect -1008 5544 -984 5600
rect -928 5544 -904 5600
rect -848 5544 -824 5600
rect -768 5544 -756 5600
rect -1076 3936 -756 5544
rect -1076 3880 -1064 3936
rect -1008 3880 -984 3936
rect -928 3880 -904 3936
rect -848 3880 -824 3936
rect -768 3880 -756 3936
rect -1076 3856 -756 3880
rect -1076 3800 -1064 3856
rect -1008 3800 -984 3856
rect -928 3800 -904 3856
rect -848 3800 -824 3856
rect -768 3800 -756 3856
rect -1076 3776 -756 3800
rect -1076 3720 -1064 3776
rect -1008 3720 -984 3776
rect -928 3720 -904 3776
rect -848 3720 -824 3776
rect -768 3720 -756 3776
rect -1076 3696 -756 3720
rect -1076 3640 -1064 3696
rect -1008 3640 -984 3696
rect -928 3640 -904 3696
rect -848 3640 -824 3696
rect -768 3640 -756 3696
rect -1076 304 -756 3640
rect -416 11300 -96 11312
rect -416 11244 -404 11300
rect -348 11244 -324 11300
rect -268 11244 -244 11300
rect -188 11244 -164 11300
rect -108 11244 -96 11300
rect -416 11220 -96 11244
rect -416 11164 -404 11220
rect -348 11164 -324 11220
rect -268 11164 -244 11220
rect -188 11164 -164 11220
rect -108 11164 -96 11220
rect -416 11140 -96 11164
rect -416 11084 -404 11140
rect -348 11084 -324 11140
rect -268 11084 -244 11140
rect -188 11084 -164 11140
rect -108 11084 -96 11140
rect -416 11060 -96 11084
rect -416 11004 -404 11060
rect -348 11004 -324 11060
rect -268 11004 -244 11060
rect -188 11004 -164 11060
rect -108 11004 -96 11060
rect -416 8988 -96 11004
rect 66908 11300 67228 11972
rect 66908 11244 66920 11300
rect 66976 11244 67000 11300
rect 67056 11244 67080 11300
rect 67136 11244 67160 11300
rect 67216 11244 67228 11300
rect 66908 11220 67228 11244
rect 66908 11164 66920 11220
rect 66976 11164 67000 11220
rect 67056 11164 67080 11220
rect 67136 11164 67160 11220
rect 67216 11164 67228 11220
rect 66908 11140 67228 11164
rect 66908 11084 66920 11140
rect 66976 11084 67000 11140
rect 67056 11084 67080 11140
rect 67136 11084 67160 11140
rect 67216 11084 67228 11140
rect 66908 11060 67228 11084
rect 66908 11004 66920 11060
rect 66976 11004 67000 11060
rect 67056 11004 67080 11060
rect 67136 11004 67160 11060
rect 67216 11004 67228 11060
rect 56600 10328 56652 10334
rect 56600 10270 56652 10276
rect -416 8932 -404 8988
rect -348 8932 -324 8988
rect -268 8932 -244 8988
rect -188 8932 -164 8988
rect -108 8932 -96 8988
rect -416 8908 -96 8932
rect -416 8852 -404 8908
rect -348 8852 -324 8908
rect -268 8852 -244 8908
rect -188 8852 -164 8908
rect -108 8852 -96 8908
rect -416 8828 -96 8852
rect 43812 8900 43864 8906
rect 43812 8842 43864 8848
rect -416 8772 -404 8828
rect -348 8772 -324 8828
rect -268 8772 -244 8828
rect -188 8772 -164 8828
rect -108 8772 -96 8828
rect -416 8748 -96 8772
rect -416 8692 -404 8748
rect -348 8692 -324 8748
rect -268 8692 -244 8748
rect -188 8692 -164 8748
rect -108 8692 -96 8748
rect -416 7084 -96 8692
rect 36084 8424 36136 8430
rect 36084 8366 36136 8372
rect 33508 8356 33560 8362
rect 33508 8298 33560 8304
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect -416 7028 -404 7084
rect -348 7028 -324 7084
rect -268 7028 -244 7084
rect -188 7028 -164 7084
rect -108 7028 -96 7084
rect -416 7004 -96 7028
rect -416 6948 -404 7004
rect -348 6948 -324 7004
rect -268 6948 -244 7004
rect -188 6948 -164 7004
rect -108 6948 -96 7004
rect -416 6924 -96 6948
rect -416 6868 -404 6924
rect -348 6868 -324 6924
rect -268 6868 -244 6924
rect -188 6868 -164 6924
rect -108 6868 -96 6924
rect -416 6844 -96 6868
rect -416 6788 -404 6844
rect -348 6788 -324 6844
rect -268 6788 -244 6844
rect -188 6788 -164 6844
rect -108 6788 -96 6844
rect -416 5180 -96 6788
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect -416 5124 -404 5180
rect -348 5124 -324 5180
rect -268 5124 -244 5180
rect -188 5124 -164 5180
rect -108 5124 -96 5180
rect -416 5100 -96 5124
rect -416 5044 -404 5100
rect -348 5044 -324 5100
rect -268 5044 -244 5100
rect -188 5044 -164 5100
rect -108 5044 -96 5100
rect -416 5020 -96 5044
rect -416 4964 -404 5020
rect -348 4964 -324 5020
rect -268 4964 -244 5020
rect -188 4964 -164 5020
rect -108 4964 -96 5020
rect -416 4940 -96 4964
rect -416 4884 -404 4940
rect -348 4884 -324 4940
rect -268 4884 -244 4940
rect -188 4884 -164 4940
rect -108 4884 -96 4940
rect -416 3276 -96 4884
rect 1872 3738 1900 6122
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4448 3738 4476 3946
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect -416 3220 -404 3276
rect -348 3220 -324 3276
rect -268 3220 -244 3276
rect -188 3220 -164 3276
rect -108 3220 -96 3276
rect -416 3196 -96 3220
rect -416 3140 -404 3196
rect -348 3140 -324 3196
rect -268 3140 -244 3196
rect -188 3140 -164 3196
rect -108 3140 -96 3196
rect -416 3116 -96 3140
rect -416 3060 -404 3116
rect -348 3060 -324 3116
rect -268 3060 -244 3116
rect -188 3060 -164 3116
rect -108 3060 -96 3116
rect -416 3036 -96 3060
rect -416 2980 -404 3036
rect -348 2980 -324 3036
rect -268 2980 -244 3036
rect -188 2980 -164 3036
rect -108 2980 -96 3036
rect -416 964 -96 2980
rect 1320 2854 1348 3402
rect 3988 2854 4016 3402
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 848 2372 900 2378
rect 848 2314 900 2320
rect -416 908 -404 964
rect -348 908 -324 964
rect -268 908 -244 964
rect -188 908 -164 964
rect -108 908 -96 964
rect -416 884 -96 908
rect -416 828 -404 884
rect -348 828 -324 884
rect -268 828 -244 884
rect -188 828 -164 884
rect -108 828 -96 884
rect -416 804 -96 828
rect 860 814 888 2314
rect 1320 814 1348 2790
rect 3988 814 4016 2790
rect 5184 2650 5212 5170
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 3738 6868 5102
rect 9600 3738 9628 5238
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12176 3738 12204 4762
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5184 2446 5212 2586
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4172 882 4200 2246
rect 6012 882 6040 2314
rect 4160 876 4212 882
rect 4160 818 4212 824
rect 6000 876 6052 882
rect 6000 818 6052 824
rect 6196 814 6224 3334
rect 9140 2854 9168 3402
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 6564 2378 6592 2790
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 6748 814 6776 2382
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7024 1766 7052 2246
rect 7012 1760 7064 1766
rect 7012 1702 7064 1708
rect 8496 814 8524 2790
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9600 814 9628 2246
rect -416 748 -404 804
rect -348 748 -324 804
rect -268 748 -244 804
rect -188 748 -164 804
rect -108 748 -96 804
rect 848 808 900 814
rect 848 750 900 756
rect 1308 808 1360 814
rect 1308 750 1360 756
rect 3976 808 4028 814
rect 3976 750 4028 756
rect 6184 808 6236 814
rect 6184 750 6236 756
rect 6736 808 6788 814
rect 6736 750 6788 756
rect 8484 808 8536 814
rect 8484 750 8536 756
rect 9588 808 9640 814
rect 9588 750 9640 756
rect -416 724 -96 748
rect 10796 746 10824 2314
rect 11348 882 11376 3334
rect 12912 2582 12940 6190
rect 14752 3738 14780 7686
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17328 3738 17356 6258
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14292 2854 14320 3402
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 12900 2576 12952 2582
rect 12900 2518 12952 2524
rect 12912 2446 12940 2518
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 14292 1154 14320 2790
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14752 1834 14780 2246
rect 14740 1828 14792 1834
rect 14740 1770 14792 1776
rect 14280 1148 14332 1154
rect 14280 1090 14332 1096
rect 11336 876 11388 882
rect 11336 818 11388 824
rect 15948 814 15976 2314
rect 16592 950 16620 3334
rect 18064 2582 18092 5306
rect 19904 3738 19932 5714
rect 22480 3738 22508 7890
rect 29920 7540 29972 7546
rect 29920 7482 29972 7488
rect 29932 6322 29960 7482
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 19248 3460 19300 3466
rect 19248 3402 19300 3408
rect 19260 2854 19288 3402
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 18052 2576 18104 2582
rect 18052 2518 18104 2524
rect 18064 2446 18092 2518
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 1018 17356 2246
rect 19260 1358 19288 2790
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 19248 1352 19300 1358
rect 19248 1294 19300 1300
rect 20732 1290 20760 2246
rect 20720 1284 20772 1290
rect 20720 1226 20772 1232
rect 21652 1222 21680 3334
rect 23216 2378 23244 4558
rect 33152 3738 33180 6802
rect 33140 3732 33192 3738
rect 33140 3674 33192 3680
rect 31852 3664 31904 3670
rect 31852 3606 31904 3612
rect 29368 3528 29420 3534
rect 29368 3470 29420 3476
rect 24584 3460 24636 3466
rect 24584 3402 24636 3408
rect 28908 3460 28960 3466
rect 28908 3402 28960 3408
rect 24596 2854 24624 3402
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 27620 3392 27672 3398
rect 27620 3334 27672 3340
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 24584 2848 24636 2854
rect 24584 2790 24636 2796
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 21640 1216 21692 1222
rect 21640 1158 21692 1164
rect 23860 1086 23888 2790
rect 23940 2304 23992 2310
rect 23940 2246 23992 2252
rect 23952 1154 23980 2246
rect 24768 1284 24820 1290
rect 24768 1226 24820 1232
rect 23940 1148 23992 1154
rect 23940 1090 23992 1096
rect 23848 1080 23900 1086
rect 23848 1022 23900 1028
rect 17316 1012 17368 1018
rect 17316 954 17368 960
rect 16580 944 16632 950
rect 16580 886 16632 892
rect 24780 814 24808 1226
rect 24872 882 24900 3334
rect 27632 3058 27660 3334
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 28920 2854 28948 3402
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 28354 2408 28410 2417
rect 28354 2343 28356 2352
rect 28408 2343 28410 2352
rect 28356 2314 28408 2320
rect 25044 2304 25096 2310
rect 25044 2246 25096 2252
rect 27620 2304 27672 2310
rect 27620 2246 27672 2252
rect 28264 2304 28316 2310
rect 28264 2246 28316 2252
rect 25056 1698 25084 2246
rect 25044 1692 25096 1698
rect 25044 1634 25096 1640
rect 27632 1222 27660 2246
rect 28276 1290 28304 2246
rect 28264 1284 28316 1290
rect 28264 1226 28316 1232
rect 28920 1222 28948 2790
rect 29092 1352 29144 1358
rect 29092 1294 29144 1300
rect 27620 1216 27672 1222
rect 27620 1158 27672 1164
rect 28908 1216 28960 1222
rect 28908 1158 28960 1164
rect 24860 876 24912 882
rect 24860 818 24912 824
rect 29104 814 29132 1294
rect 29380 950 29408 3470
rect 30196 2304 30248 2310
rect 30196 2246 30248 2252
rect 30208 2038 30236 2246
rect 30196 2032 30248 2038
rect 30196 1974 30248 1980
rect 31864 1018 31892 3606
rect 32770 3496 32826 3505
rect 32770 3431 32826 3440
rect 33140 3460 33192 3466
rect 32784 3398 32812 3431
rect 33140 3402 33192 3408
rect 32772 3392 32824 3398
rect 32772 3334 32824 3340
rect 32772 2304 32824 2310
rect 32772 2246 32824 2252
rect 32784 1154 32812 2246
rect 32772 1148 32824 1154
rect 32772 1090 32824 1096
rect 31852 1012 31904 1018
rect 31852 954 31904 960
rect 33152 950 33180 3402
rect 33520 2514 33548 8298
rect 35900 8084 35952 8090
rect 35900 8026 35952 8032
rect 35912 3602 35940 8026
rect 36096 3738 36124 8366
rect 42984 7812 43036 7818
rect 42984 7754 43036 7760
rect 40408 6452 40460 6458
rect 40408 6394 40460 6400
rect 36084 3732 36136 3738
rect 36084 3674 36136 3680
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 36096 3534 36124 3674
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 39120 3392 39172 3398
rect 39120 3334 39172 3340
rect 36820 2916 36872 2922
rect 36820 2858 36872 2864
rect 34888 2848 34940 2854
rect 34888 2790 34940 2796
rect 33508 2508 33560 2514
rect 33508 2450 33560 2456
rect 34900 2378 34928 2790
rect 34888 2372 34940 2378
rect 34888 2314 34940 2320
rect 34900 2122 34928 2314
rect 35348 2304 35400 2310
rect 35348 2246 35400 2252
rect 34808 2094 34928 2122
rect 33508 1352 33560 1358
rect 33508 1294 33560 1300
rect 29368 944 29420 950
rect 29368 886 29420 892
rect 33140 944 33192 950
rect 33140 886 33192 892
rect 15936 808 15988 814
rect 15936 750 15988 756
rect 24768 808 24820 814
rect 24768 750 24820 756
rect 29092 808 29144 814
rect 29092 750 29144 756
rect 33520 746 33548 1294
rect 34808 1290 34836 2094
rect 35360 1970 35388 2246
rect 35348 1964 35400 1970
rect 35348 1906 35400 1912
rect 34796 1284 34848 1290
rect 34796 1226 34848 1232
rect 35716 1284 35768 1290
rect 35716 1226 35768 1232
rect 35728 814 35756 1226
rect 36832 950 36860 2858
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 37476 2378 37504 2790
rect 37464 2372 37516 2378
rect 37464 2314 37516 2320
rect 37476 1086 37504 2314
rect 37924 2304 37976 2310
rect 37924 2246 37976 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 37936 2106 37964 2246
rect 37924 2100 37976 2106
rect 37924 2042 37976 2048
rect 38672 1358 38700 2246
rect 38660 1352 38712 1358
rect 38660 1294 38712 1300
rect 37832 1148 37884 1154
rect 37832 1090 37884 1096
rect 37464 1080 37516 1086
rect 37464 1022 37516 1028
rect 36820 944 36872 950
rect 36820 886 36872 892
rect 37844 814 37872 1090
rect 39132 1086 39160 3334
rect 40420 2446 40448 6394
rect 42996 6254 43024 7754
rect 42984 6248 43036 6254
rect 42984 6190 43036 6196
rect 42892 6112 42944 6118
rect 42892 6054 42944 6060
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 40696 2922 40724 3470
rect 40684 2916 40736 2922
rect 40684 2858 40736 2864
rect 41328 2916 41380 2922
rect 41328 2858 41380 2864
rect 41234 2544 41290 2553
rect 41234 2479 41236 2488
rect 41288 2479 41290 2488
rect 41236 2450 41288 2456
rect 40408 2440 40460 2446
rect 40408 2382 40460 2388
rect 39120 1080 39172 1086
rect 39120 1022 39172 1028
rect 40868 1080 40920 1086
rect 40868 1022 40920 1028
rect 40880 814 40908 1022
rect 41340 1018 41368 2858
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 42812 2446 42840 2790
rect 42904 2582 42932 6054
rect 43824 3738 43852 8842
rect 46940 6996 46992 7002
rect 46940 6938 46992 6944
rect 46952 6186 46980 6938
rect 46940 6180 46992 6186
rect 46940 6122 46992 6128
rect 48780 5908 48832 5914
rect 48780 5850 48832 5856
rect 47400 5636 47452 5642
rect 47400 5578 47452 5584
rect 45652 5024 45704 5030
rect 45652 4966 45704 4972
rect 45664 3738 45692 4966
rect 43812 3732 43864 3738
rect 43812 3674 43864 3680
rect 45652 3732 45704 3738
rect 45652 3674 45704 3680
rect 43824 3534 43852 3674
rect 47412 3602 47440 5578
rect 48228 4072 48280 4078
rect 48228 4014 48280 4020
rect 48240 3738 48268 4014
rect 48228 3732 48280 3738
rect 48228 3674 48280 3680
rect 47400 3596 47452 3602
rect 47400 3538 47452 3544
rect 43812 3528 43864 3534
rect 43812 3470 43864 3476
rect 45836 3528 45888 3534
rect 45836 3470 45888 3476
rect 43168 3392 43220 3398
rect 43168 3334 43220 3340
rect 42892 2576 42944 2582
rect 42892 2518 42944 2524
rect 42800 2440 42852 2446
rect 42800 2382 42852 2388
rect 42812 1426 42840 2382
rect 42800 1420 42852 1426
rect 42800 1362 42852 1368
rect 42156 1352 42208 1358
rect 42156 1294 42208 1300
rect 41328 1012 41380 1018
rect 41328 954 41380 960
rect 42168 814 42196 1294
rect 43180 1086 43208 3334
rect 45848 2922 45876 3470
rect 45836 2916 45888 2922
rect 45836 2858 45888 2864
rect 44088 2304 44140 2310
rect 44088 2246 44140 2252
rect 46020 2304 46072 2310
rect 46020 2246 46072 2252
rect 43260 1284 43312 1290
rect 43260 1226 43312 1232
rect 43168 1080 43220 1086
rect 43168 1022 43220 1028
rect 43272 814 43300 1226
rect 44100 1154 44128 2246
rect 44088 1148 44140 1154
rect 44088 1090 44140 1096
rect 46032 1018 46060 2246
rect 48792 2038 48820 5850
rect 56508 5568 56560 5574
rect 56508 5510 56560 5516
rect 55128 3528 55180 3534
rect 55128 3470 55180 3476
rect 49700 3392 49752 3398
rect 49700 3334 49752 3340
rect 51540 3392 51592 3398
rect 51540 3334 51592 3340
rect 52736 3392 52788 3398
rect 52736 3334 52788 3340
rect 48962 2680 49018 2689
rect 48962 2615 49018 2624
rect 48976 2446 49004 2615
rect 48964 2440 49016 2446
rect 48964 2382 49016 2388
rect 48780 2032 48832 2038
rect 48780 1974 48832 1980
rect 49712 1426 49740 3334
rect 51552 2990 51580 3334
rect 51540 2984 51592 2990
rect 51540 2926 51592 2932
rect 50528 2848 50580 2854
rect 50528 2790 50580 2796
rect 50540 2446 50568 2790
rect 50528 2440 50580 2446
rect 50528 2382 50580 2388
rect 50540 1494 50568 2382
rect 52644 2372 52696 2378
rect 52644 2314 52696 2320
rect 50804 2304 50856 2310
rect 50804 2246 50856 2252
rect 50816 1630 50844 2246
rect 50804 1624 50856 1630
rect 50804 1566 50856 1572
rect 50528 1488 50580 1494
rect 50528 1430 50580 1436
rect 51908 1488 51960 1494
rect 51908 1430 51960 1436
rect 49700 1420 49752 1426
rect 49700 1362 49752 1368
rect 49056 1352 49108 1358
rect 48976 1312 49056 1340
rect 48976 1154 49004 1312
rect 49056 1294 49108 1300
rect 49792 1284 49844 1290
rect 49792 1226 49844 1232
rect 47676 1148 47728 1154
rect 47676 1090 47728 1096
rect 48964 1148 49016 1154
rect 48964 1090 49016 1096
rect 49056 1148 49108 1154
rect 49056 1090 49108 1096
rect 46020 1012 46072 1018
rect 46020 954 46072 960
rect 47688 814 47716 1090
rect 47860 1080 47912 1086
rect 47912 1028 48084 1034
rect 47860 1022 48084 1028
rect 47872 1018 48084 1022
rect 47872 1012 48096 1018
rect 47872 1006 48044 1012
rect 48044 954 48096 960
rect 49068 898 49096 1090
rect 48884 882 49096 898
rect 48872 876 49096 882
rect 48924 870 49096 876
rect 48872 818 48924 824
rect 49804 814 49832 1226
rect 51920 882 51948 1430
rect 52656 950 52684 2314
rect 52748 1018 52776 3334
rect 55140 2854 55168 3470
rect 55956 3392 56008 3398
rect 55956 3334 56008 3340
rect 53104 2848 53156 2854
rect 53104 2790 53156 2796
rect 53840 2848 53892 2854
rect 53840 2790 53892 2796
rect 55128 2848 55180 2854
rect 55968 2825 55996 3334
rect 55128 2790 55180 2796
rect 55954 2816 56010 2825
rect 53116 2446 53144 2790
rect 53104 2440 53156 2446
rect 53104 2382 53156 2388
rect 53564 2440 53616 2446
rect 53564 2382 53616 2388
rect 53380 2304 53432 2310
rect 53380 2246 53432 2252
rect 53392 2038 53420 2246
rect 53380 2032 53432 2038
rect 53380 1974 53432 1980
rect 53576 1222 53604 2382
rect 53852 1426 53880 2790
rect 55954 2751 56010 2760
rect 56520 1970 56548 5510
rect 56612 2446 56640 10270
rect 66908 9274 67228 11004
rect 66908 9222 66914 9274
rect 66966 9222 66978 9274
rect 67030 9222 67042 9274
rect 67094 9222 67106 9274
rect 67158 9222 67170 9274
rect 67222 9222 67228 9274
rect 66908 8988 67228 9222
rect 66908 8932 66920 8988
rect 66976 8932 67000 8988
rect 67056 8932 67080 8988
rect 67136 8932 67160 8988
rect 67216 8932 67228 8988
rect 66908 8908 67228 8932
rect 66908 8852 66920 8908
rect 66976 8852 67000 8908
rect 67056 8852 67080 8908
rect 67136 8852 67160 8908
rect 67216 8852 67228 8908
rect 66908 8828 67228 8852
rect 66908 8772 66920 8828
rect 66976 8772 67000 8828
rect 67056 8772 67080 8828
rect 67136 8772 67160 8828
rect 67216 8772 67228 8828
rect 66908 8748 67228 8772
rect 66908 8692 66920 8748
rect 66976 8692 67000 8748
rect 67056 8692 67080 8748
rect 67136 8692 67160 8748
rect 67216 8692 67228 8748
rect 66908 8186 67228 8692
rect 67568 11960 67888 11972
rect 67568 11904 67580 11960
rect 67636 11904 67660 11960
rect 67716 11904 67740 11960
rect 67796 11904 67820 11960
rect 67876 11904 67888 11960
rect 67568 11880 67888 11904
rect 92204 11960 92256 11966
rect 92204 11902 92256 11908
rect 67568 11824 67580 11880
rect 67636 11824 67660 11880
rect 67716 11824 67740 11880
rect 67796 11824 67820 11880
rect 67876 11824 67888 11880
rect 67568 11800 67888 11824
rect 67568 11744 67580 11800
rect 67636 11744 67660 11800
rect 67716 11744 67740 11800
rect 67796 11744 67820 11800
rect 67876 11744 67888 11800
rect 67568 11720 67888 11744
rect 67568 11664 67580 11720
rect 67636 11664 67660 11720
rect 67716 11664 67740 11720
rect 67796 11664 67820 11720
rect 67876 11664 67888 11720
rect 67568 9818 67888 11664
rect 92112 9988 92164 9994
rect 92112 9930 92164 9936
rect 67568 9766 67574 9818
rect 67626 9766 67638 9818
rect 67690 9766 67702 9818
rect 67754 9766 67766 9818
rect 67818 9766 67830 9818
rect 67882 9766 67888 9818
rect 67568 9648 67888 9766
rect 67568 9592 67580 9648
rect 67636 9592 67660 9648
rect 67716 9592 67740 9648
rect 67796 9592 67820 9648
rect 67876 9592 67888 9648
rect 67568 9568 67888 9592
rect 67568 9512 67580 9568
rect 67636 9512 67660 9568
rect 67716 9512 67740 9568
rect 67796 9512 67820 9568
rect 67876 9512 67888 9568
rect 67568 9488 67888 9512
rect 67568 9432 67580 9488
rect 67636 9432 67660 9488
rect 67716 9432 67740 9488
rect 67796 9432 67820 9488
rect 67876 9432 67888 9488
rect 82452 9512 82504 9518
rect 82452 9454 82504 9460
rect 67568 9408 67888 9432
rect 67568 9352 67580 9408
rect 67636 9352 67660 9408
rect 67716 9352 67740 9408
rect 67796 9352 67820 9408
rect 67876 9352 67888 9408
rect 74724 9444 74776 9450
rect 74724 9386 74776 9392
rect 67568 8730 67888 9352
rect 67568 8678 67574 8730
rect 67626 8678 67638 8730
rect 67690 8678 67702 8730
rect 67754 8678 67766 8730
rect 67818 8678 67830 8730
rect 67882 8678 67888 8730
rect 67270 8528 67326 8537
rect 67270 8463 67326 8472
rect 66908 8134 66914 8186
rect 66966 8134 66978 8186
rect 67030 8134 67042 8186
rect 67094 8134 67106 8186
rect 67158 8134 67170 8186
rect 67222 8134 67228 8186
rect 59268 8016 59320 8022
rect 59268 7958 59320 7964
rect 59176 4752 59228 4758
rect 59176 4694 59228 4700
rect 56692 3392 56744 3398
rect 56692 3334 56744 3340
rect 56600 2440 56652 2446
rect 56600 2382 56652 2388
rect 56508 1964 56560 1970
rect 56508 1906 56560 1912
rect 53840 1420 53892 1426
rect 53840 1362 53892 1368
rect 56140 1352 56192 1358
rect 56140 1294 56192 1300
rect 53748 1284 53800 1290
rect 53748 1226 53800 1232
rect 53564 1216 53616 1222
rect 53564 1158 53616 1164
rect 53760 1170 53788 1226
rect 53760 1154 54064 1170
rect 53760 1148 54076 1154
rect 53760 1142 54024 1148
rect 54024 1090 54076 1096
rect 52736 1012 52788 1018
rect 52736 954 52788 960
rect 56152 950 56180 1294
rect 56232 1284 56284 1290
rect 56232 1226 56284 1232
rect 52644 944 52696 950
rect 52644 886 52696 892
rect 56140 944 56192 950
rect 56140 886 56192 892
rect 56244 882 56272 1226
rect 56704 1154 56732 3334
rect 58256 2848 58308 2854
rect 58256 2790 58308 2796
rect 58268 2446 58296 2790
rect 59188 2650 59216 4694
rect 59280 3738 59308 7958
rect 63500 7472 63552 7478
rect 63500 7414 63552 7420
rect 62120 6384 62172 6390
rect 62120 6326 62172 6332
rect 62132 3738 62160 6326
rect 63512 4826 63540 7414
rect 66908 7098 67228 8134
rect 66908 7046 66914 7098
rect 66966 7084 66978 7098
rect 67030 7084 67042 7098
rect 67094 7084 67106 7098
rect 67158 7084 67170 7098
rect 66976 7046 66978 7084
rect 67158 7046 67160 7084
rect 67222 7046 67228 7098
rect 66908 7028 66920 7046
rect 66976 7028 67000 7046
rect 67056 7028 67080 7046
rect 67136 7028 67160 7046
rect 67216 7028 67228 7046
rect 66908 7004 67228 7028
rect 66908 6948 66920 7004
rect 66976 6948 67000 7004
rect 67056 6948 67080 7004
rect 67136 6948 67160 7004
rect 67216 6948 67228 7004
rect 66908 6924 67228 6948
rect 66908 6868 66920 6924
rect 66976 6868 67000 6924
rect 67056 6868 67080 6924
rect 67136 6868 67160 6924
rect 67216 6868 67228 6924
rect 66908 6844 67228 6868
rect 66908 6788 66920 6844
rect 66976 6788 67000 6844
rect 67056 6788 67080 6844
rect 67136 6788 67160 6844
rect 67216 6788 67228 6844
rect 66908 6010 67228 6788
rect 66908 5958 66914 6010
rect 66966 5958 66978 6010
rect 67030 5958 67042 6010
rect 67094 5958 67106 6010
rect 67158 5958 67170 6010
rect 67222 5958 67228 6010
rect 66908 5180 67228 5958
rect 66908 5124 66920 5180
rect 66976 5124 67000 5180
rect 67056 5124 67080 5180
rect 67136 5124 67160 5180
rect 67216 5124 67228 5180
rect 66908 5100 67228 5124
rect 66908 5044 66920 5100
rect 66976 5044 67000 5100
rect 67056 5044 67080 5100
rect 67136 5044 67160 5100
rect 67216 5044 67228 5100
rect 66908 5020 67228 5044
rect 66908 4964 66920 5020
rect 66976 4964 67000 5020
rect 67056 4964 67080 5020
rect 67136 4964 67160 5020
rect 67216 4964 67228 5020
rect 66908 4940 67228 4964
rect 66908 4922 66920 4940
rect 66976 4922 67000 4940
rect 67056 4922 67080 4940
rect 67136 4922 67160 4940
rect 67216 4922 67228 4940
rect 66908 4870 66914 4922
rect 66976 4884 66978 4922
rect 67158 4884 67160 4922
rect 66966 4870 66978 4884
rect 67030 4870 67042 4884
rect 67094 4870 67106 4884
rect 67158 4870 67170 4884
rect 67222 4870 67228 4922
rect 63500 4820 63552 4826
rect 63500 4762 63552 4768
rect 66908 3834 67228 4870
rect 66908 3782 66914 3834
rect 66966 3782 66978 3834
rect 67030 3782 67042 3834
rect 67094 3782 67106 3834
rect 67158 3782 67170 3834
rect 67222 3782 67228 3834
rect 59268 3732 59320 3738
rect 59268 3674 59320 3680
rect 62120 3732 62172 3738
rect 62120 3674 62172 3680
rect 63500 3732 63552 3738
rect 63500 3674 63552 3680
rect 59280 3534 59308 3674
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 60660 2854 60688 3470
rect 62960 3466 63172 3482
rect 62948 3460 63184 3466
rect 63000 3454 63132 3460
rect 62948 3402 63000 3408
rect 63132 3402 63184 3408
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 59360 2848 59412 2854
rect 59360 2790 59412 2796
rect 60648 2848 60700 2854
rect 60648 2790 60700 2796
rect 59176 2644 59228 2650
rect 59176 2586 59228 2592
rect 57980 2440 58032 2446
rect 57980 2382 58032 2388
rect 58256 2440 58308 2446
rect 58256 2382 58308 2388
rect 57888 2372 57940 2378
rect 57888 2314 57940 2320
rect 57900 1494 57928 2314
rect 57888 1488 57940 1494
rect 57888 1430 57940 1436
rect 57992 1222 58020 2382
rect 58532 2304 58584 2310
rect 58532 2246 58584 2252
rect 58544 1970 58572 2246
rect 58532 1964 58584 1970
rect 58532 1906 58584 1912
rect 58992 1284 59044 1290
rect 58992 1226 59044 1232
rect 57980 1216 58032 1222
rect 57980 1158 58032 1164
rect 58532 1216 58584 1222
rect 58532 1158 58584 1164
rect 56692 1148 56744 1154
rect 56692 1090 56744 1096
rect 57428 1148 57480 1154
rect 57428 1090 57480 1096
rect 51908 876 51960 882
rect 51908 818 51960 824
rect 56232 876 56284 882
rect 56232 818 56284 824
rect 35716 808 35768 814
rect 35716 750 35768 756
rect 37832 808 37884 814
rect 37832 750 37884 756
rect 40868 808 40920 814
rect 40868 750 40920 756
rect 42156 808 42208 814
rect 42156 750 42208 756
rect 43260 808 43312 814
rect 43260 750 43312 756
rect 47676 808 47728 814
rect 47676 750 47728 756
rect 49792 808 49844 814
rect 49792 750 49844 756
rect 57440 746 57468 1090
rect 58544 814 58572 1158
rect 59004 882 59032 1226
rect 59372 1086 59400 2790
rect 60752 1442 60780 3334
rect 61108 3188 61160 3194
rect 61108 3130 61160 3136
rect 61120 2650 61148 3130
rect 61108 2644 61160 2650
rect 61108 2586 61160 2592
rect 60556 1420 60608 1426
rect 60556 1362 60608 1368
rect 60660 1414 60780 1442
rect 62764 1488 62816 1494
rect 62764 1430 62816 1436
rect 59636 1284 59688 1290
rect 59636 1226 59688 1232
rect 59360 1080 59412 1086
rect 59360 1022 59412 1028
rect 58992 876 59044 882
rect 58992 818 59044 824
rect 58532 808 58584 814
rect 58532 750 58584 756
rect 59648 746 59676 1226
rect 60568 1018 60596 1362
rect 60660 1358 60688 1414
rect 60648 1352 60700 1358
rect 60648 1294 60700 1300
rect 60740 1352 60792 1358
rect 60740 1294 60792 1300
rect 60556 1012 60608 1018
rect 60556 954 60608 960
rect 60752 814 60780 1294
rect 62776 1222 62804 1430
rect 63224 1284 63276 1290
rect 63224 1226 63276 1232
rect 62764 1216 62816 1222
rect 62764 1158 62816 1164
rect 61844 1080 61896 1086
rect 61844 1022 61896 1028
rect 61856 814 61884 1022
rect 63236 1018 63264 1226
rect 63224 1012 63276 1018
rect 63224 954 63276 960
rect 63512 950 63540 3674
rect 64880 3392 64932 3398
rect 64880 3334 64932 3340
rect 63684 2304 63736 2310
rect 63684 2246 63736 2252
rect 64420 2304 64472 2310
rect 64420 2246 64472 2252
rect 63696 1562 63724 2246
rect 64432 2145 64460 2246
rect 64418 2136 64474 2145
rect 64418 2071 64474 2080
rect 63684 1556 63736 1562
rect 63684 1498 63736 1504
rect 64892 1494 64920 3334
rect 66908 3276 67228 3782
rect 67284 3738 67312 8463
rect 67568 7744 67888 8678
rect 71044 7880 71096 7886
rect 71044 7822 71096 7828
rect 67568 7688 67580 7744
rect 67636 7688 67660 7744
rect 67716 7688 67740 7744
rect 67796 7688 67820 7744
rect 67876 7688 67888 7744
rect 67568 7664 67888 7688
rect 67568 7642 67580 7664
rect 67636 7642 67660 7664
rect 67716 7642 67740 7664
rect 67796 7642 67820 7664
rect 67876 7642 67888 7664
rect 67568 7590 67574 7642
rect 67636 7608 67638 7642
rect 67818 7608 67820 7642
rect 67626 7590 67638 7608
rect 67690 7590 67702 7608
rect 67754 7590 67766 7608
rect 67818 7590 67830 7608
rect 67882 7590 67888 7642
rect 67568 7584 67888 7590
rect 67568 7528 67580 7584
rect 67636 7528 67660 7584
rect 67716 7528 67740 7584
rect 67796 7528 67820 7584
rect 67876 7528 67888 7584
rect 67568 7504 67888 7528
rect 67568 7448 67580 7504
rect 67636 7448 67660 7504
rect 67716 7448 67740 7504
rect 67796 7448 67820 7504
rect 67876 7448 67888 7504
rect 67568 6554 67888 7448
rect 67568 6502 67574 6554
rect 67626 6502 67638 6554
rect 67690 6502 67702 6554
rect 67754 6502 67766 6554
rect 67818 6502 67830 6554
rect 67882 6502 67888 6554
rect 67568 5840 67888 6502
rect 68928 6180 68980 6186
rect 68928 6122 68980 6128
rect 67568 5784 67580 5840
rect 67636 5784 67660 5840
rect 67716 5784 67740 5840
rect 67796 5784 67820 5840
rect 67876 5784 67888 5840
rect 67568 5760 67888 5784
rect 67568 5704 67580 5760
rect 67636 5704 67660 5760
rect 67716 5704 67740 5760
rect 67796 5704 67820 5760
rect 67876 5704 67888 5760
rect 67568 5680 67888 5704
rect 67568 5624 67580 5680
rect 67636 5624 67660 5680
rect 67716 5624 67740 5680
rect 67796 5624 67820 5680
rect 67876 5624 67888 5680
rect 67568 5600 67888 5624
rect 67568 5544 67580 5600
rect 67636 5544 67660 5600
rect 67716 5544 67740 5600
rect 67796 5544 67820 5600
rect 67876 5544 67888 5600
rect 67568 5466 67888 5544
rect 67568 5414 67574 5466
rect 67626 5414 67638 5466
rect 67690 5414 67702 5466
rect 67754 5414 67766 5466
rect 67818 5414 67830 5466
rect 67882 5414 67888 5466
rect 67568 4378 67888 5414
rect 68836 5092 68888 5098
rect 68836 5034 68888 5040
rect 67568 4326 67574 4378
rect 67626 4326 67638 4378
rect 67690 4326 67702 4378
rect 67754 4326 67766 4378
rect 67818 4326 67830 4378
rect 67882 4326 67888 4378
rect 67568 3936 67888 4326
rect 67568 3880 67580 3936
rect 67636 3880 67660 3936
rect 67716 3880 67740 3936
rect 67796 3880 67820 3936
rect 67876 3880 67888 3936
rect 67568 3856 67888 3880
rect 67568 3800 67580 3856
rect 67636 3800 67660 3856
rect 67716 3800 67740 3856
rect 67796 3800 67820 3856
rect 67876 3800 67888 3856
rect 67568 3776 67888 3800
rect 67272 3732 67324 3738
rect 67272 3674 67324 3680
rect 67568 3720 67580 3776
rect 67636 3720 67660 3776
rect 67716 3720 67740 3776
rect 67796 3720 67820 3776
rect 67876 3720 67888 3776
rect 67568 3696 67888 3720
rect 67284 3534 67312 3674
rect 67568 3640 67580 3696
rect 67636 3640 67660 3696
rect 67716 3640 67740 3696
rect 67796 3640 67820 3696
rect 67876 3640 67888 3696
rect 67272 3528 67324 3534
rect 67272 3470 67324 3476
rect 66908 3220 66920 3276
rect 66976 3220 67000 3276
rect 67056 3220 67080 3276
rect 67136 3220 67160 3276
rect 67216 3220 67228 3276
rect 66908 3196 67228 3220
rect 66908 3140 66920 3196
rect 66976 3140 67000 3196
rect 67056 3140 67080 3196
rect 67136 3140 67160 3196
rect 67216 3140 67228 3196
rect 66908 3116 67228 3140
rect 66908 3060 66920 3116
rect 66976 3060 67000 3116
rect 67056 3060 67080 3116
rect 67136 3060 67160 3116
rect 67216 3060 67228 3116
rect 66908 3036 67228 3060
rect 66908 2980 66920 3036
rect 66976 2980 67000 3036
rect 67056 2980 67080 3036
rect 67136 2980 67160 3036
rect 67216 2980 67228 3036
rect 65248 2848 65300 2854
rect 65248 2790 65300 2796
rect 65260 2446 65288 2790
rect 66908 2746 67228 2980
rect 66908 2694 66914 2746
rect 66966 2694 66978 2746
rect 67030 2694 67042 2746
rect 67094 2694 67106 2746
rect 67158 2694 67170 2746
rect 67222 2694 67228 2746
rect 65248 2440 65300 2446
rect 65248 2382 65300 2388
rect 64880 1488 64932 1494
rect 64880 1430 64932 1436
rect 63592 1216 63644 1222
rect 63592 1158 63644 1164
rect 63500 944 63552 950
rect 63500 886 63552 892
rect 60740 808 60792 814
rect 60740 750 60792 756
rect 61844 808 61896 814
rect 63604 762 63632 1158
rect 63960 1148 64012 1154
rect 63960 1090 64012 1096
rect 63972 814 64000 1090
rect 65064 1012 65116 1018
rect 65064 954 65116 960
rect 65076 814 65104 954
rect 65260 882 65288 2382
rect 66260 2304 66312 2310
rect 66260 2246 66312 2252
rect 66272 1494 66300 2246
rect 66720 1896 66772 1902
rect 66720 1838 66772 1844
rect 66260 1488 66312 1494
rect 66260 1430 66312 1436
rect 66168 1352 66220 1358
rect 66168 1294 66220 1300
rect 65248 876 65300 882
rect 65248 818 65300 824
rect 66180 814 66208 1294
rect 66732 1222 66760 1838
rect 66720 1216 66772 1222
rect 66720 1158 66772 1164
rect 66812 1216 66864 1222
rect 66812 1158 66864 1164
rect 66824 814 66852 1158
rect 66908 964 67228 2694
rect 66908 908 66920 964
rect 66976 908 67000 964
rect 67056 908 67080 964
rect 67136 908 67160 964
rect 67216 908 67228 964
rect 66908 884 67228 908
rect 66908 828 66920 884
rect 66976 828 67000 884
rect 67056 828 67080 884
rect 67136 828 67160 884
rect 67216 828 67228 884
rect 61844 750 61896 756
rect 62868 746 63632 762
rect 63960 808 64012 814
rect 63960 750 64012 756
rect 65064 808 65116 814
rect 65064 750 65116 756
rect 66168 808 66220 814
rect 66168 750 66220 756
rect 66812 808 66864 814
rect 66812 750 66864 756
rect 66908 804 67228 828
rect -416 668 -404 724
rect -348 668 -324 724
rect -268 668 -244 724
rect -188 668 -164 724
rect -108 668 -96 724
rect 10784 740 10836 746
rect 10784 682 10836 688
rect 33508 740 33560 746
rect 33508 682 33560 688
rect 57428 740 57480 746
rect 57428 682 57480 688
rect 59636 740 59688 746
rect 59636 682 59688 688
rect 62856 740 63632 746
rect 62908 734 63632 740
rect 66908 748 66920 804
rect 66976 748 67000 804
rect 67056 748 67080 804
rect 67136 748 67160 804
rect 67216 748 67228 804
rect 62856 682 62908 688
rect 66908 724 67228 748
rect -416 656 -96 668
rect 66908 668 66920 724
rect 66976 668 67000 724
rect 67056 668 67080 724
rect 67136 668 67160 724
rect 67216 668 67228 724
rect -1076 248 -1064 304
rect -1008 248 -984 304
rect -928 248 -904 304
rect -848 248 -824 304
rect -768 248 -756 304
rect -1076 224 -756 248
rect -1076 168 -1064 224
rect -1008 168 -984 224
rect -928 168 -904 224
rect -848 168 -824 224
rect -768 168 -756 224
rect -1076 144 -756 168
rect -1076 88 -1064 144
rect -1008 88 -984 144
rect -928 88 -904 144
rect -848 88 -824 144
rect -768 88 -756 144
rect -1076 64 -756 88
rect -1076 8 -1064 64
rect -1008 8 -984 64
rect -928 8 -904 64
rect -848 8 -824 64
rect -768 8 -756 64
rect -1076 -4 -756 8
rect 66908 -4 67228 668
rect 67568 3290 67888 3640
rect 67568 3238 67574 3290
rect 67626 3238 67638 3290
rect 67690 3238 67702 3290
rect 67754 3238 67766 3290
rect 67818 3238 67830 3290
rect 67882 3238 67888 3290
rect 67568 2202 67888 3238
rect 67916 2916 67968 2922
rect 67916 2858 67968 2864
rect 67568 2150 67574 2202
rect 67626 2150 67638 2202
rect 67690 2150 67702 2202
rect 67754 2150 67766 2202
rect 67818 2150 67830 2202
rect 67882 2150 67888 2202
rect 67568 304 67888 2150
rect 67928 1426 67956 2858
rect 68560 2848 68612 2854
rect 68560 2790 68612 2796
rect 68572 2446 68600 2790
rect 68848 2650 68876 5034
rect 68940 5030 68968 6122
rect 68928 5024 68980 5030
rect 68928 4966 68980 4972
rect 71056 4010 71084 7822
rect 73988 4820 74040 4826
rect 73988 4762 74040 4768
rect 71044 4004 71096 4010
rect 71044 3946 71096 3952
rect 71412 3936 71464 3942
rect 71412 3878 71464 3884
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 71228 3528 71280 3534
rect 71228 3470 71280 3476
rect 69032 3398 69060 3470
rect 69020 3392 69072 3398
rect 69020 3334 69072 3340
rect 71240 3126 71268 3470
rect 71424 3398 71452 3878
rect 71412 3392 71464 3398
rect 71412 3334 71464 3340
rect 71504 3392 71556 3398
rect 71504 3334 71556 3340
rect 71228 3120 71280 3126
rect 71228 3062 71280 3068
rect 71240 2922 71268 3062
rect 71228 2916 71280 2922
rect 71228 2858 71280 2864
rect 71516 2854 71544 3334
rect 71780 2916 71832 2922
rect 71780 2858 71832 2864
rect 70400 2848 70452 2854
rect 70400 2790 70452 2796
rect 71504 2848 71556 2854
rect 71504 2790 71556 2796
rect 68836 2644 68888 2650
rect 68836 2586 68888 2592
rect 68560 2440 68612 2446
rect 68560 2382 68612 2388
rect 67916 1420 67968 1426
rect 67916 1362 67968 1368
rect 68572 1290 68600 2382
rect 70412 1902 70440 2790
rect 71412 2304 71464 2310
rect 71412 2246 71464 2252
rect 70400 1896 70452 1902
rect 70400 1838 70452 1844
rect 69480 1556 69532 1562
rect 69480 1498 69532 1504
rect 68560 1284 68612 1290
rect 68560 1226 68612 1232
rect 69492 1222 69520 1498
rect 69480 1216 69532 1222
rect 68098 1184 68154 1193
rect 69480 1158 69532 1164
rect 69664 1216 69716 1222
rect 69664 1158 69716 1164
rect 69846 1184 69902 1193
rect 68098 1119 68154 1128
rect 68112 1018 68140 1119
rect 68284 1080 68336 1086
rect 68284 1022 68336 1028
rect 68100 1012 68152 1018
rect 68100 954 68152 960
rect 68296 814 68324 1022
rect 68468 1012 68520 1018
rect 68468 954 68520 960
rect 68480 898 68508 954
rect 68480 882 68784 898
rect 68480 876 68796 882
rect 68480 870 68744 876
rect 68744 818 68796 824
rect 68284 808 68336 814
rect 69676 762 69704 1158
rect 69846 1119 69902 1128
rect 70492 1148 70544 1154
rect 69860 1018 69888 1119
rect 70492 1090 70544 1096
rect 69848 1012 69900 1018
rect 69848 954 69900 960
rect 68284 750 68336 756
rect 69400 746 69704 762
rect 70504 746 70532 1090
rect 71424 950 71452 2246
rect 71504 1352 71556 1358
rect 71504 1294 71556 1300
rect 71412 944 71464 950
rect 71412 886 71464 892
rect 71516 814 71544 1294
rect 71792 1018 71820 2858
rect 73160 2848 73212 2854
rect 73160 2790 73212 2796
rect 73172 2446 73200 2790
rect 74000 2650 74028 4762
rect 74736 3534 74764 9386
rect 78680 6928 78732 6934
rect 78680 6870 78732 6876
rect 75920 5840 75972 5846
rect 75920 5782 75972 5788
rect 75932 4078 75960 5782
rect 78692 5166 78720 6870
rect 78680 5160 78732 5166
rect 78680 5102 78732 5108
rect 76564 5092 76616 5098
rect 76564 5034 76616 5040
rect 75920 4072 75972 4078
rect 75920 4014 75972 4020
rect 76472 4004 76524 4010
rect 76472 3946 76524 3952
rect 74724 3528 74776 3534
rect 74724 3470 74776 3476
rect 76484 3466 76512 3946
rect 76472 3460 76524 3466
rect 76472 3402 76524 3408
rect 74540 3120 74592 3126
rect 74540 3062 74592 3068
rect 73988 2644 74040 2650
rect 73988 2586 74040 2592
rect 73160 2440 73212 2446
rect 73160 2382 73212 2388
rect 72148 2304 72200 2310
rect 72148 2246 72200 2252
rect 72160 1737 72188 2246
rect 72146 1728 72202 1737
rect 72146 1663 72202 1672
rect 73172 1170 73200 2382
rect 74552 1562 74580 3062
rect 76576 2650 76604 5034
rect 81714 4720 81770 4729
rect 79232 4684 79284 4690
rect 81714 4655 81770 4664
rect 79232 4626 79284 4632
rect 79048 4072 79100 4078
rect 79048 4014 79100 4020
rect 79060 3466 79088 4014
rect 76656 3460 76708 3466
rect 76656 3402 76708 3408
rect 79048 3460 79100 3466
rect 79048 3402 79100 3408
rect 76668 2922 76696 3402
rect 78496 3392 78548 3398
rect 78496 3334 78548 3340
rect 78508 3126 78536 3334
rect 78496 3120 78548 3126
rect 78496 3062 78548 3068
rect 78680 3120 78732 3126
rect 78680 3062 78732 3068
rect 76656 2916 76708 2922
rect 76656 2858 76708 2864
rect 76564 2644 76616 2650
rect 76564 2586 76616 2592
rect 75552 2440 75604 2446
rect 75552 2382 75604 2388
rect 75460 2304 75512 2310
rect 75460 2246 75512 2252
rect 74908 1896 74960 1902
rect 74908 1838 74960 1844
rect 74540 1556 74592 1562
rect 74540 1498 74592 1504
rect 73356 1426 73660 1442
rect 73356 1420 73672 1426
rect 73356 1414 73620 1420
rect 73356 1358 73384 1414
rect 73620 1362 73672 1368
rect 74920 1358 74948 1838
rect 73344 1352 73396 1358
rect 74908 1352 74960 1358
rect 73344 1294 73396 1300
rect 73448 1290 73660 1306
rect 74908 1294 74960 1300
rect 75000 1352 75052 1358
rect 75000 1294 75052 1300
rect 73436 1284 73672 1290
rect 73488 1278 73620 1284
rect 73436 1226 73488 1232
rect 73620 1226 73672 1232
rect 73080 1142 73200 1170
rect 73080 1034 73108 1142
rect 72896 1018 73108 1034
rect 73160 1080 73212 1086
rect 73160 1022 73212 1028
rect 71780 1012 71832 1018
rect 71780 954 71832 960
rect 72884 1012 73108 1018
rect 72936 1006 73108 1012
rect 72884 954 72936 960
rect 73068 944 73120 950
rect 72896 892 73068 898
rect 72896 886 73120 892
rect 72896 882 73108 886
rect 73172 882 73200 1022
rect 72884 876 73108 882
rect 72936 870 73108 876
rect 73160 876 73212 882
rect 72884 818 72936 824
rect 73160 818 73212 824
rect 71504 808 71556 814
rect 71504 750 71556 756
rect 69388 740 69704 746
rect 69440 734 69704 740
rect 70492 740 70544 746
rect 69388 682 69440 688
rect 70492 682 70544 688
rect 67568 248 67580 304
rect 67636 248 67660 304
rect 67716 248 67740 304
rect 67796 248 67820 304
rect 67876 248 67888 304
rect 67568 224 67888 248
rect 67568 168 67580 224
rect 67636 168 67660 224
rect 67716 168 67740 224
rect 67796 168 67820 224
rect 67876 168 67888 224
rect 67568 144 67888 168
rect 67568 88 67580 144
rect 67636 88 67660 144
rect 67716 88 67740 144
rect 67796 88 67820 144
rect 67876 88 67888 144
rect 67568 64 67888 88
rect 75012 66 75040 1294
rect 75472 1290 75500 2246
rect 75564 1766 75592 2382
rect 77300 2304 77352 2310
rect 77300 2246 77352 2252
rect 75552 1760 75604 1766
rect 75552 1702 75604 1708
rect 75644 1760 75696 1766
rect 75644 1702 75696 1708
rect 75460 1284 75512 1290
rect 75460 1226 75512 1232
rect 75656 1086 75684 1702
rect 75736 1556 75788 1562
rect 75736 1498 75788 1504
rect 75748 1154 75776 1498
rect 77312 1306 77340 2246
rect 78692 1902 78720 3062
rect 79244 2446 79272 4626
rect 81532 3392 81584 3398
rect 81532 3334 81584 3340
rect 80060 2916 80112 2922
rect 80060 2858 80112 2864
rect 79232 2440 79284 2446
rect 79232 2382 79284 2388
rect 79876 2304 79928 2310
rect 79876 2246 79928 2252
rect 78680 1896 78732 1902
rect 78680 1838 78732 1844
rect 79888 1601 79916 2246
rect 79874 1592 79930 1601
rect 79874 1527 79930 1536
rect 77220 1290 77340 1306
rect 78036 1352 78088 1358
rect 78036 1294 78088 1300
rect 77208 1284 77340 1290
rect 77260 1278 77340 1284
rect 77208 1226 77260 1232
rect 75736 1148 75788 1154
rect 75736 1090 75788 1096
rect 75828 1148 75880 1154
rect 75828 1090 75880 1096
rect 75644 1080 75696 1086
rect 75840 1034 75868 1090
rect 75644 1022 75696 1028
rect 75748 1006 75868 1034
rect 75748 814 75776 1006
rect 75840 882 76604 898
rect 75828 876 76616 882
rect 75880 870 76564 876
rect 75828 818 75880 824
rect 76564 818 76616 824
rect 78048 814 78076 1294
rect 79140 1284 79192 1290
rect 79140 1226 79192 1232
rect 79152 814 79180 1226
rect 80072 1086 80100 2858
rect 81440 2848 81492 2854
rect 81440 2790 81492 2796
rect 81452 2378 81480 2790
rect 81440 2372 81492 2378
rect 81440 2314 81492 2320
rect 80244 1896 80296 1902
rect 80244 1838 80296 1844
rect 80152 1760 80204 1766
rect 80152 1702 80204 1708
rect 80164 1290 80192 1702
rect 80152 1284 80204 1290
rect 80152 1226 80204 1232
rect 80060 1080 80112 1086
rect 80060 1022 80112 1028
rect 80256 814 80284 1838
rect 80336 1760 80388 1766
rect 80336 1702 80388 1708
rect 80348 950 80376 1702
rect 81346 1184 81402 1193
rect 81346 1119 81348 1128
rect 81400 1119 81402 1128
rect 81348 1090 81400 1096
rect 81452 950 81480 2314
rect 81544 1562 81572 3334
rect 81728 2650 81756 4655
rect 81900 3528 81952 3534
rect 81900 3470 81952 3476
rect 81912 3398 81940 3470
rect 82464 3466 82492 9454
rect 90180 9376 90232 9382
rect 90180 9318 90232 9324
rect 87604 9172 87656 9178
rect 87604 9114 87656 9120
rect 85580 8288 85632 8294
rect 85580 8230 85632 8236
rect 82820 5160 82872 5166
rect 82820 5102 82872 5108
rect 82452 3460 82504 3466
rect 82452 3402 82504 3408
rect 81900 3392 81952 3398
rect 81900 3334 81952 3340
rect 82832 3194 82860 5102
rect 84292 4140 84344 4146
rect 84292 4082 84344 4088
rect 84304 3398 84332 4082
rect 83648 3392 83700 3398
rect 83648 3334 83700 3340
rect 84292 3392 84344 3398
rect 84292 3334 84344 3340
rect 82820 3188 82872 3194
rect 82820 3130 82872 3136
rect 83660 3126 83688 3334
rect 83648 3120 83700 3126
rect 83648 3062 83700 3068
rect 85592 2990 85620 8230
rect 86316 7880 86368 7886
rect 86368 7828 86632 7834
rect 86316 7822 86632 7828
rect 86328 7806 86632 7822
rect 86604 7750 86632 7806
rect 86592 7744 86644 7750
rect 86592 7686 86644 7692
rect 86960 3460 87012 3466
rect 86960 3402 87012 3408
rect 86868 3392 86920 3398
rect 86868 3334 86920 3340
rect 86880 3126 86908 3334
rect 86868 3120 86920 3126
rect 86868 3062 86920 3068
rect 85580 2984 85632 2990
rect 85580 2926 85632 2932
rect 86972 2922 87000 3402
rect 87420 3392 87472 3398
rect 87420 3334 87472 3340
rect 86960 2916 87012 2922
rect 86960 2858 87012 2864
rect 84016 2848 84068 2854
rect 84016 2790 84068 2796
rect 81716 2644 81768 2650
rect 81716 2586 81768 2592
rect 84028 2394 84056 2790
rect 84028 2378 84148 2394
rect 84028 2372 84160 2378
rect 84028 2366 84108 2372
rect 84108 2314 84160 2320
rect 86776 2372 86828 2378
rect 86776 2314 86828 2320
rect 81532 1556 81584 1562
rect 81532 1498 81584 1504
rect 84120 1290 84148 2314
rect 84292 2304 84344 2310
rect 84292 2246 84344 2252
rect 84476 2304 84528 2310
rect 84476 2246 84528 2252
rect 84304 1562 84332 2246
rect 84292 1556 84344 1562
rect 84292 1498 84344 1504
rect 84108 1284 84160 1290
rect 84108 1226 84160 1232
rect 84014 1184 84070 1193
rect 84488 1154 84516 2246
rect 86788 1426 86816 2314
rect 86960 2304 87012 2310
rect 86960 2246 87012 2252
rect 86972 1766 87000 2246
rect 86960 1760 87012 1766
rect 86960 1702 87012 1708
rect 87052 1760 87104 1766
rect 87052 1702 87104 1708
rect 86776 1420 86828 1426
rect 86776 1362 86828 1368
rect 86866 1320 86922 1329
rect 85764 1284 85816 1290
rect 86866 1255 86922 1264
rect 85764 1226 85816 1232
rect 84014 1119 84070 1128
rect 84476 1148 84528 1154
rect 82452 1080 82504 1086
rect 82452 1022 82504 1028
rect 80336 944 80388 950
rect 80336 886 80388 892
rect 81440 944 81492 950
rect 81440 886 81492 892
rect 82464 814 82492 1022
rect 84028 882 84056 1119
rect 84476 1090 84528 1096
rect 84660 1148 84712 1154
rect 84660 1090 84712 1096
rect 84016 876 84068 882
rect 84016 818 84068 824
rect 75736 808 75788 814
rect 75736 750 75788 756
rect 78036 808 78088 814
rect 78036 750 78088 756
rect 79140 808 79192 814
rect 79140 750 79192 756
rect 80244 808 80296 814
rect 80244 750 80296 756
rect 82452 808 82504 814
rect 82452 750 82504 756
rect 84672 746 84700 1090
rect 85776 814 85804 1226
rect 86880 1086 86908 1255
rect 87064 1222 87092 1702
rect 87326 1456 87382 1465
rect 87326 1391 87382 1400
rect 87052 1216 87104 1222
rect 87052 1158 87104 1164
rect 86868 1080 86920 1086
rect 86868 1022 86920 1028
rect 86960 1012 87012 1018
rect 87340 1000 87368 1391
rect 87012 972 87368 1000
rect 86960 954 87012 960
rect 86914 876 86966 882
rect 87432 864 87460 3334
rect 87616 2650 87644 9114
rect 90192 3534 90220 9318
rect 91296 7942 91876 7970
rect 91296 7818 91324 7942
rect 91376 7880 91428 7886
rect 91376 7822 91428 7828
rect 91284 7812 91336 7818
rect 91284 7754 91336 7760
rect 91388 7698 91416 7822
rect 91848 7818 91876 7942
rect 91836 7812 91888 7818
rect 91836 7754 91888 7760
rect 91744 7744 91796 7750
rect 91388 7692 91744 7698
rect 91388 7686 91796 7692
rect 91388 7670 91784 7686
rect 90548 7200 90600 7206
rect 90548 7142 90600 7148
rect 90560 7002 90588 7142
rect 90548 6996 90600 7002
rect 90548 6938 90600 6944
rect 92124 6798 92152 9930
rect 92216 7410 92244 11902
rect 100668 11892 100720 11898
rect 100668 11834 100720 11840
rect 99932 11688 99984 11694
rect 99932 11630 99984 11636
rect 97448 11484 97500 11490
rect 97448 11426 97500 11432
rect 92848 11280 92900 11286
rect 92848 11222 92900 11228
rect 92860 7818 92888 11222
rect 97264 10940 97316 10946
rect 97264 10882 97316 10888
rect 96068 10804 96120 10810
rect 96068 10746 96120 10752
rect 95148 10260 95200 10266
rect 95148 10202 95200 10208
rect 93768 10056 93820 10062
rect 93768 9998 93820 10004
rect 93490 7984 93546 7993
rect 93490 7919 93546 7928
rect 92848 7812 92900 7818
rect 92848 7754 92900 7760
rect 93504 7410 93532 7919
rect 92204 7404 92256 7410
rect 92204 7346 92256 7352
rect 93492 7404 93544 7410
rect 93492 7346 93544 7352
rect 92388 7336 92440 7342
rect 92388 7278 92440 7284
rect 92296 7200 92348 7206
rect 92296 7142 92348 7148
rect 92308 6934 92336 7142
rect 92296 6928 92348 6934
rect 92296 6870 92348 6876
rect 92112 6792 92164 6798
rect 92112 6734 92164 6740
rect 90916 6656 90968 6662
rect 90916 6598 90968 6604
rect 90928 6458 90956 6598
rect 90916 6452 90968 6458
rect 90916 6394 90968 6400
rect 92400 5302 92428 7278
rect 93780 6798 93808 9998
rect 94044 7744 94096 7750
rect 94044 7686 94096 7692
rect 94056 7342 94084 7686
rect 94044 7336 94096 7342
rect 94044 7278 94096 7284
rect 94872 7336 94924 7342
rect 94872 7278 94924 7284
rect 94884 7002 94912 7278
rect 94872 6996 94924 7002
rect 94872 6938 94924 6944
rect 94504 6928 94556 6934
rect 94504 6870 94556 6876
rect 93768 6792 93820 6798
rect 93768 6734 93820 6740
rect 94320 6792 94372 6798
rect 94320 6734 94372 6740
rect 92756 6656 92808 6662
rect 92756 6598 92808 6604
rect 92388 5296 92440 5302
rect 92388 5238 92440 5244
rect 92768 4690 92796 6598
rect 94332 6118 94360 6734
rect 94320 6112 94372 6118
rect 94320 6054 94372 6060
rect 94332 4758 94360 6054
rect 94516 5234 94544 6870
rect 95160 6798 95188 10202
rect 95240 7744 95292 7750
rect 95240 7686 95292 7692
rect 95252 7478 95280 7686
rect 96080 7478 96108 10746
rect 96712 7880 96764 7886
rect 96712 7822 96764 7828
rect 95240 7472 95292 7478
rect 95240 7414 95292 7420
rect 96068 7472 96120 7478
rect 96068 7414 96120 7420
rect 96724 7410 96752 7822
rect 97276 7478 97304 10882
rect 97264 7472 97316 7478
rect 97264 7414 97316 7420
rect 96712 7404 96764 7410
rect 96712 7346 96764 7352
rect 96620 7336 96672 7342
rect 96620 7278 96672 7284
rect 95148 6792 95200 6798
rect 95148 6734 95200 6740
rect 96632 5370 96660 7278
rect 96712 7200 96764 7206
rect 96712 7142 96764 7148
rect 96620 5364 96672 5370
rect 96620 5306 96672 5312
rect 94504 5228 94556 5234
rect 94504 5170 94556 5176
rect 94320 4752 94372 4758
rect 94320 4694 94372 4700
rect 92756 4684 92808 4690
rect 92756 4626 92808 4632
rect 94136 4684 94188 4690
rect 94136 4626 94188 4632
rect 92386 4584 92442 4593
rect 91560 4548 91612 4554
rect 92386 4519 92442 4528
rect 91560 4490 91612 4496
rect 89628 3528 89680 3534
rect 89720 3528 89772 3534
rect 89680 3476 89720 3482
rect 89628 3470 89772 3476
rect 90180 3528 90232 3534
rect 90180 3470 90232 3476
rect 89640 3454 89760 3470
rect 91572 3126 91600 4490
rect 92112 3460 92164 3466
rect 92112 3402 92164 3408
rect 92020 3392 92072 3398
rect 92020 3334 92072 3340
rect 91560 3120 91612 3126
rect 91560 3062 91612 3068
rect 92032 2922 92060 3334
rect 92020 2916 92072 2922
rect 92020 2858 92072 2864
rect 92124 2854 92152 3402
rect 89536 2848 89588 2854
rect 89536 2790 89588 2796
rect 89720 2848 89772 2854
rect 89720 2790 89772 2796
rect 92112 2848 92164 2854
rect 92112 2790 92164 2796
rect 87604 2644 87656 2650
rect 87604 2586 87656 2592
rect 87616 2446 87644 2586
rect 87604 2440 87656 2446
rect 87604 2382 87656 2388
rect 89548 2378 89576 2790
rect 89536 2372 89588 2378
rect 89536 2314 89588 2320
rect 89732 1358 89760 2790
rect 92400 2650 92428 4519
rect 92572 3392 92624 3398
rect 92572 3334 92624 3340
rect 92388 2644 92440 2650
rect 92388 2586 92440 2592
rect 91284 2304 91336 2310
rect 91284 2246 91336 2252
rect 92296 2304 92348 2310
rect 92296 2246 92348 2252
rect 89812 1896 89864 1902
rect 89812 1838 89864 1844
rect 89824 1358 89852 1838
rect 89720 1352 89772 1358
rect 89720 1294 89772 1300
rect 89812 1352 89864 1358
rect 89812 1294 89864 1300
rect 89904 1284 89956 1290
rect 89904 1226 89956 1232
rect 89812 1216 89864 1222
rect 89916 1170 89944 1226
rect 89864 1164 89944 1170
rect 89812 1158 89944 1164
rect 89824 1142 89944 1158
rect 90178 1184 90234 1193
rect 90178 1119 90234 1128
rect 87880 1080 87932 1086
rect 87880 1022 87932 1028
rect 86966 836 87460 864
rect 86914 818 86966 824
rect 87892 814 87920 1022
rect 90192 1018 90220 1119
rect 90180 1012 90232 1018
rect 90180 954 90232 960
rect 90272 1012 90324 1018
rect 90272 954 90324 960
rect 90284 898 90312 954
rect 91296 950 91324 2246
rect 91836 1896 91888 1902
rect 91836 1838 91888 1844
rect 90100 870 90312 898
rect 91284 944 91336 950
rect 91284 886 91336 892
rect 91376 944 91428 950
rect 91376 886 91428 892
rect 90100 814 90128 870
rect 91388 814 91416 886
rect 91848 882 91876 1838
rect 92308 1766 92336 2246
rect 92296 1760 92348 1766
rect 92296 1702 92348 1708
rect 92584 1358 92612 3334
rect 94148 2446 94176 4626
rect 96724 4622 96752 7142
rect 97460 6798 97488 11426
rect 98460 11144 98512 11150
rect 98460 11086 98512 11092
rect 97632 7744 97684 7750
rect 97632 7686 97684 7692
rect 97644 7546 97672 7686
rect 97632 7540 97684 7546
rect 97632 7482 97684 7488
rect 98472 7478 98500 11086
rect 99472 7948 99524 7954
rect 99472 7890 99524 7896
rect 98460 7472 98512 7478
rect 98460 7414 98512 7420
rect 99484 7410 99512 7890
rect 99472 7404 99524 7410
rect 99472 7346 99524 7352
rect 96804 6792 96856 6798
rect 96804 6734 96856 6740
rect 97448 6792 97500 6798
rect 97448 6734 97500 6740
rect 96816 6118 96844 6734
rect 98368 6656 98420 6662
rect 98368 6598 98420 6604
rect 96804 6112 96856 6118
rect 96804 6054 96856 6060
rect 96712 4616 96764 4622
rect 96712 4558 96764 4564
rect 94596 3392 94648 3398
rect 94596 3334 94648 3340
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 94608 3194 94636 3334
rect 94596 3188 94648 3194
rect 94596 3130 94648 3136
rect 94136 2440 94188 2446
rect 94136 2382 94188 2388
rect 94596 1692 94648 1698
rect 94596 1634 94648 1640
rect 94608 1442 94636 1634
rect 94136 1420 94188 1426
rect 94136 1362 94188 1368
rect 94332 1414 94636 1442
rect 92572 1352 92624 1358
rect 92572 1294 92624 1300
rect 93308 1148 93360 1154
rect 93308 1090 93360 1096
rect 92204 1080 92256 1086
rect 92204 1022 92256 1028
rect 91836 876 91888 882
rect 91836 818 91888 824
rect 92216 814 92244 1022
rect 93320 814 93348 1090
rect 94148 1018 94176 1362
rect 94332 1086 94360 1414
rect 94792 1329 94820 3334
rect 96712 3120 96764 3126
rect 96712 3062 96764 3068
rect 96620 2848 96672 2854
rect 96620 2790 96672 2796
rect 95332 2440 95384 2446
rect 95332 2382 95384 2388
rect 95344 1873 95372 2382
rect 96632 2378 96660 2790
rect 96620 2372 96672 2378
rect 96620 2314 96672 2320
rect 95330 1864 95386 1873
rect 95330 1799 95386 1808
rect 96632 1465 96660 2314
rect 96618 1456 96674 1465
rect 96618 1391 96674 1400
rect 95516 1352 95568 1358
rect 94778 1320 94834 1329
rect 95516 1294 95568 1300
rect 94778 1255 94834 1264
rect 94320 1080 94372 1086
rect 94320 1022 94372 1028
rect 94688 1080 94740 1086
rect 94688 1022 94740 1028
rect 94136 1012 94188 1018
rect 94136 954 94188 960
rect 94320 944 94372 950
rect 94596 944 94648 950
rect 94372 904 94596 932
rect 94320 886 94372 892
rect 94596 886 94648 892
rect 85764 808 85816 814
rect 85764 750 85816 756
rect 87880 808 87932 814
rect 87880 750 87932 756
rect 90088 808 90140 814
rect 90088 750 90140 756
rect 91376 808 91428 814
rect 91376 750 91428 756
rect 92204 808 92256 814
rect 92204 750 92256 756
rect 93308 808 93360 814
rect 93308 750 93360 756
rect 84660 740 84712 746
rect 84660 682 84712 688
rect 87236 740 87288 746
rect 87236 682 87288 688
rect 87248 626 87276 682
rect 86880 610 87276 626
rect 86868 604 87276 610
rect 86920 598 87276 604
rect 86868 546 86920 552
rect 89168 536 89220 542
rect 89166 504 89168 513
rect 94700 513 94728 1022
rect 95528 814 95556 1294
rect 96724 1193 96752 3062
rect 96816 1834 96844 6054
rect 98380 5778 98408 6598
rect 99944 6390 99972 11630
rect 100680 7410 100708 11834
rect 175464 11824 175516 11830
rect 175464 11766 175516 11772
rect 195244 11824 195296 11830
rect 195244 11766 195296 11772
rect 107568 11756 107620 11762
rect 107568 11698 107620 11704
rect 104072 11076 104124 11082
rect 104072 11018 104124 11024
rect 102876 10872 102928 10878
rect 102876 10814 102928 10820
rect 101956 10736 102008 10742
rect 101956 10678 102008 10684
rect 101862 8120 101918 8129
rect 101312 8084 101364 8090
rect 101862 8055 101918 8064
rect 101312 8026 101364 8032
rect 101324 7410 101352 8026
rect 101876 7478 101904 8055
rect 101864 7472 101916 7478
rect 101864 7414 101916 7420
rect 100668 7404 100720 7410
rect 100668 7346 100720 7352
rect 101312 7404 101364 7410
rect 101312 7346 101364 7352
rect 100668 6724 100720 6730
rect 100668 6666 100720 6672
rect 99932 6384 99984 6390
rect 99932 6326 99984 6332
rect 100576 6316 100628 6322
rect 100576 6258 100628 6264
rect 100588 6118 100616 6258
rect 99564 6112 99616 6118
rect 99564 6054 99616 6060
rect 100576 6112 100628 6118
rect 100576 6054 100628 6060
rect 98368 5772 98420 5778
rect 98368 5714 98420 5720
rect 98644 5704 98696 5710
rect 98644 5646 98696 5652
rect 97172 4752 97224 4758
rect 97172 4694 97224 4700
rect 97184 2650 97212 4694
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 97920 3398 97948 3470
rect 97908 3392 97960 3398
rect 97908 3334 97960 3340
rect 97172 2644 97224 2650
rect 97172 2586 97224 2592
rect 96804 1828 96856 1834
rect 96804 1770 96856 1776
rect 97448 1828 97500 1834
rect 97448 1770 97500 1776
rect 96710 1184 96766 1193
rect 96710 1119 96766 1128
rect 97460 882 97488 1770
rect 97538 1320 97594 1329
rect 97538 1255 97594 1264
rect 97552 950 97580 1255
rect 97920 1193 97948 3334
rect 98656 2106 98684 5646
rect 99104 3392 99156 3398
rect 99104 3334 99156 3340
rect 99116 3126 99144 3334
rect 99104 3120 99156 3126
rect 99104 3062 99156 3068
rect 99472 2848 99524 2854
rect 99472 2790 99524 2796
rect 99104 2644 99156 2650
rect 99104 2586 99156 2592
rect 99010 2272 99066 2281
rect 99010 2207 99066 2216
rect 98644 2100 98696 2106
rect 98644 2042 98696 2048
rect 98826 1456 98882 1465
rect 98826 1391 98882 1400
rect 97906 1184 97962 1193
rect 97906 1119 97962 1128
rect 97540 944 97592 950
rect 97540 886 97592 892
rect 97448 876 97500 882
rect 97448 818 97500 824
rect 98840 814 98868 1391
rect 99024 1358 99052 2207
rect 99012 1352 99064 1358
rect 99012 1294 99064 1300
rect 99116 1290 99144 2586
rect 99196 2440 99248 2446
rect 99196 2382 99248 2388
rect 99104 1284 99156 1290
rect 99104 1226 99156 1232
rect 99208 1222 99236 2382
rect 99484 2378 99512 2790
rect 99472 2372 99524 2378
rect 99472 2314 99524 2320
rect 99378 2000 99434 2009
rect 99378 1935 99434 1944
rect 99196 1216 99248 1222
rect 99196 1158 99248 1164
rect 99392 1018 99420 1935
rect 99576 1766 99604 6054
rect 99748 3392 99800 3398
rect 99748 3334 99800 3340
rect 99760 3126 99788 3334
rect 99748 3120 99800 3126
rect 99748 3062 99800 3068
rect 99748 2304 99800 2310
rect 99748 2246 99800 2252
rect 99760 2106 99788 2246
rect 99748 2100 99800 2106
rect 99748 2042 99800 2048
rect 99564 1760 99616 1766
rect 99564 1702 99616 1708
rect 100024 1216 100076 1222
rect 100024 1158 100076 1164
rect 100680 1170 100708 6666
rect 101220 6656 101272 6662
rect 101220 6598 101272 6604
rect 100852 3052 100904 3058
rect 100852 2994 100904 3000
rect 100864 2774 100892 2994
rect 101232 2990 101260 6598
rect 101968 6390 101996 10678
rect 102232 7268 102284 7274
rect 102232 7210 102284 7216
rect 102244 6934 102272 7210
rect 102232 6928 102284 6934
rect 102232 6870 102284 6876
rect 102888 6866 102916 10814
rect 103058 9208 103114 9217
rect 103058 9143 103114 9152
rect 102876 6860 102928 6866
rect 102876 6802 102928 6808
rect 101956 6384 102008 6390
rect 101956 6326 102008 6332
rect 102600 6316 102652 6322
rect 102600 6258 102652 6264
rect 102612 6118 102640 6258
rect 102600 6112 102652 6118
rect 102600 6054 102652 6060
rect 102612 5914 102640 6054
rect 102600 5908 102652 5914
rect 102600 5850 102652 5856
rect 102324 4480 102376 4486
rect 102324 4422 102376 4428
rect 102140 3460 102192 3466
rect 102140 3402 102192 3408
rect 101220 2984 101272 2990
rect 101220 2926 101272 2932
rect 102152 2854 102180 3402
rect 102336 3398 102364 4422
rect 102324 3392 102376 3398
rect 102324 3334 102376 3340
rect 102508 3392 102560 3398
rect 102508 3334 102560 3340
rect 102140 2848 102192 2854
rect 102140 2790 102192 2796
rect 100772 2746 100892 2774
rect 100772 1329 100800 2746
rect 102152 1902 102180 2790
rect 102140 1896 102192 1902
rect 102140 1838 102192 1844
rect 102232 1896 102284 1902
rect 102232 1838 102284 1844
rect 102244 1578 102272 1838
rect 102060 1550 102272 1578
rect 101126 1456 101182 1465
rect 101126 1391 101182 1400
rect 101140 1358 101168 1391
rect 101128 1352 101180 1358
rect 100758 1320 100814 1329
rect 100758 1255 100814 1264
rect 100942 1320 100998 1329
rect 101128 1294 101180 1300
rect 100942 1255 100998 1264
rect 100956 1170 100984 1255
rect 100036 1034 100064 1158
rect 100680 1142 100984 1170
rect 99380 1012 99432 1018
rect 99380 954 99432 960
rect 99852 1006 100064 1034
rect 100944 1012 100996 1018
rect 99852 898 99880 1006
rect 100944 954 100996 960
rect 99760 870 99880 898
rect 99760 814 99788 870
rect 95516 808 95568 814
rect 95516 750 95568 756
rect 98828 808 98880 814
rect 98828 750 98880 756
rect 99748 808 99800 814
rect 99748 750 99800 756
rect 100956 746 100984 954
rect 102060 814 102088 1550
rect 102520 1086 102548 3334
rect 103072 2650 103100 9143
rect 103244 7200 103296 7206
rect 103244 7142 103296 7148
rect 103256 6798 103284 7142
rect 104084 6866 104112 11018
rect 106188 10600 106240 10606
rect 106188 10542 106240 10548
rect 104072 6860 104124 6866
rect 104072 6802 104124 6808
rect 103244 6792 103296 6798
rect 103244 6734 103296 6740
rect 104440 6792 104492 6798
rect 104440 6734 104492 6740
rect 103704 6656 103756 6662
rect 103704 6598 103756 6604
rect 103716 6254 103744 6598
rect 103704 6248 103756 6254
rect 103704 6190 103756 6196
rect 103796 6248 103848 6254
rect 103796 6190 103848 6196
rect 103808 5846 103836 6190
rect 104452 6118 104480 6734
rect 106200 6390 106228 10542
rect 107292 6724 107344 6730
rect 107292 6666 107344 6672
rect 107304 6458 107332 6666
rect 107292 6452 107344 6458
rect 107292 6394 107344 6400
rect 106188 6384 106240 6390
rect 106188 6326 106240 6332
rect 106924 6316 106976 6322
rect 106924 6258 106976 6264
rect 104440 6112 104492 6118
rect 104440 6054 104492 6060
rect 105084 6112 105136 6118
rect 105084 6054 105136 6060
rect 103796 5840 103848 5846
rect 103796 5782 103848 5788
rect 104452 3505 104480 6054
rect 105096 5574 105124 6054
rect 106936 5642 106964 6258
rect 107580 5778 107608 11698
rect 157892 11552 157944 11558
rect 157892 11494 157944 11500
rect 123116 11212 123168 11218
rect 123116 11154 123168 11160
rect 109868 10532 109920 10538
rect 109868 10474 109920 10480
rect 109500 6860 109552 6866
rect 109500 6802 109552 6808
rect 109512 6254 109540 6802
rect 109776 6316 109828 6322
rect 109776 6258 109828 6264
rect 109500 6248 109552 6254
rect 109500 6190 109552 6196
rect 109788 6118 109816 6258
rect 109776 6112 109828 6118
rect 109776 6054 109828 6060
rect 107568 5772 107620 5778
rect 107568 5714 107620 5720
rect 106924 5636 106976 5642
rect 106924 5578 106976 5584
rect 105084 5568 105136 5574
rect 105084 5510 105136 5516
rect 107660 5568 107712 5574
rect 108764 5568 108816 5574
rect 107660 5510 107712 5516
rect 108684 5528 108764 5556
rect 105084 3528 105136 3534
rect 104438 3496 104494 3505
rect 104438 3431 104494 3440
rect 105082 3496 105084 3505
rect 105136 3496 105138 3505
rect 105082 3431 105138 3440
rect 105634 3496 105690 3505
rect 105634 3431 105636 3440
rect 105688 3431 105690 3440
rect 107568 3460 107620 3466
rect 105636 3402 105688 3408
rect 107568 3402 107620 3408
rect 107476 3392 107528 3398
rect 107476 3334 107528 3340
rect 107488 2990 107516 3334
rect 107580 3058 107608 3402
rect 107568 3052 107620 3058
rect 107568 2994 107620 3000
rect 107476 2984 107528 2990
rect 107476 2926 107528 2932
rect 104624 2848 104676 2854
rect 104624 2790 104676 2796
rect 107384 2848 107436 2854
rect 107384 2790 107436 2796
rect 103060 2644 103112 2650
rect 103060 2586 103112 2592
rect 103428 2644 103480 2650
rect 103428 2586 103480 2592
rect 103072 2446 103100 2586
rect 103060 2440 103112 2446
rect 103060 2382 103112 2388
rect 103440 1766 103468 2586
rect 104164 2576 104216 2582
rect 103992 2524 104164 2530
rect 103992 2518 104216 2524
rect 103992 2514 104204 2518
rect 103980 2508 104204 2514
rect 104032 2502 104204 2508
rect 103980 2450 104032 2456
rect 104636 2378 104664 2790
rect 107396 2582 107424 2790
rect 107384 2576 107436 2582
rect 107384 2518 107436 2524
rect 107672 2514 107700 5510
rect 107844 2644 107896 2650
rect 107844 2586 107896 2592
rect 107936 2644 107988 2650
rect 107936 2586 107988 2592
rect 107856 2514 107884 2586
rect 107660 2508 107712 2514
rect 107660 2450 107712 2456
rect 107844 2508 107896 2514
rect 107844 2450 107896 2456
rect 104624 2372 104676 2378
rect 104624 2314 104676 2320
rect 104900 2304 104952 2310
rect 104900 2246 104952 2252
rect 106372 2304 106424 2310
rect 106372 2246 106424 2252
rect 107752 2304 107804 2310
rect 107752 2246 107804 2252
rect 103428 1760 103480 1766
rect 103428 1702 103480 1708
rect 104912 1630 104940 2246
rect 104900 1624 104952 1630
rect 104900 1566 104952 1572
rect 105268 1420 105320 1426
rect 105268 1362 105320 1368
rect 102508 1080 102560 1086
rect 102508 1022 102560 1028
rect 104164 1080 104216 1086
rect 104164 1022 104216 1028
rect 103612 876 103664 882
rect 103612 818 103664 824
rect 102048 808 102100 814
rect 102048 750 102100 756
rect 100944 740 100996 746
rect 100944 682 100996 688
rect 103624 513 103652 818
rect 104176 814 104204 1022
rect 105280 814 105308 1362
rect 106384 1290 106412 2246
rect 107476 1760 107528 1766
rect 107476 1702 107528 1708
rect 106372 1284 106424 1290
rect 106372 1226 106424 1232
rect 106556 1284 106608 1290
rect 106556 1226 106608 1232
rect 106568 814 106596 1226
rect 107488 814 107516 1702
rect 107764 1426 107792 2246
rect 107948 1902 107976 2586
rect 108684 2038 108712 5528
rect 108764 5510 108816 5516
rect 109684 3596 109736 3602
rect 109684 3538 109736 3544
rect 109132 3392 109184 3398
rect 109132 3334 109184 3340
rect 109040 2644 109092 2650
rect 109040 2586 109092 2592
rect 108672 2032 108724 2038
rect 108672 1974 108724 1980
rect 108764 2032 108816 2038
rect 108764 1974 108816 1980
rect 107936 1896 107988 1902
rect 107936 1838 107988 1844
rect 108302 1456 108358 1465
rect 107752 1420 107804 1426
rect 108302 1391 108358 1400
rect 107752 1362 107804 1368
rect 108316 882 108344 1391
rect 108304 876 108356 882
rect 108304 818 108356 824
rect 108776 814 108804 1974
rect 109052 1358 109080 2586
rect 109040 1352 109092 1358
rect 108854 1320 108910 1329
rect 108910 1278 108988 1306
rect 109040 1294 109092 1300
rect 108854 1255 108910 1264
rect 108960 1154 108988 1278
rect 108856 1148 108908 1154
rect 108856 1090 108908 1096
rect 108948 1148 109000 1154
rect 108948 1090 109000 1096
rect 104164 808 104216 814
rect 104164 750 104216 756
rect 105268 808 105320 814
rect 105268 750 105320 756
rect 106556 808 106608 814
rect 106556 750 106608 756
rect 107476 808 107528 814
rect 107476 750 107528 756
rect 108764 808 108816 814
rect 108764 750 108816 756
rect 108868 513 108896 1090
rect 109144 513 109172 3334
rect 109696 3058 109724 3538
rect 109684 3052 109736 3058
rect 109684 2994 109736 3000
rect 109788 2446 109816 6054
rect 109880 5710 109908 10474
rect 122564 10464 122616 10470
rect 122564 10406 122616 10412
rect 112812 10124 112864 10130
rect 112812 10066 112864 10072
rect 110788 9104 110840 9110
rect 110788 9046 110840 9052
rect 109868 5704 109920 5710
rect 109868 5646 109920 5652
rect 109960 4276 110012 4282
rect 109960 4218 110012 4224
rect 109972 3670 110000 4218
rect 109960 3664 110012 3670
rect 109960 3606 110012 3612
rect 110800 2650 110828 9046
rect 112824 6866 112852 10066
rect 122576 8090 122604 10406
rect 122564 8084 122616 8090
rect 122564 8026 122616 8032
rect 121000 7948 121052 7954
rect 121000 7890 121052 7896
rect 114836 7880 114888 7886
rect 114836 7822 114888 7828
rect 113640 7812 113692 7818
rect 113640 7754 113692 7760
rect 113652 7274 113680 7754
rect 114848 7750 114876 7822
rect 114836 7744 114888 7750
rect 114836 7686 114888 7692
rect 114848 7410 114876 7686
rect 114836 7404 114888 7410
rect 114836 7346 114888 7352
rect 113640 7268 113692 7274
rect 113640 7210 113692 7216
rect 113364 7200 113416 7206
rect 113364 7142 113416 7148
rect 118516 7200 118568 7206
rect 118516 7142 118568 7148
rect 112812 6860 112864 6866
rect 112812 6802 112864 6808
rect 113376 6798 113404 7142
rect 112720 6792 112772 6798
rect 112720 6734 112772 6740
rect 113364 6792 113416 6798
rect 113364 6734 113416 6740
rect 114652 6792 114704 6798
rect 114652 6734 114704 6740
rect 110880 6724 110932 6730
rect 110880 6666 110932 6672
rect 110892 5846 110920 6666
rect 111524 6656 111576 6662
rect 111524 6598 111576 6604
rect 111536 5914 111564 6598
rect 111984 6316 112036 6322
rect 111984 6258 112036 6264
rect 111996 6118 112024 6258
rect 111984 6112 112036 6118
rect 111984 6054 112036 6060
rect 111524 5908 111576 5914
rect 111524 5850 111576 5856
rect 110880 5840 110932 5846
rect 110880 5782 110932 5788
rect 111064 3596 111116 3602
rect 111064 3538 111116 3544
rect 111076 3466 111104 3538
rect 111064 3460 111116 3466
rect 111064 3402 111116 3408
rect 111892 3392 111944 3398
rect 111892 3334 111944 3340
rect 111708 2848 111760 2854
rect 111708 2790 111760 2796
rect 110052 2644 110104 2650
rect 110052 2586 110104 2592
rect 110788 2644 110840 2650
rect 110788 2586 110840 2592
rect 110064 2514 110092 2586
rect 110052 2508 110104 2514
rect 110052 2450 110104 2456
rect 110328 2508 110380 2514
rect 110328 2450 110380 2456
rect 109776 2440 109828 2446
rect 109776 2382 109828 2388
rect 109224 2304 109276 2310
rect 109224 2246 109276 2252
rect 109236 1834 109264 2246
rect 109224 1828 109276 1834
rect 109224 1770 109276 1776
rect 110340 1426 110368 2450
rect 110800 2446 110828 2586
rect 111720 2582 111748 2790
rect 111708 2576 111760 2582
rect 111708 2518 111760 2524
rect 110788 2440 110840 2446
rect 110788 2382 110840 2388
rect 111904 2281 111932 3334
rect 111890 2272 111946 2281
rect 111890 2207 111946 2216
rect 111996 1698 112024 6054
rect 112628 4616 112680 4622
rect 112628 4558 112680 4564
rect 112352 2848 112404 2854
rect 112352 2790 112404 2796
rect 112364 2378 112392 2790
rect 112640 2650 112668 4558
rect 112732 3534 112760 6734
rect 114192 6724 114244 6730
rect 114192 6666 114244 6672
rect 114204 6633 114232 6666
rect 114190 6624 114246 6633
rect 114190 6559 114246 6568
rect 113192 6458 113404 6474
rect 113192 6452 113416 6458
rect 113192 6446 113364 6452
rect 113192 6322 113220 6446
rect 113364 6394 113416 6400
rect 113180 6316 113232 6322
rect 113180 6258 113232 6264
rect 113548 6316 113600 6322
rect 113548 6258 113600 6264
rect 113560 5574 113588 6258
rect 114100 6248 114152 6254
rect 114100 6190 114152 6196
rect 114112 5914 114140 6190
rect 114664 6118 114692 6734
rect 116032 6656 116084 6662
rect 116032 6598 116084 6604
rect 116676 6656 116728 6662
rect 116676 6598 116728 6604
rect 114652 6112 114704 6118
rect 114652 6054 114704 6060
rect 114100 5908 114152 5914
rect 114100 5850 114152 5856
rect 113548 5568 113600 5574
rect 113548 5510 113600 5516
rect 112720 3528 112772 3534
rect 112720 3470 112772 3476
rect 114560 3392 114612 3398
rect 114560 3334 114612 3340
rect 112996 2848 113048 2854
rect 112994 2816 112996 2825
rect 113048 2816 113050 2825
rect 112994 2751 113050 2760
rect 113178 2816 113234 2825
rect 113178 2751 113234 2760
rect 112628 2644 112680 2650
rect 112628 2586 112680 2592
rect 112352 2372 112404 2378
rect 112352 2314 112404 2320
rect 112364 2009 112392 2314
rect 112350 2000 112406 2009
rect 112350 1935 112406 1944
rect 111984 1692 112036 1698
rect 111984 1634 112036 1640
rect 112812 1692 112864 1698
rect 112812 1634 112864 1640
rect 110788 1624 110840 1630
rect 110788 1566 110840 1572
rect 110800 1426 110828 1566
rect 110328 1420 110380 1426
rect 110328 1362 110380 1368
rect 110788 1420 110840 1426
rect 110788 1362 110840 1368
rect 112824 1222 112852 1634
rect 113192 1358 113220 2751
rect 114572 1465 114600 3334
rect 114664 2854 114692 6054
rect 115388 5772 115440 5778
rect 115388 5714 115440 5720
rect 115112 5228 115164 5234
rect 115112 5170 115164 5176
rect 115124 3670 115152 5170
rect 115112 3664 115164 3670
rect 115112 3606 115164 3612
rect 114652 2848 114704 2854
rect 114652 2790 114704 2796
rect 115296 2848 115348 2854
rect 115296 2790 115348 2796
rect 115308 2378 115336 2790
rect 115296 2372 115348 2378
rect 115296 2314 115348 2320
rect 115204 2304 115256 2310
rect 115204 2246 115256 2252
rect 114928 1760 114980 1766
rect 114928 1702 114980 1708
rect 114558 1456 114614 1465
rect 114558 1391 114614 1400
rect 113180 1352 113232 1358
rect 113180 1294 113232 1300
rect 113640 1352 113692 1358
rect 113640 1294 113692 1300
rect 114742 1320 114798 1329
rect 110696 1216 110748 1222
rect 110696 1158 110748 1164
rect 110788 1216 110840 1222
rect 112812 1216 112864 1222
rect 110788 1158 110840 1164
rect 111890 1184 111946 1193
rect 110708 513 110736 1158
rect 110800 1086 110828 1158
rect 112812 1158 112864 1164
rect 113088 1216 113140 1222
rect 113088 1158 113140 1164
rect 111890 1119 111946 1128
rect 110788 1080 110840 1086
rect 110788 1022 110840 1028
rect 110880 1080 110932 1086
rect 110880 1022 110932 1028
rect 110892 814 110920 1022
rect 111904 814 111932 1119
rect 113100 814 113128 1158
rect 113652 1154 113680 1294
rect 114742 1255 114798 1264
rect 113824 1216 113876 1222
rect 113824 1158 113876 1164
rect 113640 1148 113692 1154
rect 113640 1090 113692 1096
rect 113836 1086 113864 1158
rect 113824 1080 113876 1086
rect 113824 1022 113876 1028
rect 113916 1080 113968 1086
rect 113916 1022 113968 1028
rect 114560 1080 114612 1086
rect 114560 1022 114612 1028
rect 113364 1012 113416 1018
rect 113364 954 113416 960
rect 110880 808 110932 814
rect 110880 750 110932 756
rect 111892 808 111944 814
rect 111892 750 111944 756
rect 113088 808 113140 814
rect 113088 750 113140 756
rect 113376 610 113404 954
rect 113928 950 113956 1022
rect 113916 944 113968 950
rect 113916 886 113968 892
rect 114008 944 114060 950
rect 114008 886 114060 892
rect 114020 678 114048 886
rect 114008 672 114060 678
rect 114008 614 114060 620
rect 113364 604 113416 610
rect 113364 546 113416 552
rect 114192 604 114244 610
rect 114468 604 114520 610
rect 114244 564 114468 592
rect 114192 546 114244 552
rect 114468 546 114520 552
rect 89220 504 89222 513
rect 89166 439 89222 448
rect 94686 504 94742 513
rect 94686 439 94742 448
rect 97906 504 97962 513
rect 97906 439 97908 448
rect 97960 439 97962 448
rect 103610 504 103666 513
rect 103610 439 103666 448
rect 108854 504 108910 513
rect 108854 439 108910 448
rect 109130 504 109186 513
rect 109130 439 109186 448
rect 110694 504 110750 513
rect 110694 439 110750 448
rect 97908 410 97960 416
rect 114572 270 114600 1022
rect 114756 746 114784 1255
rect 114744 740 114796 746
rect 114744 682 114796 688
rect 114940 542 114968 1702
rect 115216 1630 115244 2246
rect 115308 1902 115336 2314
rect 115296 1896 115348 1902
rect 115296 1838 115348 1844
rect 115204 1624 115256 1630
rect 115204 1566 115256 1572
rect 115020 1216 115072 1222
rect 115112 1216 115164 1222
rect 115020 1158 115072 1164
rect 115110 1184 115112 1193
rect 115164 1184 115166 1193
rect 115032 1086 115060 1158
rect 115110 1119 115166 1128
rect 115204 1148 115256 1154
rect 115204 1090 115256 1096
rect 115020 1080 115072 1086
rect 115020 1022 115072 1028
rect 115216 1018 115244 1090
rect 115204 1012 115256 1018
rect 115204 954 115256 960
rect 115400 678 115428 5714
rect 115480 5568 115532 5574
rect 115480 5510 115532 5516
rect 115492 1970 115520 5510
rect 115480 1964 115532 1970
rect 115480 1906 115532 1912
rect 115388 672 115440 678
rect 115388 614 115440 620
rect 114928 536 114980 542
rect 114742 504 114798 513
rect 116044 513 116072 6598
rect 116688 3058 116716 6598
rect 117504 6316 117556 6322
rect 117504 6258 117556 6264
rect 117516 6118 117544 6258
rect 118528 6254 118556 7142
rect 118792 6860 118844 6866
rect 118792 6802 118844 6808
rect 117964 6248 118016 6254
rect 117964 6190 118016 6196
rect 118516 6248 118568 6254
rect 118516 6190 118568 6196
rect 117504 6112 117556 6118
rect 117504 6054 117556 6060
rect 117136 5704 117188 5710
rect 117136 5646 117188 5652
rect 117148 5166 117176 5646
rect 117136 5160 117188 5166
rect 117136 5102 117188 5108
rect 117516 3534 117544 6054
rect 117504 3528 117556 3534
rect 117504 3470 117556 3476
rect 117596 3460 117648 3466
rect 117596 3402 117648 3408
rect 117608 3058 117636 3402
rect 116676 3052 116728 3058
rect 116676 2994 116728 3000
rect 117596 3052 117648 3058
rect 117596 2994 117648 3000
rect 117608 2774 117636 2994
rect 117516 2746 117636 2774
rect 116492 1012 116544 1018
rect 116492 954 116544 960
rect 116504 814 116532 954
rect 116492 808 116544 814
rect 116492 750 116544 756
rect 114928 478 114980 484
rect 116030 504 116086 513
rect 114742 439 114744 448
rect 114796 439 114798 448
rect 117516 474 117544 2746
rect 117976 1329 118004 6190
rect 118804 5710 118832 6802
rect 120448 6656 120500 6662
rect 120448 6598 120500 6604
rect 120460 6322 120488 6598
rect 121012 6322 121040 7890
rect 122576 7886 122604 8026
rect 122564 7880 122616 7886
rect 122564 7822 122616 7828
rect 121644 6656 121696 6662
rect 121644 6598 121696 6604
rect 122104 6656 122156 6662
rect 122104 6598 122156 6604
rect 121656 6322 121684 6598
rect 122116 6458 122144 6598
rect 122104 6452 122156 6458
rect 122104 6394 122156 6400
rect 120448 6316 120500 6322
rect 120448 6258 120500 6264
rect 121000 6316 121052 6322
rect 121000 6258 121052 6264
rect 121644 6316 121696 6322
rect 121644 6258 121696 6264
rect 120172 5840 120224 5846
rect 120172 5782 120224 5788
rect 118792 5704 118844 5710
rect 118792 5646 118844 5652
rect 118884 5568 118936 5574
rect 118884 5510 118936 5516
rect 118606 2000 118662 2009
rect 118606 1935 118662 1944
rect 117962 1320 118018 1329
rect 117962 1255 118018 1264
rect 118514 1184 118570 1193
rect 118514 1119 118570 1128
rect 118528 678 118556 1119
rect 118620 1086 118648 1935
rect 118700 1760 118752 1766
rect 118700 1702 118752 1708
rect 118712 1562 118740 1702
rect 118700 1556 118752 1562
rect 118700 1498 118752 1504
rect 118792 1556 118844 1562
rect 118792 1498 118844 1504
rect 118804 1306 118832 1498
rect 118896 1494 118924 5510
rect 119344 3392 119396 3398
rect 119344 3334 119396 3340
rect 119356 2825 119384 3334
rect 120080 2848 120132 2854
rect 119342 2816 119398 2825
rect 120080 2790 120132 2796
rect 119342 2751 119398 2760
rect 119436 2440 119488 2446
rect 119436 2382 119488 2388
rect 118884 1488 118936 1494
rect 118884 1430 118936 1436
rect 118712 1290 118832 1306
rect 118700 1284 118832 1290
rect 118752 1278 118832 1284
rect 118700 1226 118752 1232
rect 118790 1184 118846 1193
rect 118790 1119 118846 1128
rect 118804 1086 118832 1119
rect 118608 1080 118660 1086
rect 118608 1022 118660 1028
rect 118792 1080 118844 1086
rect 118792 1022 118844 1028
rect 118516 672 118568 678
rect 118516 614 118568 620
rect 118608 672 118660 678
rect 118608 614 118660 620
rect 118620 542 118648 614
rect 118608 536 118660 542
rect 118608 478 118660 484
rect 116030 439 116086 448
rect 117504 468 117556 474
rect 114744 410 114796 416
rect 117504 410 117556 416
rect 119448 270 119476 2382
rect 120092 2378 120120 2790
rect 120080 2372 120132 2378
rect 120080 2314 120132 2320
rect 119620 1488 119672 1494
rect 119526 1456 119582 1465
rect 119620 1430 119672 1436
rect 119526 1391 119582 1400
rect 119540 678 119568 1391
rect 119632 882 119660 1430
rect 119620 876 119672 882
rect 119620 818 119672 824
rect 119528 672 119580 678
rect 120092 626 120120 2314
rect 120184 1193 120212 5782
rect 120460 3738 120488 6258
rect 120724 5704 120776 5710
rect 120724 5646 120776 5652
rect 120736 5030 120764 5646
rect 120724 5024 120776 5030
rect 120724 4966 120776 4972
rect 121656 3942 121684 6258
rect 123128 6186 123156 11154
rect 145748 10396 145800 10402
rect 145748 10338 145800 10344
rect 127808 9716 127860 9722
rect 127808 9658 127860 9664
rect 123392 9648 123444 9654
rect 123392 9590 123444 9596
rect 123300 8084 123352 8090
rect 123300 8026 123352 8032
rect 123116 6180 123168 6186
rect 123116 6122 123168 6128
rect 123208 6112 123260 6118
rect 123208 6054 123260 6060
rect 122840 5704 122892 5710
rect 122840 5646 122892 5652
rect 122852 5030 122880 5646
rect 122840 5024 122892 5030
rect 122840 4966 122892 4972
rect 122852 4826 122880 4966
rect 122840 4820 122892 4826
rect 122840 4762 122892 4768
rect 123220 4010 123248 6054
rect 123312 5914 123340 8026
rect 123404 6662 123432 9590
rect 126336 7812 126388 7818
rect 126336 7754 126388 7760
rect 126348 7546 126376 7754
rect 127716 7744 127768 7750
rect 127716 7686 127768 7692
rect 127728 7546 127756 7686
rect 126336 7540 126388 7546
rect 126336 7482 126388 7488
rect 127716 7540 127768 7546
rect 127716 7482 127768 7488
rect 123484 7268 123536 7274
rect 123484 7210 123536 7216
rect 123392 6656 123444 6662
rect 123392 6598 123444 6604
rect 123496 6322 123524 7210
rect 125140 6928 125192 6934
rect 125140 6870 125192 6876
rect 124036 6656 124088 6662
rect 124036 6598 124088 6604
rect 123484 6316 123536 6322
rect 123484 6258 123536 6264
rect 123300 5908 123352 5914
rect 123300 5850 123352 5856
rect 124048 5710 124076 6598
rect 125152 6322 125180 6870
rect 125506 6352 125562 6361
rect 125140 6316 125192 6322
rect 127820 6322 127848 9658
rect 135260 8628 135312 8634
rect 135260 8570 135312 8576
rect 135272 8022 135300 8570
rect 145760 8566 145788 10338
rect 145840 10328 145892 10334
rect 145840 10270 145892 10276
rect 149704 10328 149756 10334
rect 149704 10270 149756 10276
rect 145852 8566 145880 10270
rect 145748 8560 145800 8566
rect 145748 8502 145800 8508
rect 145840 8560 145892 8566
rect 145840 8502 145892 8508
rect 149716 8498 149744 10270
rect 157904 8498 157932 11494
rect 173072 10192 173124 10198
rect 173072 10134 173124 10140
rect 171784 9580 171836 9586
rect 171784 9522 171836 9528
rect 167368 9512 167420 9518
rect 167104 9460 167368 9466
rect 167104 9454 167420 9460
rect 167104 9450 167408 9454
rect 167092 9444 167408 9450
rect 167144 9438 167408 9444
rect 167092 9386 167144 9392
rect 168748 9036 168800 9042
rect 168748 8978 168800 8984
rect 160100 8900 160152 8906
rect 160100 8842 160152 8848
rect 167552 8900 167604 8906
rect 167552 8842 167604 8848
rect 149704 8492 149756 8498
rect 149704 8434 149756 8440
rect 157892 8492 157944 8498
rect 157892 8434 157944 8440
rect 149060 8424 149112 8430
rect 149060 8366 149112 8372
rect 135260 8016 135312 8022
rect 135260 7958 135312 7964
rect 139032 8016 139084 8022
rect 139032 7958 139084 7964
rect 132040 7880 132092 7886
rect 132040 7822 132092 7828
rect 131396 7812 131448 7818
rect 131396 7754 131448 7760
rect 131408 7478 131436 7754
rect 131396 7472 131448 7478
rect 131396 7414 131448 7420
rect 131396 6452 131448 6458
rect 131396 6394 131448 6400
rect 128188 6322 128400 6338
rect 131408 6322 131436 6394
rect 125506 6287 125508 6296
rect 125140 6258 125192 6264
rect 125560 6287 125562 6296
rect 126612 6316 126664 6322
rect 125508 6258 125560 6264
rect 126612 6258 126664 6264
rect 127808 6316 127860 6322
rect 127808 6258 127860 6264
rect 128188 6316 128412 6322
rect 128188 6310 128360 6316
rect 124680 6180 124732 6186
rect 124680 6122 124732 6128
rect 124692 5778 124720 6122
rect 124680 5772 124732 5778
rect 124680 5714 124732 5720
rect 124036 5704 124088 5710
rect 124036 5646 124088 5652
rect 124128 5704 124180 5710
rect 124128 5646 124180 5652
rect 124140 5098 124168 5646
rect 124128 5092 124180 5098
rect 124128 5034 124180 5040
rect 123392 4820 123444 4826
rect 123392 4762 123444 4768
rect 123404 4554 123432 4762
rect 123392 4548 123444 4554
rect 123392 4490 123444 4496
rect 125152 4078 125180 6258
rect 126624 6118 126652 6258
rect 126612 6112 126664 6118
rect 126612 6054 126664 6060
rect 125692 5228 125744 5234
rect 125692 5170 125744 5176
rect 125704 5030 125732 5170
rect 125692 5024 125744 5030
rect 125692 4966 125744 4972
rect 125704 4729 125732 4966
rect 125690 4720 125746 4729
rect 125690 4655 125746 4664
rect 126624 4146 126652 6054
rect 127348 5908 127400 5914
rect 127348 5850 127400 5856
rect 127360 5710 127388 5850
rect 127348 5704 127400 5710
rect 127348 5646 127400 5652
rect 128188 5574 128216 6310
rect 128360 6258 128412 6264
rect 131396 6316 131448 6322
rect 131396 6258 131448 6264
rect 130934 6216 130990 6225
rect 130934 6151 130990 6160
rect 130948 5710 130976 6151
rect 131764 6112 131816 6118
rect 131764 6054 131816 6060
rect 131776 5710 131804 6054
rect 132052 5710 132080 7822
rect 136640 7812 136692 7818
rect 136640 7754 136692 7760
rect 132868 7744 132920 7750
rect 132868 7686 132920 7692
rect 130660 5704 130712 5710
rect 130660 5646 130712 5652
rect 130936 5704 130988 5710
rect 130936 5646 130988 5652
rect 131764 5704 131816 5710
rect 131764 5646 131816 5652
rect 132040 5704 132092 5710
rect 132040 5646 132092 5652
rect 130672 5574 130700 5646
rect 128176 5568 128228 5574
rect 128176 5510 128228 5516
rect 130108 5568 130160 5574
rect 130108 5510 130160 5516
rect 130660 5568 130712 5574
rect 130660 5510 130712 5516
rect 127624 5228 127676 5234
rect 127624 5170 127676 5176
rect 127636 4486 127664 5170
rect 128084 5160 128136 5166
rect 128084 5102 128136 5108
rect 127624 4480 127676 4486
rect 127624 4422 127676 4428
rect 127716 4480 127768 4486
rect 127716 4422 127768 4428
rect 126612 4140 126664 4146
rect 126612 4082 126664 4088
rect 126888 4140 126940 4146
rect 126888 4082 126940 4088
rect 125140 4072 125192 4078
rect 125140 4014 125192 4020
rect 123208 4004 123260 4010
rect 123208 3946 123260 3952
rect 121644 3936 121696 3942
rect 121644 3878 121696 3884
rect 122932 3936 122984 3942
rect 122932 3878 122984 3884
rect 122944 3738 122972 3878
rect 120448 3732 120500 3738
rect 120448 3674 120500 3680
rect 122932 3732 122984 3738
rect 122932 3674 122984 3680
rect 122656 3460 122708 3466
rect 122656 3402 122708 3408
rect 121092 3392 121144 3398
rect 121092 3334 121144 3340
rect 121104 2825 121132 3334
rect 122668 2854 122696 3402
rect 124220 3392 124272 3398
rect 124220 3334 124272 3340
rect 125692 3392 125744 3398
rect 125692 3334 125744 3340
rect 121460 2848 121512 2854
rect 121090 2816 121146 2825
rect 121460 2790 121512 2796
rect 122656 2848 122708 2854
rect 122656 2790 122708 2796
rect 121090 2751 121146 2760
rect 120356 2304 120408 2310
rect 120356 2246 120408 2252
rect 120368 1902 120396 2246
rect 120356 1896 120408 1902
rect 120356 1838 120408 1844
rect 121472 1698 121500 2790
rect 122932 2304 122984 2310
rect 122932 2246 122984 2252
rect 122944 1970 122972 2246
rect 122932 1964 122984 1970
rect 122932 1906 122984 1912
rect 121460 1692 121512 1698
rect 121460 1634 121512 1640
rect 121736 1692 121788 1698
rect 121736 1634 121788 1640
rect 120170 1184 120226 1193
rect 121748 1154 121776 1634
rect 124232 1562 124260 3334
rect 125508 2304 125560 2310
rect 125508 2246 125560 2252
rect 124494 2000 124550 2009
rect 124494 1935 124550 1944
rect 124220 1556 124272 1562
rect 124220 1498 124272 1504
rect 123576 1216 123628 1222
rect 123576 1158 123628 1164
rect 120170 1119 120226 1128
rect 121736 1148 121788 1154
rect 121736 1090 121788 1096
rect 122104 1148 122156 1154
rect 122104 1090 122156 1096
rect 122116 814 122144 1090
rect 123588 882 123616 1158
rect 123576 876 123628 882
rect 123576 818 123628 824
rect 122104 808 122156 814
rect 122104 750 122156 756
rect 119528 614 119580 620
rect 119724 610 120120 626
rect 119712 604 120120 610
rect 119764 598 120120 604
rect 119712 546 119764 552
rect 124508 270 124536 1935
rect 125520 1834 125548 2246
rect 125508 1828 125560 1834
rect 125508 1770 125560 1776
rect 125704 1494 125732 3334
rect 126900 2650 126928 4082
rect 126888 2644 126940 2650
rect 126888 2586 126940 2592
rect 126428 2508 126480 2514
rect 126428 2450 126480 2456
rect 126244 2304 126296 2310
rect 126244 2246 126296 2252
rect 126256 2009 126284 2246
rect 126242 2000 126298 2009
rect 126242 1935 126298 1944
rect 125692 1488 125744 1494
rect 125692 1430 125744 1436
rect 126152 1488 126204 1494
rect 126152 1430 126204 1436
rect 126164 1222 126192 1430
rect 126152 1216 126204 1222
rect 126152 1158 126204 1164
rect 126244 1216 126296 1222
rect 126244 1158 126296 1164
rect 126256 814 126284 1158
rect 126244 808 126296 814
rect 126244 750 126296 756
rect 126440 270 126468 2450
rect 127072 2372 127124 2378
rect 127072 2314 127124 2320
rect 126980 1488 127032 1494
rect 127084 1465 127112 2314
rect 127636 1766 127664 4422
rect 127728 2106 127756 4422
rect 128096 4214 128124 5102
rect 128188 4826 128216 5510
rect 129556 5024 129608 5030
rect 129556 4966 129608 4972
rect 128176 4820 128228 4826
rect 128176 4762 128228 4768
rect 129568 4690 129596 4966
rect 129556 4684 129608 4690
rect 129556 4626 129608 4632
rect 128084 4208 128136 4214
rect 128084 4150 128136 4156
rect 128360 3392 128412 3398
rect 128360 3334 128412 3340
rect 128372 3058 128400 3334
rect 128360 3052 128412 3058
rect 128360 2994 128412 3000
rect 130120 2922 130148 5510
rect 131212 5228 131264 5234
rect 131212 5170 131264 5176
rect 130844 5160 130896 5166
rect 130844 5102 130896 5108
rect 130856 4826 130884 5102
rect 130844 4820 130896 4826
rect 130844 4762 130896 4768
rect 130384 4684 130436 4690
rect 130384 4626 130436 4632
rect 130396 4554 130424 4626
rect 130844 4616 130896 4622
rect 131028 4616 131080 4622
rect 130896 4564 131028 4570
rect 131224 4593 131252 5170
rect 130844 4558 131080 4564
rect 131210 4584 131266 4593
rect 130384 4548 130436 4554
rect 130856 4542 131068 4558
rect 131210 4519 131212 4528
rect 130384 4490 130436 4496
rect 131264 4519 131266 4528
rect 131212 4490 131264 4496
rect 130844 4004 130896 4010
rect 130844 3946 130896 3952
rect 130856 3738 130884 3946
rect 130844 3732 130896 3738
rect 130844 3674 130896 3680
rect 130476 3528 130528 3534
rect 130476 3470 130528 3476
rect 130108 2916 130160 2922
rect 130108 2858 130160 2864
rect 128176 2848 128228 2854
rect 128176 2790 128228 2796
rect 128188 2378 128216 2790
rect 130488 2514 130516 3470
rect 131776 3194 131804 5646
rect 132684 5228 132736 5234
rect 132684 5170 132736 5176
rect 132696 5030 132724 5170
rect 132684 5024 132736 5030
rect 132684 4966 132736 4972
rect 132696 4758 132724 4966
rect 132684 4752 132736 4758
rect 132684 4694 132736 4700
rect 132500 3528 132552 3534
rect 132500 3470 132552 3476
rect 131764 3188 131816 3194
rect 131764 3130 131816 3136
rect 130476 2508 130528 2514
rect 130476 2450 130528 2456
rect 128268 2440 128320 2446
rect 128268 2382 128320 2388
rect 130660 2440 130712 2446
rect 130660 2382 130712 2388
rect 128176 2372 128228 2378
rect 128176 2314 128228 2320
rect 128084 2304 128136 2310
rect 128084 2246 128136 2252
rect 127716 2100 127768 2106
rect 127716 2042 127768 2048
rect 127992 2100 128044 2106
rect 127992 2042 128044 2048
rect 127624 1760 127676 1766
rect 127624 1702 127676 1708
rect 126980 1430 127032 1436
rect 127070 1456 127126 1465
rect 126992 1290 127020 1430
rect 127070 1391 127126 1400
rect 126888 1284 126940 1290
rect 126888 1226 126940 1232
rect 126980 1284 127032 1290
rect 126980 1226 127032 1232
rect 126900 678 126928 1226
rect 128004 882 128032 2042
rect 128096 1494 128124 2246
rect 128176 1760 128228 1766
rect 128176 1702 128228 1708
rect 128084 1488 128136 1494
rect 128084 1430 128136 1436
rect 127992 876 128044 882
rect 127992 818 128044 824
rect 128188 814 128216 1702
rect 128280 950 128308 2382
rect 128360 2372 128412 2378
rect 128360 2314 128412 2320
rect 128268 944 128320 950
rect 128268 886 128320 892
rect 128176 808 128228 814
rect 128176 750 128228 756
rect 128372 678 128400 2314
rect 130672 2038 130700 2382
rect 130844 2304 130896 2310
rect 130844 2246 130896 2252
rect 130660 2032 130712 2038
rect 130660 1974 130712 1980
rect 130856 1834 130884 2246
rect 130844 1828 130896 1834
rect 130844 1770 130896 1776
rect 132512 1698 132540 3470
rect 132880 3194 132908 7686
rect 134432 6112 134484 6118
rect 134432 6054 134484 6060
rect 135534 6080 135590 6089
rect 134444 5710 134472 6054
rect 135534 6015 135590 6024
rect 135548 5778 135576 6015
rect 135536 5772 135588 5778
rect 135536 5714 135588 5720
rect 134432 5704 134484 5710
rect 134432 5646 134484 5652
rect 135352 5704 135404 5710
rect 135352 5646 135404 5652
rect 133604 5568 133656 5574
rect 133604 5510 133656 5516
rect 133512 5160 133564 5166
rect 133512 5102 133564 5108
rect 133524 4729 133552 5102
rect 133510 4720 133566 4729
rect 133510 4655 133566 4664
rect 133052 4072 133104 4078
rect 133052 4014 133104 4020
rect 133064 3602 133092 4014
rect 133144 3936 133196 3942
rect 133144 3878 133196 3884
rect 133156 3738 133184 3878
rect 133144 3732 133196 3738
rect 133144 3674 133196 3680
rect 133052 3596 133104 3602
rect 133052 3538 133104 3544
rect 132868 3188 132920 3194
rect 132868 3130 132920 3136
rect 133616 3126 133644 5510
rect 134340 5228 134392 5234
rect 134340 5170 134392 5176
rect 134352 4486 134380 5170
rect 135364 5030 135392 5646
rect 135352 5024 135404 5030
rect 135352 4966 135404 4972
rect 135364 4758 135392 4966
rect 135352 4752 135404 4758
rect 135352 4694 135404 4700
rect 134340 4480 134392 4486
rect 134340 4422 134392 4428
rect 136180 4480 136232 4486
rect 136180 4422 136232 4428
rect 134340 3664 134392 3670
rect 134340 3606 134392 3612
rect 135260 3664 135312 3670
rect 135260 3606 135312 3612
rect 133604 3120 133656 3126
rect 133604 3062 133656 3068
rect 134352 3058 134380 3606
rect 134340 3052 134392 3058
rect 134340 2994 134392 3000
rect 133972 2304 134024 2310
rect 133972 2246 134024 2252
rect 132592 1760 132644 1766
rect 132592 1702 132644 1708
rect 132500 1692 132552 1698
rect 132500 1634 132552 1640
rect 132224 1488 132276 1494
rect 130474 1456 130530 1465
rect 132500 1488 132552 1494
rect 132276 1448 132500 1476
rect 132224 1430 132276 1436
rect 132500 1430 132552 1436
rect 132604 1426 132632 1702
rect 133984 1698 134012 2246
rect 133972 1692 134024 1698
rect 133972 1634 134024 1640
rect 135272 1465 135300 3606
rect 136088 3460 136140 3466
rect 136088 3402 136140 3408
rect 136100 3126 136128 3402
rect 136088 3120 136140 3126
rect 136088 3062 136140 3068
rect 136192 1562 136220 4422
rect 136652 2417 136680 7754
rect 138296 5704 138348 5710
rect 138216 5652 138296 5658
rect 138216 5646 138348 5652
rect 138216 5630 138336 5646
rect 139044 5642 139072 7958
rect 141240 7880 141292 7886
rect 141240 7822 141292 7828
rect 141252 7478 141280 7822
rect 141240 7472 141292 7478
rect 141240 7414 141292 7420
rect 139032 5636 139084 5642
rect 138216 5574 138244 5630
rect 139032 5578 139084 5584
rect 138204 5568 138256 5574
rect 138204 5510 138256 5516
rect 141700 5568 141752 5574
rect 141700 5510 141752 5516
rect 137008 5296 137060 5302
rect 137008 5238 137060 5244
rect 137020 5030 137048 5238
rect 137100 5228 137152 5234
rect 137100 5170 137152 5176
rect 137112 5030 137140 5170
rect 137836 5160 137888 5166
rect 137836 5102 137888 5108
rect 137008 5024 137060 5030
rect 137008 4966 137060 4972
rect 137100 5024 137152 5030
rect 137100 4966 137152 4972
rect 137020 2990 137048 4966
rect 137848 4457 137876 5102
rect 138112 4820 138164 4826
rect 138112 4762 138164 4768
rect 138124 4690 138152 4762
rect 138112 4684 138164 4690
rect 138112 4626 138164 4632
rect 137928 4616 137980 4622
rect 137928 4558 137980 4564
rect 137834 4448 137890 4457
rect 137834 4383 137890 4392
rect 137940 4146 137968 4558
rect 138216 4282 138244 5510
rect 141330 5400 141386 5409
rect 141330 5335 141386 5344
rect 141344 5234 141372 5335
rect 141712 5234 141740 5510
rect 145840 5296 145892 5302
rect 145840 5238 145892 5244
rect 140504 5228 140556 5234
rect 140504 5170 140556 5176
rect 141332 5228 141384 5234
rect 141332 5170 141384 5176
rect 141700 5228 141752 5234
rect 141700 5170 141752 5176
rect 144552 5228 144604 5234
rect 144552 5170 144604 5176
rect 145472 5228 145524 5234
rect 145472 5170 145524 5176
rect 140516 5030 140544 5170
rect 140504 5024 140556 5030
rect 140504 4966 140556 4972
rect 140688 5024 140740 5030
rect 140688 4966 140740 4972
rect 138204 4276 138256 4282
rect 138204 4218 138256 4224
rect 137928 4140 137980 4146
rect 137928 4082 137980 4088
rect 140700 3738 140728 4966
rect 141608 4752 141660 4758
rect 141608 4694 141660 4700
rect 141056 4616 141108 4622
rect 141056 4558 141108 4564
rect 141068 3942 141096 4558
rect 141620 4554 141648 4694
rect 141608 4548 141660 4554
rect 141608 4490 141660 4496
rect 141712 4146 141740 5170
rect 142436 5160 142488 5166
rect 142436 5102 142488 5108
rect 142448 4282 142476 5102
rect 144564 5030 144592 5170
rect 144828 5160 144880 5166
rect 144828 5102 144880 5108
rect 144552 5024 144604 5030
rect 144552 4966 144604 4972
rect 144644 5024 144696 5030
rect 144644 4966 144696 4972
rect 142436 4276 142488 4282
rect 142436 4218 142488 4224
rect 141700 4140 141752 4146
rect 141700 4082 141752 4088
rect 144000 4072 144052 4078
rect 144000 4014 144052 4020
rect 143172 4004 143224 4010
rect 143172 3946 143224 3952
rect 140964 3936 141016 3942
rect 140964 3878 141016 3884
rect 141056 3936 141108 3942
rect 141056 3878 141108 3884
rect 141700 3936 141752 3942
rect 141700 3878 141752 3884
rect 140976 3738 141004 3878
rect 140688 3732 140740 3738
rect 140688 3674 140740 3680
rect 140964 3732 141016 3738
rect 140964 3674 141016 3680
rect 137008 2984 137060 2990
rect 137008 2926 137060 2932
rect 138020 2848 138072 2854
rect 138020 2790 138072 2796
rect 138032 2530 138060 2790
rect 138032 2502 138152 2530
rect 138124 2446 138152 2502
rect 138112 2440 138164 2446
rect 136638 2408 136694 2417
rect 138112 2382 138164 2388
rect 136638 2343 136694 2352
rect 136456 2304 136508 2310
rect 136456 2246 136508 2252
rect 136468 2106 136496 2246
rect 136456 2100 136508 2106
rect 136456 2042 136508 2048
rect 138124 1630 138152 2382
rect 139124 2032 139176 2038
rect 139124 1974 139176 1980
rect 137008 1624 137060 1630
rect 137008 1566 137060 1572
rect 138112 1624 138164 1630
rect 138112 1566 138164 1572
rect 136180 1556 136232 1562
rect 136180 1498 136232 1504
rect 135258 1456 135314 1465
rect 130474 1391 130530 1400
rect 132592 1420 132644 1426
rect 130488 882 130516 1391
rect 135258 1391 135314 1400
rect 132592 1362 132644 1368
rect 133144 1284 133196 1290
rect 133144 1226 133196 1232
rect 133236 1284 133288 1290
rect 133236 1226 133288 1232
rect 130752 1148 130804 1154
rect 130752 1090 130804 1096
rect 132960 1148 133012 1154
rect 132960 1090 133012 1096
rect 130764 1034 130792 1090
rect 130764 1006 131068 1034
rect 131040 950 131068 1006
rect 131028 944 131080 950
rect 131028 886 131080 892
rect 130476 876 130528 882
rect 130476 818 130528 824
rect 132972 814 133000 1090
rect 133156 1018 133184 1226
rect 133052 1012 133104 1018
rect 133052 954 133104 960
rect 133144 1012 133196 1018
rect 133144 954 133196 960
rect 133064 898 133092 954
rect 133248 898 133276 1226
rect 134892 1012 134944 1018
rect 134892 954 134944 960
rect 133064 870 133276 898
rect 134904 814 134932 954
rect 137020 882 137048 1566
rect 137744 1216 137796 1222
rect 137796 1164 137876 1170
rect 137744 1158 137876 1164
rect 137756 1142 137876 1158
rect 137848 882 137876 1142
rect 139136 882 139164 1974
rect 141068 1766 141096 3878
rect 141148 2644 141200 2650
rect 141148 2586 141200 2592
rect 141160 2446 141188 2586
rect 141148 2440 141200 2446
rect 141148 2382 141200 2388
rect 141712 1970 141740 3878
rect 143080 2848 143132 2854
rect 143080 2790 143132 2796
rect 143092 2446 143120 2790
rect 143080 2440 143132 2446
rect 143080 2382 143132 2388
rect 143092 2038 143120 2382
rect 143080 2032 143132 2038
rect 143080 1974 143132 1980
rect 141700 1964 141752 1970
rect 141700 1906 141752 1912
rect 143184 1902 143212 3946
rect 144012 2990 144040 4014
rect 144656 3738 144684 4966
rect 144840 4321 144868 5102
rect 145484 4486 145512 5170
rect 145852 4690 145880 5238
rect 145932 5228 145984 5234
rect 145932 5170 145984 5176
rect 148048 5228 148100 5234
rect 148048 5170 148100 5176
rect 145840 4684 145892 4690
rect 145840 4626 145892 4632
rect 145944 4593 145972 5170
rect 148060 5030 148088 5170
rect 148968 5160 149020 5166
rect 148968 5102 149020 5108
rect 148048 5024 148100 5030
rect 148048 4966 148100 4972
rect 145930 4584 145986 4593
rect 145930 4519 145986 4528
rect 145472 4480 145524 4486
rect 145472 4422 145524 4428
rect 144826 4312 144882 4321
rect 144826 4247 144882 4256
rect 144736 4004 144788 4010
rect 144736 3946 144788 3952
rect 144644 3732 144696 3738
rect 144644 3674 144696 3680
rect 144000 2984 144052 2990
rect 144000 2926 144052 2932
rect 143448 2372 143500 2378
rect 143448 2314 143500 2320
rect 143460 2106 143488 2314
rect 143448 2100 143500 2106
rect 143448 2042 143500 2048
rect 143172 1896 143224 1902
rect 143172 1838 143224 1844
rect 141056 1760 141108 1766
rect 141056 1702 141108 1708
rect 144748 1630 144776 3946
rect 145484 3602 145512 4422
rect 148140 4140 148192 4146
rect 148140 4082 148192 4088
rect 148152 3602 148180 4082
rect 148692 4072 148744 4078
rect 148692 4014 148744 4020
rect 148704 3738 148732 4014
rect 148692 3732 148744 3738
rect 148692 3674 148744 3680
rect 145472 3596 145524 3602
rect 145472 3538 145524 3544
rect 148140 3596 148192 3602
rect 148140 3538 148192 3544
rect 146850 2408 146906 2417
rect 146850 2343 146852 2352
rect 146904 2343 146906 2352
rect 146852 2314 146904 2320
rect 144920 2304 144972 2310
rect 144920 2246 144972 2252
rect 146668 2304 146720 2310
rect 146668 2246 146720 2252
rect 144736 1624 144788 1630
rect 144736 1566 144788 1572
rect 141424 1556 141476 1562
rect 141424 1498 141476 1504
rect 141436 1290 141464 1498
rect 143724 1488 143776 1494
rect 143724 1430 143776 1436
rect 141424 1284 141476 1290
rect 141424 1226 141476 1232
rect 141516 1284 141568 1290
rect 141516 1226 141568 1232
rect 139308 1216 139360 1222
rect 139308 1158 139360 1164
rect 139216 1148 139268 1154
rect 139216 1090 139268 1096
rect 139228 882 139256 1090
rect 139320 1018 139348 1158
rect 139400 1148 139452 1154
rect 139400 1090 139452 1096
rect 139308 1012 139360 1018
rect 139308 954 139360 960
rect 137008 876 137060 882
rect 137008 818 137060 824
rect 137836 876 137888 882
rect 137836 818 137888 824
rect 139124 876 139176 882
rect 139124 818 139176 824
rect 139216 876 139268 882
rect 139216 818 139268 824
rect 132960 808 133012 814
rect 132960 750 133012 756
rect 134892 808 134944 814
rect 134892 750 134944 756
rect 139412 746 139440 1090
rect 139492 944 139544 950
rect 139492 886 139544 892
rect 139400 740 139452 746
rect 139400 682 139452 688
rect 126888 672 126940 678
rect 126888 614 126940 620
rect 128360 672 128412 678
rect 139504 626 139532 886
rect 141528 814 141556 1226
rect 142712 1080 142764 1086
rect 142764 1028 142936 1034
rect 142712 1022 142936 1028
rect 142724 1018 142936 1022
rect 142724 1012 142948 1018
rect 142724 1006 142896 1012
rect 142896 954 142948 960
rect 143736 882 143764 1430
rect 144932 1426 144960 2246
rect 145840 1760 145892 1766
rect 145840 1702 145892 1708
rect 144920 1420 144972 1426
rect 144920 1362 144972 1368
rect 143724 876 143776 882
rect 143724 818 143776 824
rect 141516 808 141568 814
rect 141516 750 141568 756
rect 145852 678 145880 1702
rect 146208 1624 146260 1630
rect 146208 1566 146260 1572
rect 146220 950 146248 1566
rect 146390 1456 146446 1465
rect 146680 1426 146708 2246
rect 148152 1834 148180 3538
rect 148232 2848 148284 2854
rect 148232 2790 148284 2796
rect 148244 2446 148272 2790
rect 148232 2440 148284 2446
rect 148232 2382 148284 2388
rect 148140 1828 148192 1834
rect 148140 1770 148192 1776
rect 148244 1562 148272 2382
rect 148600 2372 148652 2378
rect 148600 2314 148652 2320
rect 148508 1760 148560 1766
rect 148508 1702 148560 1708
rect 148520 1630 148548 1702
rect 148612 1630 148640 2314
rect 148980 1902 149008 5102
rect 149072 2553 149100 8366
rect 149716 7886 149744 8434
rect 156696 8424 156748 8430
rect 156696 8366 156748 8372
rect 149704 7880 149756 7886
rect 149704 7822 149756 7828
rect 149704 5908 149756 5914
rect 149704 5850 149756 5856
rect 149716 5778 149744 5850
rect 149704 5772 149756 5778
rect 149704 5714 149756 5720
rect 149152 4616 149204 4622
rect 149152 4558 149204 4564
rect 149164 3058 149192 4558
rect 150808 4140 150860 4146
rect 150808 4082 150860 4088
rect 149152 3052 149204 3058
rect 149152 2994 149204 3000
rect 149058 2544 149114 2553
rect 150820 2514 150848 4082
rect 150900 4072 150952 4078
rect 150952 4020 151216 4026
rect 150900 4014 151216 4020
rect 150912 4010 151216 4014
rect 150912 4004 151228 4010
rect 150912 3998 151176 4004
rect 151176 3946 151228 3952
rect 153384 2848 153436 2854
rect 153384 2790 153436 2796
rect 149058 2479 149114 2488
rect 150808 2508 150860 2514
rect 150808 2450 150860 2456
rect 153396 2446 153424 2790
rect 156708 2689 156736 8366
rect 160112 8294 160140 8842
rect 167564 8634 167592 8842
rect 168760 8838 168788 8978
rect 171796 8974 171824 9522
rect 173084 8974 173112 10134
rect 175372 10124 175424 10130
rect 175372 10066 175424 10072
rect 171784 8968 171836 8974
rect 171784 8910 171836 8916
rect 173072 8968 173124 8974
rect 173072 8910 173124 8916
rect 171232 8900 171284 8906
rect 171232 8842 171284 8848
rect 175280 8900 175332 8906
rect 175280 8842 175332 8848
rect 168748 8832 168800 8838
rect 168748 8774 168800 8780
rect 167552 8628 167604 8634
rect 167552 8570 167604 8576
rect 160100 8288 160152 8294
rect 160100 8230 160152 8236
rect 158720 3596 158772 3602
rect 158720 3538 158772 3544
rect 158536 2848 158588 2854
rect 158536 2790 158588 2796
rect 156694 2680 156750 2689
rect 156694 2615 156750 2624
rect 153384 2440 153436 2446
rect 153384 2382 153436 2388
rect 151268 2304 151320 2310
rect 151268 2246 151320 2252
rect 152004 2304 152056 2310
rect 152004 2246 152056 2252
rect 148968 1896 149020 1902
rect 148968 1838 149020 1844
rect 148508 1624 148560 1630
rect 148508 1566 148560 1572
rect 148600 1624 148652 1630
rect 148600 1566 148652 1572
rect 148232 1556 148284 1562
rect 148232 1498 148284 1504
rect 150348 1556 150400 1562
rect 150348 1498 150400 1504
rect 147772 1488 147824 1494
rect 147772 1430 147824 1436
rect 147864 1488 147916 1494
rect 147864 1430 147916 1436
rect 146390 1391 146446 1400
rect 146668 1420 146720 1426
rect 146404 1154 146432 1391
rect 146668 1362 146720 1368
rect 147784 1290 147812 1430
rect 146484 1284 146536 1290
rect 146484 1226 146536 1232
rect 147772 1284 147824 1290
rect 147772 1226 147824 1232
rect 146392 1148 146444 1154
rect 146392 1090 146444 1096
rect 146496 950 146524 1226
rect 147876 1222 147904 1430
rect 147864 1216 147916 1222
rect 147864 1158 147916 1164
rect 148140 1216 148192 1222
rect 148140 1158 148192 1164
rect 148048 1148 148100 1154
rect 148048 1090 148100 1096
rect 148060 950 148088 1090
rect 146208 944 146260 950
rect 146208 886 146260 892
rect 146484 944 146536 950
rect 146484 886 146536 892
rect 148048 944 148100 950
rect 148048 886 148100 892
rect 146300 876 146352 882
rect 146300 818 146352 824
rect 128360 614 128412 620
rect 139320 610 139532 626
rect 145840 672 145892 678
rect 145840 614 145892 620
rect 139308 604 139532 610
rect 139360 598 139532 604
rect 139308 546 139360 552
rect 114560 264 114612 270
rect 114560 206 114612 212
rect 119436 264 119488 270
rect 119436 206 119488 212
rect 124496 264 124548 270
rect 124496 206 124548 212
rect 126428 264 126480 270
rect 126428 206 126480 212
rect 67568 8 67580 64
rect 67636 8 67660 64
rect 67716 8 67740 64
rect 67796 8 67820 64
rect 67876 8 67888 64
rect 67568 -4 67888 8
rect 75000 60 75052 66
rect 146312 48 146340 818
rect 148152 218 148180 1158
rect 150360 1154 150388 1498
rect 150530 1456 150586 1465
rect 150530 1391 150586 1400
rect 150348 1148 150400 1154
rect 150348 1090 150400 1096
rect 150440 1148 150492 1154
rect 150440 1090 150492 1096
rect 150452 950 150480 1090
rect 150544 950 150572 1391
rect 151280 1290 151308 2246
rect 152016 2038 152044 2246
rect 152004 2032 152056 2038
rect 152004 1974 152056 1980
rect 153396 1494 153424 2382
rect 158548 2378 158576 2790
rect 158536 2372 158588 2378
rect 158536 2314 158588 2320
rect 156420 2304 156472 2310
rect 156420 2246 156472 2252
rect 157156 2304 157208 2310
rect 157156 2246 157208 2252
rect 156432 1494 156460 2246
rect 157168 1970 157196 2246
rect 157156 1964 157208 1970
rect 157156 1906 157208 1912
rect 157248 1896 157300 1902
rect 157248 1838 157300 1844
rect 153384 1488 153436 1494
rect 153384 1430 153436 1436
rect 154580 1488 154632 1494
rect 156420 1488 156472 1494
rect 154580 1430 154632 1436
rect 154670 1456 154726 1465
rect 151268 1284 151320 1290
rect 151268 1226 151320 1232
rect 151360 1216 151412 1222
rect 151544 1216 151596 1222
rect 151412 1164 151544 1170
rect 151360 1158 151596 1164
rect 151372 1142 151584 1158
rect 152372 1148 152424 1154
rect 152372 1090 152424 1096
rect 150440 944 150492 950
rect 150440 886 150492 892
rect 150532 944 150584 950
rect 150532 886 150584 892
rect 152384 746 152412 1090
rect 154592 950 154620 1430
rect 156420 1430 156472 1436
rect 156970 1456 157026 1465
rect 154670 1391 154726 1400
rect 156970 1391 157026 1400
rect 157154 1456 157210 1465
rect 157154 1391 157210 1400
rect 154580 944 154632 950
rect 154580 886 154632 892
rect 154580 808 154632 814
rect 154684 796 154712 1391
rect 156984 1222 157012 1391
rect 157168 1290 157196 1391
rect 157260 1290 157288 1838
rect 158548 1766 158576 2314
rect 158536 1760 158588 1766
rect 158732 1737 158760 3538
rect 166908 2916 166960 2922
rect 166908 2858 166960 2864
rect 163688 2848 163740 2854
rect 163688 2790 163740 2796
rect 158902 2544 158958 2553
rect 158902 2479 158958 2488
rect 158916 2446 158944 2479
rect 158904 2440 158956 2446
rect 158904 2382 158956 2388
rect 161940 2440 161992 2446
rect 161940 2382 161992 2388
rect 161572 2304 161624 2310
rect 161572 2246 161624 2252
rect 158996 1896 159048 1902
rect 158996 1838 159048 1844
rect 158536 1702 158588 1708
rect 158718 1728 158774 1737
rect 158718 1663 158774 1672
rect 157432 1420 157484 1426
rect 157352 1380 157432 1408
rect 157156 1284 157208 1290
rect 157156 1226 157208 1232
rect 157248 1284 157300 1290
rect 157248 1226 157300 1232
rect 156880 1216 156932 1222
rect 156880 1158 156932 1164
rect 156972 1216 157024 1222
rect 156972 1158 157024 1164
rect 156788 1148 156840 1154
rect 156788 1090 156840 1096
rect 156696 1080 156748 1086
rect 156696 1022 156748 1028
rect 154632 768 154712 796
rect 154580 750 154632 756
rect 152372 740 152424 746
rect 152372 682 152424 688
rect 156708 354 156736 1022
rect 156800 490 156828 1090
rect 156892 796 156920 1158
rect 156984 1018 157196 1034
rect 157352 1018 157380 1380
rect 157432 1362 157484 1368
rect 158904 1148 158956 1154
rect 158904 1090 158956 1096
rect 157524 1080 157576 1086
rect 157524 1022 157576 1028
rect 156972 1012 157196 1018
rect 157024 1006 157196 1012
rect 156972 954 157024 960
rect 157168 864 157196 1006
rect 157340 1012 157392 1018
rect 157340 954 157392 960
rect 157432 1012 157484 1018
rect 157432 954 157484 960
rect 157444 864 157472 954
rect 157168 836 157472 864
rect 156892 768 157196 796
rect 157168 610 157196 768
rect 157156 604 157208 610
rect 157156 546 157208 552
rect 157248 536 157300 542
rect 156800 484 157248 490
rect 157536 490 157564 1022
rect 158916 542 158944 1090
rect 159008 610 159036 1838
rect 161204 1760 161256 1766
rect 161204 1702 161256 1708
rect 159088 876 159140 882
rect 159088 818 159140 824
rect 158996 604 159048 610
rect 158996 546 159048 552
rect 156800 478 157300 484
rect 156800 462 157288 478
rect 157352 462 157564 490
rect 158904 536 158956 542
rect 159100 490 159128 818
rect 161216 746 161244 1702
rect 161584 1562 161612 2246
rect 161952 1834 161980 2382
rect 163700 2378 163728 2790
rect 164146 2680 164202 2689
rect 164146 2615 164202 2624
rect 163688 2372 163740 2378
rect 163688 2314 163740 2320
rect 162308 2304 162360 2310
rect 162308 2246 162360 2252
rect 162320 1902 162348 2246
rect 162308 1896 162360 1902
rect 162308 1838 162360 1844
rect 163700 1834 163728 2314
rect 164160 2310 164188 2615
rect 164148 2304 164200 2310
rect 164148 2246 164200 2252
rect 161940 1828 161992 1834
rect 161940 1770 161992 1776
rect 163688 1828 163740 1834
rect 163688 1770 163740 1776
rect 163964 1828 164016 1834
rect 163964 1770 164016 1776
rect 163976 1698 164004 1770
rect 163964 1692 164016 1698
rect 163964 1634 164016 1640
rect 161572 1556 161624 1562
rect 161572 1498 161624 1504
rect 161756 1556 161808 1562
rect 161756 1498 161808 1504
rect 166816 1556 166868 1562
rect 166816 1498 166868 1504
rect 161768 814 161796 1498
rect 166828 1426 166856 1498
rect 166724 1420 166776 1426
rect 166724 1362 166776 1368
rect 166816 1420 166868 1426
rect 166816 1362 166868 1368
rect 166736 1306 166764 1362
rect 166736 1278 166856 1306
rect 166828 1154 166856 1278
rect 166724 1148 166776 1154
rect 166724 1090 166776 1096
rect 166816 1148 166868 1154
rect 166816 1090 166868 1096
rect 161756 808 161808 814
rect 161756 750 161808 756
rect 166736 746 166764 1090
rect 161204 740 161256 746
rect 161204 682 161256 688
rect 166724 740 166776 746
rect 166724 682 166776 688
rect 164056 672 164108 678
rect 164332 672 164384 678
rect 164108 632 164332 660
rect 164056 614 164108 620
rect 164332 614 164384 620
rect 166264 672 166316 678
rect 166632 672 166684 678
rect 166316 632 166632 660
rect 166264 614 166316 620
rect 166632 614 166684 620
rect 158904 478 158956 484
rect 159008 474 159128 490
rect 166264 536 166316 542
rect 166540 536 166592 542
rect 166316 496 166540 524
rect 166264 478 166316 484
rect 166540 478 166592 484
rect 158996 468 159128 474
rect 157352 354 157380 462
rect 159048 462 159128 468
rect 158996 410 159048 416
rect 166920 406 166948 2858
rect 168380 2848 168432 2854
rect 168380 2790 168432 2796
rect 168392 2378 168420 2790
rect 168380 2372 168432 2378
rect 168380 2314 168432 2320
rect 167460 2304 167512 2310
rect 167460 2246 167512 2252
rect 167472 1834 167500 2246
rect 167460 1828 167512 1834
rect 167460 1770 167512 1776
rect 168194 1728 168250 1737
rect 167196 1686 167500 1714
rect 167000 1420 167052 1426
rect 167052 1380 167132 1408
rect 167000 1362 167052 1368
rect 167104 1222 167132 1380
rect 167000 1216 167052 1222
rect 167000 1158 167052 1164
rect 167092 1216 167144 1222
rect 167092 1158 167144 1164
rect 167012 1034 167040 1158
rect 167196 1154 167224 1686
rect 167472 1562 167500 1686
rect 168104 1692 168156 1698
rect 168194 1663 168250 1672
rect 168288 1692 168340 1698
rect 168104 1634 168156 1640
rect 167460 1556 167512 1562
rect 167460 1498 167512 1504
rect 168116 1154 168144 1634
rect 167184 1148 167236 1154
rect 167184 1090 167236 1096
rect 168104 1148 168156 1154
rect 168104 1090 168156 1096
rect 167012 1018 167224 1034
rect 167012 1012 167236 1018
rect 167012 1006 167184 1012
rect 167184 954 167236 960
rect 168104 944 168156 950
rect 168104 886 168156 892
rect 168116 542 168144 886
rect 168208 814 168236 1663
rect 168288 1634 168340 1640
rect 168300 882 168328 1634
rect 168392 1465 168420 2314
rect 169300 2304 169352 2310
rect 169298 2272 169300 2281
rect 171140 2304 171192 2310
rect 169352 2272 169354 2281
rect 171140 2246 171192 2252
rect 169298 2207 169354 2216
rect 168656 1488 168708 1494
rect 168378 1456 168434 1465
rect 168378 1391 168434 1400
rect 168562 1456 168618 1465
rect 168656 1430 168708 1436
rect 168562 1391 168618 1400
rect 168288 876 168340 882
rect 168288 818 168340 824
rect 168196 808 168248 814
rect 168196 750 168248 756
rect 168288 740 168340 746
rect 168576 728 168604 1391
rect 168340 700 168604 728
rect 168288 682 168340 688
rect 168472 604 168524 610
rect 168668 592 168696 1430
rect 170864 1148 170916 1154
rect 170864 1090 170916 1096
rect 170956 1148 171008 1154
rect 170956 1090 171008 1096
rect 170876 678 170904 1090
rect 170968 950 170996 1090
rect 171152 1018 171180 2246
rect 171244 2145 171272 8842
rect 175292 8537 175320 8842
rect 175384 8634 175412 10066
rect 175476 8838 175504 11766
rect 194968 11756 195020 11762
rect 194968 11698 195020 11704
rect 184388 11620 184440 11626
rect 184388 11562 184440 11568
rect 184204 11212 184256 11218
rect 184204 11154 184256 11160
rect 176660 10260 176712 10266
rect 176660 10202 176712 10208
rect 176292 10124 176344 10130
rect 176292 10066 176344 10072
rect 176304 8974 176332 10066
rect 176292 8968 176344 8974
rect 176292 8910 176344 8916
rect 175464 8832 175516 8838
rect 175464 8774 175516 8780
rect 175372 8628 175424 8634
rect 175372 8570 175424 8576
rect 175278 8528 175334 8537
rect 175278 8463 175334 8472
rect 172518 8392 172574 8401
rect 172518 8327 172574 8336
rect 172532 2582 172560 8327
rect 176672 8265 176700 10202
rect 178040 9920 178092 9926
rect 178040 9862 178092 9868
rect 178052 9586 178080 9862
rect 178040 9580 178092 9586
rect 178040 9522 178092 9528
rect 176752 9036 176804 9042
rect 176752 8978 176804 8984
rect 176658 8256 176714 8265
rect 176658 8191 176714 8200
rect 173992 2848 174044 2854
rect 173992 2790 174044 2796
rect 172520 2576 172572 2582
rect 172520 2518 172572 2524
rect 172612 2576 172664 2582
rect 172612 2518 172664 2524
rect 172624 2394 172652 2518
rect 172532 2366 172652 2394
rect 174004 2378 174032 2790
rect 176764 2582 176792 8978
rect 179420 8900 179472 8906
rect 179420 8842 179472 8848
rect 179432 3602 179460 8842
rect 184216 8537 184244 11154
rect 184400 9586 184428 11562
rect 186688 11348 186740 11354
rect 186688 11290 186740 11296
rect 186240 10118 186544 10146
rect 186240 10062 186268 10118
rect 186228 10056 186280 10062
rect 186228 9998 186280 10004
rect 186320 10056 186372 10062
rect 186320 9998 186372 10004
rect 184388 9580 184440 9586
rect 184388 9522 184440 9528
rect 184202 8528 184258 8537
rect 184202 8463 184258 8472
rect 186332 8362 186360 9998
rect 186412 8900 186464 8906
rect 186412 8842 186464 8848
rect 186320 8356 186372 8362
rect 186320 8298 186372 8304
rect 182914 7304 182970 7313
rect 182914 7239 182970 7248
rect 179420 3596 179472 3602
rect 179420 3538 179472 3544
rect 180800 3596 180852 3602
rect 180800 3538 180852 3544
rect 178040 2848 178092 2854
rect 178040 2790 178092 2796
rect 179144 2848 179196 2854
rect 179144 2790 179196 2796
rect 176752 2576 176804 2582
rect 176752 2518 176804 2524
rect 177212 2576 177264 2582
rect 177212 2518 177264 2524
rect 177224 2446 177252 2518
rect 177212 2440 177264 2446
rect 177212 2382 177264 2388
rect 173992 2372 174044 2378
rect 171230 2136 171286 2145
rect 171230 2071 171286 2080
rect 172532 1766 172560 2366
rect 173992 2314 174044 2320
rect 175004 2372 175056 2378
rect 175004 2314 175056 2320
rect 172612 2304 172664 2310
rect 172612 2246 172664 2252
rect 172624 1766 172652 2246
rect 172520 1760 172572 1766
rect 172520 1702 172572 1708
rect 172612 1760 172664 1766
rect 172612 1702 172664 1708
rect 173070 1456 173126 1465
rect 173070 1391 173126 1400
rect 172244 1080 172296 1086
rect 172244 1022 172296 1028
rect 172336 1080 172388 1086
rect 172336 1022 172388 1028
rect 171140 1012 171192 1018
rect 171140 954 171192 960
rect 172256 950 172284 1022
rect 170956 944 171008 950
rect 170956 886 171008 892
rect 172244 944 172296 950
rect 172244 886 172296 892
rect 171048 808 171100 814
rect 170968 768 171048 796
rect 170864 672 170916 678
rect 170864 614 170916 620
rect 168524 564 168696 592
rect 168472 546 168524 552
rect 168104 536 168156 542
rect 168104 478 168156 484
rect 170404 536 170456 542
rect 170968 524 170996 768
rect 171048 750 171100 756
rect 172348 746 172376 1022
rect 172336 740 172388 746
rect 172336 682 172388 688
rect 172796 672 172848 678
rect 172796 614 172848 620
rect 170456 496 170996 524
rect 170404 478 170456 484
rect 172808 490 172836 614
rect 173084 610 173112 1391
rect 173256 1148 173308 1154
rect 173256 1090 173308 1096
rect 173348 1148 173400 1154
rect 173348 1090 173400 1096
rect 173164 740 173216 746
rect 173164 682 173216 688
rect 173072 604 173124 610
rect 173072 546 173124 552
rect 173176 490 173204 682
rect 172808 462 173204 490
rect 156708 326 157380 354
rect 166908 400 166960 406
rect 166908 342 166960 348
rect 147968 190 148180 218
rect 147968 66 147996 190
rect 173268 66 173296 1090
rect 173360 814 173388 1090
rect 173348 808 173400 814
rect 173348 750 173400 756
rect 174004 610 174032 2314
rect 174452 2304 174504 2310
rect 174452 2246 174504 2252
rect 174636 2304 174688 2310
rect 174636 2246 174688 2252
rect 174464 2145 174492 2246
rect 174450 2136 174506 2145
rect 174450 2071 174506 2080
rect 174648 1562 174676 2246
rect 174636 1556 174688 1562
rect 174636 1498 174688 1504
rect 174820 1556 174872 1562
rect 174820 1498 174872 1504
rect 173992 604 174044 610
rect 173992 546 174044 552
rect 174832 66 174860 1498
rect 175016 746 175044 2314
rect 178052 1737 178080 2790
rect 179156 2446 179184 2790
rect 180812 2582 180840 3538
rect 181076 3120 181128 3126
rect 181076 3062 181128 3068
rect 180800 2576 180852 2582
rect 180800 2518 180852 2524
rect 179144 2440 179196 2446
rect 179144 2382 179196 2388
rect 179604 2304 179656 2310
rect 179604 2246 179656 2252
rect 178038 1728 178094 1737
rect 178038 1663 178094 1672
rect 178682 1728 178738 1737
rect 178682 1663 178738 1672
rect 176752 1488 176804 1494
rect 176382 1456 176438 1465
rect 176752 1430 176804 1436
rect 176936 1488 176988 1494
rect 176936 1430 176988 1436
rect 176382 1391 176438 1400
rect 176396 1222 176424 1391
rect 176384 1216 176436 1222
rect 176568 1216 176620 1222
rect 176384 1158 176436 1164
rect 176488 1164 176568 1170
rect 176488 1158 176620 1164
rect 176488 1142 176608 1158
rect 176488 1086 176516 1142
rect 176764 1086 176792 1430
rect 176476 1080 176528 1086
rect 176476 1022 176528 1028
rect 176752 1080 176804 1086
rect 176752 1022 176804 1028
rect 176948 950 176976 1430
rect 177488 1012 177540 1018
rect 177488 954 177540 960
rect 176936 944 176988 950
rect 176936 886 176988 892
rect 177500 864 177528 954
rect 177948 944 178000 950
rect 177948 886 178000 892
rect 177672 876 177724 882
rect 177500 836 177672 864
rect 177672 818 177724 824
rect 177028 808 177080 814
rect 177960 762 177988 886
rect 178696 882 178724 1663
rect 179616 1562 179644 2246
rect 179512 1556 179564 1562
rect 179512 1498 179564 1504
rect 179604 1556 179656 1562
rect 179604 1498 179656 1504
rect 179524 1442 179552 1498
rect 181088 1494 181116 3062
rect 182928 2582 182956 7239
rect 184204 3052 184256 3058
rect 184204 2994 184256 3000
rect 183560 2848 183612 2854
rect 183560 2790 183612 2796
rect 182916 2576 182968 2582
rect 182916 2518 182968 2524
rect 182928 2446 182956 2518
rect 182916 2440 182968 2446
rect 182916 2382 182968 2388
rect 183572 2378 183600 2790
rect 183560 2372 183612 2378
rect 183560 2314 183612 2320
rect 182180 2304 182232 2310
rect 182180 2246 182232 2252
rect 183652 2304 183704 2310
rect 183652 2246 183704 2252
rect 182192 1494 182220 2246
rect 183664 1850 183692 2246
rect 183572 1822 183692 1850
rect 181076 1488 181128 1494
rect 179524 1414 179828 1442
rect 181076 1430 181128 1436
rect 181352 1488 181404 1494
rect 181352 1430 181404 1436
rect 182180 1488 182232 1494
rect 183572 1465 183600 1822
rect 183664 1550 184060 1578
rect 182180 1430 182232 1436
rect 183558 1456 183614 1465
rect 178684 876 178736 882
rect 178684 818 178736 824
rect 177080 756 177988 762
rect 177028 750 177988 756
rect 175004 740 175056 746
rect 177040 734 177988 750
rect 175004 682 175056 688
rect 179800 202 179828 1414
rect 181364 1086 181392 1430
rect 183664 1426 183692 1550
rect 183926 1456 183982 1465
rect 183558 1391 183614 1400
rect 183652 1420 183704 1426
rect 183926 1391 183982 1400
rect 183652 1362 183704 1368
rect 183812 1352 183864 1358
rect 183526 1300 183812 1306
rect 183526 1294 183864 1300
rect 183526 1290 183852 1294
rect 183514 1284 183852 1290
rect 183566 1278 183852 1284
rect 183514 1226 183566 1232
rect 181628 1216 181680 1222
rect 181548 1176 181628 1204
rect 181352 1080 181404 1086
rect 181352 1022 181404 1028
rect 181548 950 181576 1176
rect 181628 1158 181680 1164
rect 183652 1216 183704 1222
rect 183836 1216 183888 1222
rect 183704 1176 183836 1204
rect 183652 1158 183704 1164
rect 183836 1158 183888 1164
rect 183940 1154 183968 1391
rect 184032 1358 184060 1550
rect 184020 1352 184072 1358
rect 184020 1294 184072 1300
rect 183928 1148 183980 1154
rect 183928 1090 183980 1096
rect 184020 1148 184072 1154
rect 184020 1090 184072 1096
rect 183572 1040 183876 1068
rect 183572 1034 183600 1040
rect 183526 1018 183600 1034
rect 183514 1012 183600 1018
rect 183566 1006 183600 1012
rect 183848 1034 183876 1040
rect 184032 1034 184060 1090
rect 183848 1006 184060 1034
rect 184112 1080 184164 1086
rect 184112 1022 184164 1028
rect 183514 954 183566 960
rect 181536 944 181588 950
rect 181536 886 181588 892
rect 183652 944 183704 950
rect 183704 892 183784 898
rect 183652 886 183784 892
rect 183664 870 183784 886
rect 183756 864 183784 870
rect 183928 876 183980 882
rect 183756 836 183928 864
rect 183928 818 183980 824
rect 183514 808 183566 814
rect 183566 768 183784 796
rect 183514 750 183566 756
rect 183756 626 183784 768
rect 184124 626 184152 1022
rect 181260 604 181312 610
rect 181904 604 181956 610
rect 181312 564 181904 592
rect 181260 546 181312 552
rect 181904 546 181956 552
rect 183560 604 183612 610
rect 183756 598 184152 626
rect 183560 546 183612 552
rect 183572 354 183600 546
rect 184216 354 184244 2994
rect 184296 2440 184348 2446
rect 184296 2382 184348 2388
rect 183572 326 184244 354
rect 184308 218 184336 2382
rect 185492 2372 185544 2378
rect 185492 2314 185544 2320
rect 185504 1698 185532 2314
rect 185492 1692 185544 1698
rect 185492 1634 185544 1640
rect 185860 1692 185912 1698
rect 185860 1634 185912 1640
rect 185872 1154 185900 1634
rect 186134 1592 186190 1601
rect 186424 1578 186452 8842
rect 186516 8294 186544 10118
rect 186596 9716 186648 9722
rect 186596 9658 186648 9664
rect 186504 8288 186556 8294
rect 186504 8230 186556 8236
rect 186608 7750 186636 9658
rect 186596 7744 186648 7750
rect 186596 7686 186648 7692
rect 186700 7002 186728 11290
rect 187884 10260 187936 10266
rect 187884 10202 187936 10208
rect 187516 8968 187568 8974
rect 187700 8968 187752 8974
rect 187568 8916 187700 8922
rect 187516 8910 187752 8916
rect 187528 8894 187740 8910
rect 187792 8900 187844 8906
rect 187792 8842 187844 8848
rect 187516 8832 187568 8838
rect 187804 8786 187832 8842
rect 187568 8780 187832 8786
rect 187516 8774 187832 8780
rect 187528 8758 187832 8774
rect 187896 7410 187924 10202
rect 191472 9580 191524 9586
rect 191472 9522 191524 9528
rect 191484 9382 191512 9522
rect 194692 9512 194744 9518
rect 194692 9454 194744 9460
rect 191472 9376 191524 9382
rect 191472 9318 191524 9324
rect 191484 8430 191512 9318
rect 194704 9178 194732 9454
rect 194980 9178 195008 11698
rect 195060 11416 195112 11422
rect 195060 11358 195112 11364
rect 195072 9994 195100 11358
rect 195256 11218 195284 11766
rect 195612 11620 195664 11626
rect 195612 11562 195664 11568
rect 195520 11484 195572 11490
rect 195520 11426 195572 11432
rect 195244 11212 195296 11218
rect 195244 11154 195296 11160
rect 195336 11144 195388 11150
rect 195336 11086 195388 11092
rect 195244 11076 195296 11082
rect 195244 11018 195296 11024
rect 195152 10804 195204 10810
rect 195152 10746 195204 10752
rect 195164 9994 195192 10746
rect 195256 10674 195284 11018
rect 195348 10878 195376 11086
rect 195532 11014 195560 11426
rect 195624 11082 195652 11562
rect 195888 11484 195940 11490
rect 195888 11426 195940 11432
rect 195612 11076 195664 11082
rect 195612 11018 195664 11024
rect 195520 11008 195572 11014
rect 195520 10950 195572 10956
rect 195336 10872 195388 10878
rect 195336 10814 195388 10820
rect 195244 10668 195296 10674
rect 195244 10610 195296 10616
rect 195060 9988 195112 9994
rect 195060 9930 195112 9936
rect 195152 9988 195204 9994
rect 195152 9930 195204 9936
rect 195900 9586 195928 11426
rect 198836 11300 199156 11972
rect 199496 11960 199816 11972
rect 199496 11904 199508 11960
rect 199564 11904 199588 11960
rect 199644 11904 199668 11960
rect 199724 11904 199748 11960
rect 199804 11904 199816 11960
rect 199200 11892 199252 11898
rect 199200 11834 199252 11840
rect 199496 11880 199816 11904
rect 199936 11960 199988 11966
rect 199988 11908 200436 11914
rect 199936 11902 200436 11908
rect 199948 11898 200436 11902
rect 199948 11892 200448 11898
rect 199948 11886 200396 11892
rect 198836 11244 198848 11300
rect 198904 11244 198928 11300
rect 198984 11244 199008 11300
rect 199064 11244 199088 11300
rect 199144 11244 199156 11300
rect 198836 11220 199156 11244
rect 198464 11212 198516 11218
rect 198464 11154 198516 11160
rect 198836 11164 198848 11220
rect 198904 11164 198928 11220
rect 198984 11164 199008 11220
rect 199064 11164 199088 11220
rect 199144 11164 199156 11220
rect 198476 11098 198504 11154
rect 198836 11140 199156 11164
rect 198476 11070 198780 11098
rect 198556 11008 198608 11014
rect 198556 10950 198608 10956
rect 198464 10260 198516 10266
rect 198464 10202 198516 10208
rect 198370 10024 198426 10033
rect 198370 9959 198372 9968
rect 198424 9959 198426 9968
rect 198372 9930 198424 9936
rect 197818 9888 197874 9897
rect 197818 9823 197874 9832
rect 195888 9580 195940 9586
rect 195888 9522 195940 9528
rect 194692 9172 194744 9178
rect 194692 9114 194744 9120
rect 194968 9172 195020 9178
rect 194968 9114 195020 9120
rect 195612 8560 195664 8566
rect 195612 8502 195664 8508
rect 191472 8424 191524 8430
rect 191472 8366 191524 8372
rect 187884 7404 187936 7410
rect 187884 7346 187936 7352
rect 189172 7404 189224 7410
rect 189172 7346 189224 7352
rect 186688 6996 186740 7002
rect 186688 6938 186740 6944
rect 188068 3664 188120 3670
rect 188068 3606 188120 3612
rect 187332 2644 187384 2650
rect 187332 2586 187384 2592
rect 187424 2644 187476 2650
rect 187424 2586 187476 2592
rect 186780 2372 186832 2378
rect 186780 2314 186832 2320
rect 186872 2372 186924 2378
rect 186872 2314 186924 2320
rect 186190 1550 186452 1578
rect 186134 1527 186190 1536
rect 186688 1488 186740 1494
rect 186688 1430 186740 1436
rect 186148 1290 186452 1306
rect 186136 1284 186464 1290
rect 186188 1278 186412 1284
rect 186136 1226 186188 1232
rect 186412 1226 186464 1232
rect 186228 1216 186280 1222
rect 186228 1158 186280 1164
rect 185860 1148 185912 1154
rect 185860 1090 185912 1096
rect 185952 1080 186004 1086
rect 186240 1068 186268 1158
rect 186700 1086 186728 1430
rect 186792 1154 186820 2314
rect 186884 1766 186912 2314
rect 186872 1760 186924 1766
rect 187344 1737 187372 2586
rect 187436 2446 187464 2586
rect 188080 2446 188108 3606
rect 189184 3194 189212 7346
rect 194520 3862 194824 3890
rect 189172 3188 189224 3194
rect 189172 3130 189224 3136
rect 192852 3052 192904 3058
rect 192852 2994 192904 3000
rect 189080 2848 189132 2854
rect 189080 2790 189132 2796
rect 190460 2848 190512 2854
rect 190460 2790 190512 2796
rect 187424 2440 187476 2446
rect 187424 2382 187476 2388
rect 188068 2440 188120 2446
rect 188068 2382 188120 2388
rect 189092 2378 189120 2790
rect 189080 2372 189132 2378
rect 189080 2314 189132 2320
rect 188344 1760 188396 1766
rect 186872 1702 186924 1708
rect 187330 1728 187386 1737
rect 188344 1702 188396 1708
rect 187330 1663 187386 1672
rect 188356 1494 188384 1702
rect 189092 1601 189120 2314
rect 190472 1873 190500 2790
rect 191748 2440 191800 2446
rect 191748 2382 191800 2388
rect 191104 2100 191156 2106
rect 191104 2042 191156 2048
rect 191116 1873 191144 2042
rect 190458 1864 190514 1873
rect 190458 1799 190514 1808
rect 191102 1864 191158 1873
rect 191102 1799 191158 1808
rect 189078 1592 189134 1601
rect 189078 1527 189134 1536
rect 188344 1488 188396 1494
rect 188344 1430 188396 1436
rect 190184 1488 190236 1494
rect 191760 1465 191788 2382
rect 190184 1430 190236 1436
rect 191746 1456 191802 1465
rect 186780 1148 186832 1154
rect 186780 1090 186832 1096
rect 186004 1040 186268 1068
rect 186688 1080 186740 1086
rect 185952 1022 186004 1028
rect 186688 1022 186740 1028
rect 186872 1080 186924 1086
rect 186872 1022 186924 1028
rect 186884 950 186912 1022
rect 187884 1012 187936 1018
rect 187884 954 187936 960
rect 185676 944 185728 950
rect 185676 886 185728 892
rect 186872 944 186924 950
rect 186872 886 186924 892
rect 185688 814 185716 886
rect 185676 808 185728 814
rect 185676 750 185728 756
rect 187896 746 187924 954
rect 190196 814 190224 1430
rect 191746 1391 191802 1400
rect 190184 808 190236 814
rect 190184 750 190236 756
rect 187884 740 187936 746
rect 187884 682 187936 688
rect 192864 542 192892 2994
rect 194520 2650 194548 3862
rect 194796 3738 194824 3862
rect 194692 3732 194744 3738
rect 194692 3674 194744 3680
rect 194784 3732 194836 3738
rect 194784 3674 194836 3680
rect 194704 3194 194732 3674
rect 195152 3664 195204 3670
rect 195204 3612 195376 3618
rect 195152 3606 195376 3612
rect 195164 3602 195376 3606
rect 195164 3596 195388 3602
rect 195164 3590 195336 3596
rect 195336 3538 195388 3544
rect 194692 3188 194744 3194
rect 194692 3130 194744 3136
rect 195152 2916 195204 2922
rect 195152 2858 195204 2864
rect 193220 2644 193272 2650
rect 193220 2586 193272 2592
rect 194508 2644 194560 2650
rect 194508 2586 194560 2592
rect 193232 2446 193260 2586
rect 195164 2446 195192 2858
rect 193220 2440 193272 2446
rect 193220 2382 193272 2388
rect 195152 2440 195204 2446
rect 195152 2382 195204 2388
rect 195336 2372 195388 2378
rect 195336 2314 195388 2320
rect 195060 2304 195112 2310
rect 195060 2246 195112 2252
rect 195152 2304 195204 2310
rect 195152 2246 195204 2252
rect 195072 2106 195100 2246
rect 195060 2100 195112 2106
rect 195060 2042 195112 2048
rect 192944 1760 192996 1766
rect 192944 1702 192996 1708
rect 192852 536 192904 542
rect 192852 478 192904 484
rect 192220 338 192892 354
rect 192208 332 192892 338
rect 192260 326 192892 332
rect 192208 274 192260 280
rect 183664 202 184336 218
rect 179788 196 179840 202
rect 179788 138 179840 144
rect 181260 196 181312 202
rect 181904 196 181956 202
rect 181312 156 181904 184
rect 181260 138 181312 144
rect 181904 138 181956 144
rect 183652 196 184336 202
rect 183704 190 184336 196
rect 183652 138 183704 144
rect 192864 66 192892 326
rect 192956 134 192984 1702
rect 195164 1601 195192 2246
rect 195150 1592 195206 1601
rect 195150 1527 195206 1536
rect 195348 1494 195376 2314
rect 195624 2038 195652 8502
rect 196716 6928 196768 6934
rect 196716 6870 196768 6876
rect 196164 3664 196216 3670
rect 196164 3606 196216 3612
rect 196176 3505 196204 3606
rect 195978 3496 196034 3505
rect 195978 3431 196034 3440
rect 196162 3496 196218 3505
rect 196162 3431 196218 3440
rect 195992 3058 196020 3431
rect 195980 3052 196032 3058
rect 195980 2994 196032 3000
rect 195980 2304 196032 2310
rect 195980 2246 196032 2252
rect 195612 2032 195664 2038
rect 195612 1974 195664 1980
rect 195992 1766 196020 2246
rect 196072 1964 196124 1970
rect 196072 1906 196124 1912
rect 195980 1760 196032 1766
rect 195980 1702 196032 1708
rect 195244 1488 195296 1494
rect 195150 1456 195206 1465
rect 195244 1430 195296 1436
rect 195336 1488 195388 1494
rect 195336 1430 195388 1436
rect 195150 1391 195206 1400
rect 195060 1148 195112 1154
rect 195060 1090 195112 1096
rect 194968 808 195020 814
rect 194968 750 195020 756
rect 194600 672 194652 678
rect 194652 632 194916 660
rect 194600 614 194652 620
rect 194324 536 194376 542
rect 194324 478 194376 484
rect 194336 354 194364 478
rect 194888 474 194916 632
rect 194980 610 195008 750
rect 194968 604 195020 610
rect 194968 546 195020 552
rect 195072 542 195100 1090
rect 195164 678 195192 1391
rect 195256 1086 195284 1430
rect 195244 1080 195296 1086
rect 195244 1022 195296 1028
rect 195244 876 195296 882
rect 195244 818 195296 824
rect 195152 672 195204 678
rect 195152 614 195204 620
rect 195060 536 195112 542
rect 195060 478 195112 484
rect 194876 468 194928 474
rect 194876 410 194928 416
rect 194336 326 195008 354
rect 195256 338 195284 818
rect 196084 610 196112 1906
rect 196728 1902 196756 6870
rect 197832 2446 197860 9823
rect 198476 9722 198504 10202
rect 198568 9994 198596 10950
rect 198648 10940 198700 10946
rect 198648 10882 198700 10888
rect 198660 10849 198688 10882
rect 198646 10840 198702 10849
rect 198646 10775 198702 10784
rect 198752 10674 198780 11070
rect 198836 11084 198848 11140
rect 198904 11084 198928 11140
rect 198984 11084 199008 11140
rect 199064 11084 199088 11140
rect 199144 11084 199156 11140
rect 198836 11060 199156 11084
rect 199212 11082 199240 11834
rect 199496 11824 199508 11880
rect 199564 11824 199588 11880
rect 199644 11824 199668 11880
rect 199724 11824 199748 11880
rect 199804 11824 199816 11880
rect 200396 11834 200448 11840
rect 199496 11800 199816 11824
rect 199496 11744 199508 11800
rect 199564 11744 199588 11800
rect 199644 11744 199668 11800
rect 199724 11744 199748 11800
rect 199804 11744 199816 11800
rect 199496 11720 199816 11744
rect 199384 11688 199436 11694
rect 199384 11630 199436 11636
rect 199496 11664 199508 11720
rect 199564 11664 199588 11720
rect 199644 11664 199668 11720
rect 199724 11664 199748 11720
rect 199804 11664 199816 11720
rect 199396 11529 199424 11630
rect 199382 11520 199438 11529
rect 199292 11484 199344 11490
rect 199382 11455 199438 11464
rect 199292 11426 199344 11432
rect 198836 11004 198848 11060
rect 198904 11004 198928 11060
rect 198984 11004 199008 11060
rect 199064 11004 199088 11060
rect 199144 11004 199156 11060
rect 199200 11076 199252 11082
rect 199200 11018 199252 11024
rect 198648 10668 198700 10674
rect 198648 10610 198700 10616
rect 198740 10668 198792 10674
rect 198740 10610 198792 10616
rect 198660 10266 198688 10610
rect 198648 10260 198700 10266
rect 198648 10202 198700 10208
rect 198646 10160 198702 10169
rect 198646 10095 198702 10104
rect 198556 9988 198608 9994
rect 198556 9930 198608 9936
rect 198464 9716 198516 9722
rect 198464 9658 198516 9664
rect 198660 8566 198688 10095
rect 198836 9274 199156 11004
rect 199304 10713 199332 11426
rect 199384 11348 199436 11354
rect 199384 11290 199436 11296
rect 199290 10704 199346 10713
rect 199290 10639 199346 10648
rect 199290 10568 199346 10577
rect 199290 10503 199346 10512
rect 199304 10470 199332 10503
rect 199396 10470 199424 11290
rect 199292 10464 199344 10470
rect 199292 10406 199344 10412
rect 199384 10464 199436 10470
rect 199384 10406 199436 10412
rect 199496 9818 199816 11664
rect 277124 11688 277176 11694
rect 205284 11626 205680 11642
rect 277124 11630 277176 11636
rect 205284 11620 205692 11626
rect 205284 11614 205640 11620
rect 199844 11552 199896 11558
rect 199844 11494 199896 11500
rect 202050 11520 202106 11529
rect 199856 11150 199884 11494
rect 202050 11455 202106 11464
rect 200856 11280 200908 11286
rect 200856 11222 200908 11228
rect 201316 11280 201368 11286
rect 201316 11222 201368 11228
rect 201960 11280 202012 11286
rect 201960 11222 202012 11228
rect 199936 11212 199988 11218
rect 199936 11154 199988 11160
rect 199844 11144 199896 11150
rect 199844 11086 199896 11092
rect 199948 11014 199976 11154
rect 199936 11008 199988 11014
rect 199936 10950 199988 10956
rect 199496 9766 199502 9818
rect 199554 9766 199566 9818
rect 199618 9766 199630 9818
rect 199682 9766 199694 9818
rect 199746 9766 199758 9818
rect 199810 9766 199816 9818
rect 199496 9648 199816 9766
rect 200868 9722 200896 11222
rect 201328 11014 201356 11222
rect 201316 11008 201368 11014
rect 201316 10950 201368 10956
rect 201408 11008 201460 11014
rect 201408 10950 201460 10956
rect 201224 10872 201276 10878
rect 200946 10840 201002 10849
rect 201420 10826 201448 10950
rect 201500 10940 201552 10946
rect 201500 10882 201552 10888
rect 201276 10820 201448 10826
rect 201224 10814 201448 10820
rect 201236 10798 201448 10814
rect 200946 10775 201002 10784
rect 200960 9722 200988 10775
rect 201512 10674 201540 10882
rect 201500 10668 201552 10674
rect 201500 10610 201552 10616
rect 201498 10432 201554 10441
rect 201498 10367 201554 10376
rect 200856 9716 200908 9722
rect 200856 9658 200908 9664
rect 200948 9716 201000 9722
rect 200948 9658 201000 9664
rect 199496 9592 199508 9648
rect 199564 9592 199588 9648
rect 199644 9592 199668 9648
rect 199724 9592 199748 9648
rect 199804 9592 199816 9648
rect 199496 9568 199816 9592
rect 199496 9512 199508 9568
rect 199564 9512 199588 9568
rect 199644 9512 199668 9568
rect 199724 9512 199748 9568
rect 199804 9512 199816 9568
rect 199496 9488 199816 9512
rect 199496 9432 199508 9488
rect 199564 9432 199588 9488
rect 199644 9432 199668 9488
rect 199724 9432 199748 9488
rect 199804 9432 199816 9488
rect 199496 9408 199816 9432
rect 199200 9376 199252 9382
rect 199200 9318 199252 9324
rect 199496 9352 199508 9408
rect 199564 9352 199588 9408
rect 199644 9352 199668 9408
rect 199724 9352 199748 9408
rect 199804 9352 199816 9408
rect 200764 9444 200816 9450
rect 200764 9386 200816 9392
rect 198836 9222 198842 9274
rect 198894 9222 198906 9274
rect 198958 9222 198970 9274
rect 199022 9222 199034 9274
rect 199086 9222 199098 9274
rect 199150 9222 199156 9274
rect 198836 8988 199156 9222
rect 198836 8932 198848 8988
rect 198904 8932 198928 8988
rect 198984 8932 199008 8988
rect 199064 8932 199088 8988
rect 199144 8932 199156 8988
rect 198836 8908 199156 8932
rect 198836 8852 198848 8908
rect 198904 8852 198928 8908
rect 198984 8852 199008 8908
rect 199064 8852 199088 8908
rect 199144 8852 199156 8908
rect 198836 8828 199156 8852
rect 198836 8772 198848 8828
rect 198904 8772 198928 8828
rect 198984 8772 199008 8828
rect 199064 8772 199088 8828
rect 199144 8772 199156 8828
rect 198836 8748 199156 8772
rect 198836 8692 198848 8748
rect 198904 8692 198928 8748
rect 198984 8692 199008 8748
rect 199064 8692 199088 8748
rect 199144 8692 199156 8748
rect 198648 8560 198700 8566
rect 198648 8502 198700 8508
rect 198740 8356 198792 8362
rect 198740 8298 198792 8304
rect 197820 2440 197872 2446
rect 197820 2382 197872 2388
rect 196716 1896 196768 1902
rect 196716 1838 196768 1844
rect 198752 1834 198780 8298
rect 198836 8186 199156 8692
rect 199212 8566 199240 9318
rect 199496 8730 199816 9352
rect 200776 8838 200804 9386
rect 200764 8832 200816 8838
rect 200764 8774 200816 8780
rect 199496 8678 199502 8730
rect 199554 8678 199566 8730
rect 199618 8678 199630 8730
rect 199682 8678 199694 8730
rect 199746 8678 199758 8730
rect 199810 8678 199816 8730
rect 199200 8560 199252 8566
rect 199200 8502 199252 8508
rect 198836 8134 198842 8186
rect 198894 8134 198906 8186
rect 198958 8134 198970 8186
rect 199022 8134 199034 8186
rect 199086 8134 199098 8186
rect 199150 8134 199156 8186
rect 198836 7098 199156 8134
rect 198836 7046 198842 7098
rect 198894 7084 198906 7098
rect 198958 7084 198970 7098
rect 199022 7084 199034 7098
rect 199086 7084 199098 7098
rect 198904 7046 198906 7084
rect 199086 7046 199088 7084
rect 199150 7046 199156 7098
rect 198836 7028 198848 7046
rect 198904 7028 198928 7046
rect 198984 7028 199008 7046
rect 199064 7028 199088 7046
rect 199144 7028 199156 7046
rect 198836 7004 199156 7028
rect 198836 6948 198848 7004
rect 198904 6948 198928 7004
rect 198984 6948 199008 7004
rect 199064 6948 199088 7004
rect 199144 6948 199156 7004
rect 198836 6924 199156 6948
rect 198836 6868 198848 6924
rect 198904 6868 198928 6924
rect 198984 6868 199008 6924
rect 199064 6868 199088 6924
rect 199144 6868 199156 6924
rect 198836 6844 199156 6868
rect 198836 6788 198848 6844
rect 198904 6788 198928 6844
rect 198984 6788 199008 6844
rect 199064 6788 199088 6844
rect 199144 6788 199156 6844
rect 198836 6010 199156 6788
rect 198836 5958 198842 6010
rect 198894 5958 198906 6010
rect 198958 5958 198970 6010
rect 199022 5958 199034 6010
rect 199086 5958 199098 6010
rect 199150 5958 199156 6010
rect 198836 5180 199156 5958
rect 198836 5124 198848 5180
rect 198904 5124 198928 5180
rect 198984 5124 199008 5180
rect 199064 5124 199088 5180
rect 199144 5124 199156 5180
rect 198836 5100 199156 5124
rect 198836 5044 198848 5100
rect 198904 5044 198928 5100
rect 198984 5044 199008 5100
rect 199064 5044 199088 5100
rect 199144 5044 199156 5100
rect 198836 5020 199156 5044
rect 198836 4964 198848 5020
rect 198904 4964 198928 5020
rect 198984 4964 199008 5020
rect 199064 4964 199088 5020
rect 199144 4964 199156 5020
rect 198836 4940 199156 4964
rect 198836 4922 198848 4940
rect 198904 4922 198928 4940
rect 198984 4922 199008 4940
rect 199064 4922 199088 4940
rect 199144 4922 199156 4940
rect 198836 4870 198842 4922
rect 198904 4884 198906 4922
rect 199086 4884 199088 4922
rect 198894 4870 198906 4884
rect 198958 4870 198970 4884
rect 199022 4870 199034 4884
rect 199086 4870 199098 4884
rect 199150 4870 199156 4922
rect 198836 3834 199156 4870
rect 198836 3782 198842 3834
rect 198894 3782 198906 3834
rect 198958 3782 198970 3834
rect 199022 3782 199034 3834
rect 199086 3782 199098 3834
rect 199150 3782 199156 3834
rect 198836 3276 199156 3782
rect 198836 3220 198848 3276
rect 198904 3220 198928 3276
rect 198984 3220 199008 3276
rect 199064 3220 199088 3276
rect 199144 3220 199156 3276
rect 198836 3196 199156 3220
rect 198836 3140 198848 3196
rect 198904 3140 198928 3196
rect 198984 3140 199008 3196
rect 199064 3140 199088 3196
rect 199144 3140 199156 3196
rect 198836 3116 199156 3140
rect 198836 3060 198848 3116
rect 198904 3060 198928 3116
rect 198984 3060 199008 3116
rect 199064 3060 199088 3116
rect 199144 3060 199156 3116
rect 198836 3036 199156 3060
rect 198836 2980 198848 3036
rect 198904 2980 198928 3036
rect 198984 2980 199008 3036
rect 199064 2980 199088 3036
rect 199144 2980 199156 3036
rect 198836 2746 199156 2980
rect 198836 2694 198842 2746
rect 198894 2694 198906 2746
rect 198958 2694 198970 2746
rect 199022 2694 199034 2746
rect 199086 2694 199098 2746
rect 199150 2694 199156 2746
rect 198740 1828 198792 1834
rect 198740 1770 198792 1776
rect 198836 964 199156 2694
rect 198740 944 198792 950
rect 198740 886 198792 892
rect 198836 908 198848 964
rect 198904 908 198928 964
rect 198984 908 199008 964
rect 199064 908 199088 964
rect 199144 908 199156 964
rect 198004 876 198056 882
rect 198004 818 198056 824
rect 196348 808 196400 814
rect 196348 750 196400 756
rect 195980 604 196032 610
rect 195980 546 196032 552
rect 196072 604 196124 610
rect 196072 546 196124 552
rect 194980 270 195008 326
rect 195244 332 195296 338
rect 195244 274 195296 280
rect 194968 264 195020 270
rect 194520 190 194916 218
rect 194968 206 195020 212
rect 195992 202 196020 546
rect 196360 542 196388 750
rect 196348 536 196400 542
rect 196348 478 196400 484
rect 198016 474 198044 818
rect 198004 468 198056 474
rect 198004 410 198056 416
rect 198752 406 198780 886
rect 198836 884 199156 908
rect 198836 828 198848 884
rect 198904 828 198928 884
rect 198984 828 199008 884
rect 199064 828 199088 884
rect 199144 828 199156 884
rect 198836 804 199156 828
rect 198836 748 198848 804
rect 198904 748 198928 804
rect 198984 748 199008 804
rect 199064 748 199088 804
rect 199144 748 199156 804
rect 198836 724 199156 748
rect 198836 668 198848 724
rect 198904 668 198928 724
rect 198984 668 199008 724
rect 199064 668 199088 724
rect 199144 668 199156 724
rect 198740 400 198792 406
rect 198740 342 198792 348
rect 192944 128 192996 134
rect 192944 70 192996 76
rect 194520 66 194548 190
rect 194600 128 194652 134
rect 194784 128 194836 134
rect 194652 76 194784 82
rect 194600 70 194836 76
rect 146392 60 146444 66
rect 146312 20 146392 48
rect 75000 2 75052 8
rect 146392 2 146444 8
rect 147956 60 148008 66
rect 147956 2 148008 8
rect 173256 60 173308 66
rect 173256 2 173308 8
rect 174820 60 174872 66
rect 174820 2 174872 8
rect 192852 60 192904 66
rect 192852 2 192904 8
rect 194508 60 194560 66
rect 194612 54 194824 70
rect 194888 66 194916 190
rect 195980 196 196032 202
rect 195980 138 196032 144
rect 194876 60 194928 66
rect 194508 2 194560 8
rect 194876 2 194928 8
rect 198836 -4 199156 668
rect 199496 7744 199816 8678
rect 199496 7688 199508 7744
rect 199564 7688 199588 7744
rect 199644 7688 199668 7744
rect 199724 7688 199748 7744
rect 199804 7688 199816 7744
rect 199496 7664 199816 7688
rect 199496 7642 199508 7664
rect 199564 7642 199588 7664
rect 199644 7642 199668 7664
rect 199724 7642 199748 7664
rect 199804 7642 199816 7664
rect 199496 7590 199502 7642
rect 199564 7608 199566 7642
rect 199746 7608 199748 7642
rect 199554 7590 199566 7608
rect 199618 7590 199630 7608
rect 199682 7590 199694 7608
rect 199746 7590 199758 7608
rect 199810 7590 199816 7642
rect 199496 7584 199816 7590
rect 199496 7528 199508 7584
rect 199564 7528 199588 7584
rect 199644 7528 199668 7584
rect 199724 7528 199748 7584
rect 199804 7528 199816 7584
rect 201512 7546 201540 10367
rect 201972 8294 202000 11222
rect 202064 8294 202092 11455
rect 202512 11280 202564 11286
rect 202512 11222 202564 11228
rect 202972 11280 203024 11286
rect 202972 11222 203024 11228
rect 203432 11280 203484 11286
rect 203432 11222 203484 11228
rect 205088 11280 205140 11286
rect 205088 11222 205140 11228
rect 202420 9512 202472 9518
rect 202420 9454 202472 9460
rect 201960 8288 202012 8294
rect 201960 8230 202012 8236
rect 202052 8288 202104 8294
rect 202052 8230 202104 8236
rect 199496 7504 199816 7528
rect 199496 7448 199508 7504
rect 199564 7448 199588 7504
rect 199644 7448 199668 7504
rect 199724 7448 199748 7504
rect 199804 7448 199816 7504
rect 201500 7540 201552 7546
rect 201500 7482 201552 7488
rect 199496 6554 199816 7448
rect 199496 6502 199502 6554
rect 199554 6502 199566 6554
rect 199618 6502 199630 6554
rect 199682 6502 199694 6554
rect 199746 6502 199758 6554
rect 199810 6502 199816 6554
rect 199496 5840 199816 6502
rect 199496 5784 199508 5840
rect 199564 5784 199588 5840
rect 199644 5784 199668 5840
rect 199724 5784 199748 5840
rect 199804 5784 199816 5840
rect 199496 5760 199816 5784
rect 199496 5704 199508 5760
rect 199564 5704 199588 5760
rect 199644 5704 199668 5760
rect 199724 5704 199748 5760
rect 199804 5704 199816 5760
rect 199496 5680 199816 5704
rect 199496 5624 199508 5680
rect 199564 5624 199588 5680
rect 199644 5624 199668 5680
rect 199724 5624 199748 5680
rect 199804 5624 199816 5680
rect 199496 5600 199816 5624
rect 199496 5544 199508 5600
rect 199564 5544 199588 5600
rect 199644 5544 199668 5600
rect 199724 5544 199748 5600
rect 199804 5544 199816 5600
rect 199496 5466 199816 5544
rect 199496 5414 199502 5466
rect 199554 5414 199566 5466
rect 199618 5414 199630 5466
rect 199682 5414 199694 5466
rect 199746 5414 199758 5466
rect 199810 5414 199816 5466
rect 199496 4378 199816 5414
rect 199496 4326 199502 4378
rect 199554 4326 199566 4378
rect 199618 4326 199630 4378
rect 199682 4326 199694 4378
rect 199746 4326 199758 4378
rect 199810 4326 199816 4378
rect 199496 3936 199816 4326
rect 199496 3880 199508 3936
rect 199564 3880 199588 3936
rect 199644 3880 199668 3936
rect 199724 3880 199748 3936
rect 199804 3880 199816 3936
rect 199496 3856 199816 3880
rect 199496 3800 199508 3856
rect 199564 3800 199588 3856
rect 199644 3800 199668 3856
rect 199724 3800 199748 3856
rect 199804 3800 199816 3856
rect 199496 3776 199816 3800
rect 199496 3720 199508 3776
rect 199564 3720 199588 3776
rect 199644 3720 199668 3776
rect 199724 3720 199748 3776
rect 199804 3720 199816 3776
rect 199496 3696 199816 3720
rect 199496 3640 199508 3696
rect 199564 3640 199588 3696
rect 199644 3640 199668 3696
rect 199724 3640 199748 3696
rect 199804 3640 199816 3696
rect 199496 3290 199816 3640
rect 199496 3238 199502 3290
rect 199554 3238 199566 3290
rect 199618 3238 199630 3290
rect 199682 3238 199694 3290
rect 199746 3238 199758 3290
rect 199810 3238 199816 3290
rect 199496 2202 199816 3238
rect 202432 2922 202460 9454
rect 202524 7993 202552 11222
rect 202880 10668 202932 10674
rect 202880 10610 202932 10616
rect 202892 9994 202920 10610
rect 202880 9988 202932 9994
rect 202880 9930 202932 9936
rect 202984 8265 203012 11222
rect 203444 10470 203472 11222
rect 203984 11212 204036 11218
rect 203984 11154 204036 11160
rect 204536 11212 204588 11218
rect 204536 11154 204588 11160
rect 203996 10577 204024 11154
rect 203982 10568 204038 10577
rect 203982 10503 204038 10512
rect 203432 10464 203484 10470
rect 203432 10406 203484 10412
rect 203524 10464 203576 10470
rect 203524 10406 203576 10412
rect 203536 10169 203564 10406
rect 203706 10296 203762 10305
rect 203706 10231 203762 10240
rect 203522 10160 203578 10169
rect 203522 10095 203578 10104
rect 203616 9988 203668 9994
rect 203616 9930 203668 9936
rect 203628 9586 203656 9930
rect 203616 9580 203668 9586
rect 203616 9522 203668 9528
rect 202970 8256 203026 8265
rect 202970 8191 203026 8200
rect 202510 7984 202566 7993
rect 202510 7919 202566 7928
rect 202694 7984 202750 7993
rect 202694 7919 202750 7928
rect 202708 6934 202736 7919
rect 202696 6928 202748 6934
rect 202696 6870 202748 6876
rect 202420 2916 202472 2922
rect 202420 2858 202472 2864
rect 200028 2848 200080 2854
rect 200028 2790 200080 2796
rect 200040 2446 200068 2790
rect 203720 2774 203748 10231
rect 204548 10033 204576 11154
rect 205100 10674 205128 11222
rect 205088 10668 205140 10674
rect 205088 10610 205140 10616
rect 205180 10668 205232 10674
rect 205180 10610 205232 10616
rect 205192 10470 205220 10610
rect 205180 10464 205232 10470
rect 205180 10406 205232 10412
rect 204534 10024 204590 10033
rect 204534 9959 204590 9968
rect 205284 9722 205312 11614
rect 205640 11562 205692 11568
rect 258724 11552 258776 11558
rect 205454 11520 205510 11529
rect 205454 11455 205510 11464
rect 207294 11520 207350 11529
rect 207294 11455 207350 11464
rect 213642 11520 213698 11529
rect 213642 11455 213698 11464
rect 214378 11520 214434 11529
rect 258724 11494 258776 11500
rect 214378 11455 214380 11464
rect 205468 11082 205496 11455
rect 206192 11280 206244 11286
rect 205652 11206 206140 11234
rect 206192 11222 206244 11228
rect 205652 11082 205680 11206
rect 205456 11076 205508 11082
rect 205456 11018 205508 11024
rect 205548 11076 205600 11082
rect 205548 11018 205600 11024
rect 205640 11076 205692 11082
rect 205640 11018 205692 11024
rect 205560 10384 205588 11018
rect 205640 10736 205692 10742
rect 205732 10736 205784 10742
rect 205640 10678 205692 10684
rect 205730 10704 205732 10713
rect 205784 10704 205786 10713
rect 205652 10470 205680 10678
rect 205730 10639 205786 10648
rect 206112 10606 206140 11206
rect 206008 10600 206060 10606
rect 205822 10568 205878 10577
rect 206008 10542 206060 10548
rect 206100 10600 206152 10606
rect 206100 10542 206152 10548
rect 205822 10503 205878 10512
rect 205640 10464 205692 10470
rect 205640 10406 205692 10412
rect 205836 10402 205864 10503
rect 205376 10356 205588 10384
rect 205824 10396 205876 10402
rect 205376 10266 205404 10356
rect 205824 10338 205876 10344
rect 205640 10328 205692 10334
rect 205640 10270 205692 10276
rect 205364 10260 205416 10266
rect 205364 10202 205416 10208
rect 205652 10146 205680 10270
rect 206020 10266 206048 10542
rect 206204 10441 206232 11222
rect 207308 11150 207336 11455
rect 212908 11416 212960 11422
rect 212092 11364 212908 11370
rect 212092 11358 212960 11364
rect 212092 11342 212948 11358
rect 207480 11280 207532 11286
rect 207480 11222 207532 11228
rect 208124 11280 208176 11286
rect 208124 11222 208176 11228
rect 208584 11280 208636 11286
rect 208584 11222 208636 11228
rect 209964 11280 210016 11286
rect 209964 11222 210016 11228
rect 210700 11280 210752 11286
rect 210700 11222 210752 11228
rect 211160 11280 211212 11286
rect 211160 11222 211212 11228
rect 211804 11280 211856 11286
rect 211804 11222 211856 11228
rect 207296 11144 207348 11150
rect 207296 11086 207348 11092
rect 207020 11076 207072 11082
rect 207020 11018 207072 11024
rect 207388 11076 207440 11082
rect 207388 11018 207440 11024
rect 207032 10810 207060 11018
rect 207296 11008 207348 11014
rect 207296 10950 207348 10956
rect 206928 10804 206980 10810
rect 206928 10746 206980 10752
rect 207020 10804 207072 10810
rect 207020 10746 207072 10752
rect 206940 10538 206968 10746
rect 206836 10532 206888 10538
rect 206836 10474 206888 10480
rect 206928 10532 206980 10538
rect 206928 10474 206980 10480
rect 206190 10432 206246 10441
rect 206190 10367 206246 10376
rect 206742 10296 206798 10305
rect 206008 10260 206060 10266
rect 206742 10231 206798 10240
rect 206008 10202 206060 10208
rect 205652 10118 205864 10146
rect 205640 10056 205692 10062
rect 205638 10024 205640 10033
rect 205692 10024 205694 10033
rect 205836 9994 205864 10118
rect 206756 10062 206784 10231
rect 206848 10062 206876 10474
rect 206744 10056 206796 10062
rect 206744 9998 206796 10004
rect 206836 10056 206888 10062
rect 207308 10033 207336 10950
rect 207400 10577 207428 11018
rect 207386 10568 207442 10577
rect 207386 10503 207442 10512
rect 206836 9998 206888 10004
rect 207294 10024 207350 10033
rect 205638 9959 205694 9968
rect 205824 9988 205876 9994
rect 207294 9959 207350 9968
rect 205824 9930 205876 9936
rect 205546 9888 205602 9897
rect 205546 9823 205602 9832
rect 206282 9888 206338 9897
rect 206282 9823 206338 9832
rect 205560 9722 205588 9823
rect 205272 9716 205324 9722
rect 205272 9658 205324 9664
rect 205548 9716 205600 9722
rect 205548 9658 205600 9664
rect 206296 9586 206324 9823
rect 206284 9580 206336 9586
rect 206284 9522 206336 9528
rect 205456 9512 205508 9518
rect 205456 9454 205508 9460
rect 205364 4140 205416 4146
rect 205364 4082 205416 4088
rect 205088 2848 205140 2854
rect 205088 2790 205140 2796
rect 203076 2746 203748 2774
rect 203076 2446 203104 2746
rect 205100 2446 205128 2790
rect 205376 2650 205404 4082
rect 205468 3126 205496 9454
rect 207492 8294 207520 11222
rect 207480 8288 207532 8294
rect 207480 8230 207532 8236
rect 205456 3120 205508 3126
rect 205456 3062 205508 3068
rect 208136 2774 208164 11222
rect 208596 7410 208624 11222
rect 209976 10470 210004 11222
rect 210056 11212 210108 11218
rect 210056 11154 210108 11160
rect 209964 10464 210016 10470
rect 209964 10406 210016 10412
rect 208674 10160 208730 10169
rect 208674 10095 208730 10104
rect 208584 7404 208636 7410
rect 208584 7346 208636 7352
rect 208688 2774 208716 10095
rect 210068 8129 210096 11154
rect 210240 10464 210292 10470
rect 210240 10406 210292 10412
rect 210330 10432 210386 10441
rect 210148 10328 210200 10334
rect 210146 10296 210148 10305
rect 210200 10296 210202 10305
rect 210146 10231 210202 10240
rect 210252 9897 210280 10406
rect 210330 10367 210332 10376
rect 210384 10367 210386 10376
rect 210332 10338 210384 10344
rect 210238 9888 210294 9897
rect 210238 9823 210294 9832
rect 210240 9512 210292 9518
rect 210240 9454 210292 9460
rect 210252 9217 210280 9454
rect 210238 9208 210294 9217
rect 210238 9143 210294 9152
rect 210054 8120 210110 8129
rect 210054 8055 210110 8064
rect 210712 7478 210740 11222
rect 211068 11076 211120 11082
rect 211068 11018 211120 11024
rect 211080 9586 211108 11018
rect 211172 10538 211200 11222
rect 211160 10532 211212 10538
rect 211160 10474 211212 10480
rect 211252 10532 211304 10538
rect 211252 10474 211304 10480
rect 211264 9926 211292 10474
rect 211252 9920 211304 9926
rect 211252 9862 211304 9868
rect 211068 9580 211120 9586
rect 211068 9522 211120 9528
rect 210700 7472 210752 7478
rect 210700 7414 210752 7420
rect 210424 4140 210476 4146
rect 210424 4082 210476 4088
rect 210436 3738 210464 4082
rect 210424 3732 210476 3738
rect 210424 3674 210476 3680
rect 210516 3120 210568 3126
rect 210516 3062 210568 3068
rect 210240 2848 210292 2854
rect 210240 2790 210292 2796
rect 208136 2746 208256 2774
rect 205364 2644 205416 2650
rect 205364 2586 205416 2592
rect 200028 2440 200080 2446
rect 200028 2382 200080 2388
rect 203064 2440 203116 2446
rect 203064 2382 203116 2388
rect 205088 2440 205140 2446
rect 205088 2382 205140 2388
rect 200212 2304 200264 2310
rect 200212 2246 200264 2252
rect 202788 2304 202840 2310
rect 202788 2246 202840 2252
rect 199496 2150 199502 2202
rect 199554 2150 199566 2202
rect 199618 2150 199630 2202
rect 199682 2150 199694 2202
rect 199746 2150 199758 2202
rect 199810 2150 199816 2202
rect 199496 304 199816 2150
rect 200224 2038 200252 2246
rect 200212 2032 200264 2038
rect 200212 1974 200264 1980
rect 202800 338 202828 2246
rect 199496 248 199508 304
rect 199564 248 199588 304
rect 199644 248 199668 304
rect 199724 248 199748 304
rect 199804 248 199816 304
rect 202788 332 202840 338
rect 202788 274 202840 280
rect 199496 224 199816 248
rect 199496 168 199508 224
rect 199564 168 199588 224
rect 199644 168 199668 224
rect 199724 168 199748 224
rect 199804 168 199816 224
rect 199496 144 199816 168
rect 199496 88 199508 144
rect 199564 88 199588 144
rect 199644 88 199668 144
rect 199724 88 199748 144
rect 199804 88 199816 144
rect 205100 134 205128 2382
rect 207940 2304 207992 2310
rect 207940 2246 207992 2252
rect 207952 202 207980 2246
rect 208228 1358 208256 2746
rect 208596 2746 208716 2774
rect 208596 2650 208624 2746
rect 208584 2644 208636 2650
rect 208584 2586 208636 2592
rect 208596 2446 208624 2586
rect 210252 2446 210280 2790
rect 210528 2650 210556 3062
rect 211816 2774 211844 11222
rect 212092 11014 212120 11342
rect 212724 11280 212776 11286
rect 212724 11222 212776 11228
rect 212080 11008 212132 11014
rect 212080 10950 212132 10956
rect 212172 11008 212224 11014
rect 212172 10950 212224 10956
rect 212184 10742 212212 10950
rect 212356 10804 212408 10810
rect 212356 10746 212408 10752
rect 212172 10736 212224 10742
rect 212172 10678 212224 10684
rect 212368 10334 212396 10746
rect 212736 10606 212764 11222
rect 213656 11150 213684 11455
rect 214432 11455 214434 11464
rect 258632 11484 258684 11490
rect 214380 11426 214432 11432
rect 258632 11426 258684 11432
rect 258540 11416 258592 11422
rect 258540 11358 258592 11364
rect 219256 11348 219308 11354
rect 219256 11290 219308 11296
rect 254216 11348 254268 11354
rect 254216 11290 254268 11296
rect 213828 11280 213880 11286
rect 213748 11240 213828 11268
rect 213644 11144 213696 11150
rect 213644 11086 213696 11092
rect 212724 10600 212776 10606
rect 212724 10542 212776 10548
rect 213276 10600 213328 10606
rect 213276 10542 213328 10548
rect 212356 10328 212408 10334
rect 212356 10270 212408 10276
rect 212448 10328 212500 10334
rect 212448 10270 212500 10276
rect 212460 8906 212488 10270
rect 212540 9512 212592 9518
rect 212540 9454 212592 9460
rect 212448 8900 212500 8906
rect 212448 8842 212500 8848
rect 212552 3058 212580 9454
rect 212540 3052 212592 3058
rect 212540 2994 212592 3000
rect 211816 2746 212120 2774
rect 210516 2644 210568 2650
rect 210516 2586 210568 2592
rect 208584 2440 208636 2446
rect 208584 2382 208636 2388
rect 210240 2440 210292 2446
rect 210240 2382 210292 2388
rect 208216 1352 208268 1358
rect 208216 1294 208268 1300
rect 210252 270 210280 2382
rect 212092 814 212120 2746
rect 213288 2446 213316 10542
rect 213276 2440 213328 2446
rect 213276 2382 213328 2388
rect 213092 2304 213144 2310
rect 213092 2246 213144 2252
rect 213104 1222 213132 2246
rect 213092 1216 213144 1222
rect 213092 1158 213144 1164
rect 212080 808 212132 814
rect 212080 750 212132 756
rect 213748 513 213776 11240
rect 213828 11222 213880 11228
rect 213920 11280 213972 11286
rect 213920 11222 213972 11228
rect 215392 11280 215444 11286
rect 215392 11222 215444 11228
rect 215576 11280 215628 11286
rect 215576 11222 215628 11228
rect 217048 11280 217100 11286
rect 217048 11222 217100 11228
rect 217232 11280 217284 11286
rect 217232 11222 217284 11228
rect 217600 11280 217652 11286
rect 217600 11222 217652 11228
rect 218336 11280 218388 11286
rect 218336 11222 218388 11228
rect 213932 10266 213960 11222
rect 214012 11144 214064 11150
rect 214012 11086 214064 11092
rect 213920 10260 213972 10266
rect 213920 10202 213972 10208
rect 214024 9994 214052 11086
rect 214104 10260 214156 10266
rect 214104 10202 214156 10208
rect 214116 10169 214144 10202
rect 214102 10160 214158 10169
rect 214102 10095 214158 10104
rect 214012 9988 214064 9994
rect 214012 9930 214064 9936
rect 213828 9920 213880 9926
rect 213828 9862 213880 9868
rect 213840 9586 213868 9862
rect 213828 9580 213880 9586
rect 213828 9522 213880 9528
rect 215404 9178 215432 11222
rect 215392 9172 215444 9178
rect 215392 9114 215444 9120
rect 215588 8537 215616 11222
rect 216772 11144 216824 11150
rect 216772 11086 216824 11092
rect 216784 10946 216812 11086
rect 216772 10940 216824 10946
rect 216772 10882 216824 10888
rect 215574 8528 215630 8537
rect 215574 8463 215630 8472
rect 215392 2848 215444 2854
rect 215392 2790 215444 2796
rect 215404 2446 215432 2790
rect 217060 2774 217088 11222
rect 217244 10062 217272 11222
rect 217612 10334 217640 11222
rect 217876 10532 217928 10538
rect 217876 10474 217928 10480
rect 217888 10334 217916 10474
rect 217600 10328 217652 10334
rect 217600 10270 217652 10276
rect 217876 10328 217928 10334
rect 217876 10270 217928 10276
rect 217232 10056 217284 10062
rect 217232 9998 217284 10004
rect 217968 9512 218020 9518
rect 217968 9454 218020 9460
rect 217980 9110 218008 9454
rect 217968 9104 218020 9110
rect 217968 9046 218020 9052
rect 218348 7274 218376 11222
rect 218796 10532 218848 10538
rect 218796 10474 218848 10480
rect 218428 9988 218480 9994
rect 218428 9930 218480 9936
rect 218336 7268 218388 7274
rect 218336 7210 218388 7216
rect 216968 2746 217088 2774
rect 215392 2440 215444 2446
rect 215392 2382 215444 2388
rect 215404 1154 215432 2382
rect 215668 2304 215720 2310
rect 215668 2246 215720 2252
rect 215680 1970 215708 2246
rect 215668 1964 215720 1970
rect 215668 1906 215720 1912
rect 216968 1329 216996 2746
rect 218440 2446 218468 9930
rect 218808 9654 218836 10474
rect 218796 9648 218848 9654
rect 218796 9590 218848 9596
rect 219268 2774 219296 11290
rect 219440 11280 219492 11286
rect 219440 11222 219492 11228
rect 220360 11280 220412 11286
rect 220360 11222 220412 11228
rect 220912 11280 220964 11286
rect 220912 11222 220964 11228
rect 221648 11280 221700 11286
rect 221648 11222 221700 11228
rect 222200 11280 222252 11286
rect 222200 11222 222252 11228
rect 222476 11280 222528 11286
rect 222476 11222 222528 11228
rect 223212 11280 223264 11286
rect 223212 11222 223264 11228
rect 223764 11280 223816 11286
rect 223764 11222 223816 11228
rect 224960 11280 225012 11286
rect 224960 11222 225012 11228
rect 225420 11280 225472 11286
rect 225420 11222 225472 11228
rect 225788 11280 225840 11286
rect 225788 11222 225840 11228
rect 226432 11280 226484 11286
rect 226432 11222 226484 11228
rect 226984 11280 227036 11286
rect 226984 11222 227036 11228
rect 227352 11280 227404 11286
rect 227352 11222 227404 11228
rect 228088 11280 228140 11286
rect 228088 11222 228140 11228
rect 228456 11280 228508 11286
rect 228456 11222 228508 11228
rect 229192 11280 229244 11286
rect 229192 11222 229244 11228
rect 229836 11280 229888 11286
rect 229836 11222 229888 11228
rect 230388 11280 230440 11286
rect 230388 11222 230440 11228
rect 230848 11280 230900 11286
rect 230848 11222 230900 11228
rect 231400 11280 231452 11286
rect 231400 11222 231452 11228
rect 231860 11280 231912 11286
rect 231860 11222 231912 11228
rect 232320 11280 232372 11286
rect 232320 11222 232372 11228
rect 233424 11280 233476 11286
rect 233424 11222 233476 11228
rect 233608 11280 233660 11286
rect 233608 11222 233660 11228
rect 233884 11280 233936 11286
rect 233884 11222 233936 11228
rect 234712 11280 234764 11286
rect 234712 11222 234764 11228
rect 234988 11280 235040 11286
rect 234988 11222 235040 11228
rect 235724 11280 235776 11286
rect 235724 11222 235776 11228
rect 236276 11280 236328 11286
rect 236276 11222 236328 11228
rect 236920 11280 236972 11286
rect 236920 11222 236972 11228
rect 237380 11280 237432 11286
rect 237380 11222 237432 11228
rect 237932 11280 237984 11286
rect 237932 11222 237984 11228
rect 238300 11280 238352 11286
rect 238300 11222 238352 11228
rect 238944 11280 238996 11286
rect 238944 11222 238996 11228
rect 239496 11280 239548 11286
rect 239496 11222 239548 11228
rect 240140 11280 240192 11286
rect 240140 11222 240192 11228
rect 240416 11280 240468 11286
rect 240416 11222 240468 11228
rect 241152 11280 241204 11286
rect 241152 11222 241204 11228
rect 241612 11280 241664 11286
rect 241612 11222 241664 11228
rect 242900 11280 242952 11286
rect 242900 11222 242952 11228
rect 243360 11280 243412 11286
rect 243360 11222 243412 11228
rect 244464 11280 244516 11286
rect 244464 11222 244516 11228
rect 245016 11280 245068 11286
rect 245016 11222 245068 11228
rect 245384 11280 245436 11286
rect 245384 11222 245436 11228
rect 246120 11280 246172 11286
rect 246120 11222 246172 11228
rect 246672 11280 246724 11286
rect 246672 11222 246724 11228
rect 246948 11280 247000 11286
rect 246948 11222 247000 11228
rect 247684 11280 247736 11286
rect 247684 11222 247736 11228
rect 248604 11280 248656 11286
rect 248604 11222 248656 11228
rect 249340 11280 249392 11286
rect 249340 11222 249392 11228
rect 249984 11280 250036 11286
rect 249984 11222 250036 11228
rect 250260 11280 250312 11286
rect 250260 11222 250312 11228
rect 251548 11280 251600 11286
rect 251548 11222 251600 11228
rect 251916 11280 251968 11286
rect 251916 11222 251968 11228
rect 252744 11280 252796 11286
rect 252744 11222 252796 11228
rect 253112 11280 253164 11286
rect 253112 11222 253164 11228
rect 254032 11280 254084 11286
rect 254032 11222 254084 11228
rect 219452 10742 219480 11222
rect 219900 11212 219952 11218
rect 219900 11154 219952 11160
rect 219440 10736 219492 10742
rect 219440 10678 219492 10684
rect 219912 8634 219940 11154
rect 220176 10872 220228 10878
rect 220176 10814 220228 10820
rect 220084 10736 220136 10742
rect 220084 10678 220136 10684
rect 219992 10600 220044 10606
rect 219992 10542 220044 10548
rect 220004 10062 220032 10542
rect 220096 10402 220124 10678
rect 220188 10402 220216 10814
rect 220084 10396 220136 10402
rect 220084 10338 220136 10344
rect 220176 10396 220228 10402
rect 220176 10338 220228 10344
rect 219992 10056 220044 10062
rect 219992 9998 220044 10004
rect 220372 9518 220400 11222
rect 220924 10334 220952 11222
rect 221372 10872 221424 10878
rect 221372 10814 221424 10820
rect 220912 10328 220964 10334
rect 220912 10270 220964 10276
rect 221384 9654 221412 10814
rect 221372 9648 221424 9654
rect 221372 9590 221424 9596
rect 220360 9512 220412 9518
rect 220360 9454 220412 9460
rect 220544 9512 220596 9518
rect 220544 9454 220596 9460
rect 219900 8628 219952 8634
rect 219900 8570 219952 8576
rect 220556 3466 220584 9454
rect 221660 8090 221688 11222
rect 221648 8084 221700 8090
rect 221648 8026 221700 8032
rect 222212 6633 222240 11222
rect 222488 8498 222516 11222
rect 222476 8492 222528 8498
rect 222476 8434 222528 8440
rect 223224 6798 223252 11222
rect 223212 6792 223264 6798
rect 223212 6734 223264 6740
rect 222198 6624 222254 6633
rect 222198 6559 222254 6568
rect 223776 5642 223804 11222
rect 224776 11144 224828 11150
rect 224776 11086 224828 11092
rect 224788 11014 224816 11086
rect 224776 11008 224828 11014
rect 224776 10950 224828 10956
rect 224684 9512 224736 9518
rect 224684 9454 224736 9460
rect 224132 8900 224184 8906
rect 224132 8842 224184 8848
rect 223764 5636 223816 5642
rect 223764 5578 223816 5584
rect 220544 3460 220596 3466
rect 220544 3402 220596 3408
rect 220544 2848 220596 2854
rect 220544 2790 220596 2796
rect 219176 2746 219296 2774
rect 218428 2440 218480 2446
rect 218428 2382 218480 2388
rect 218244 2304 218296 2310
rect 218244 2246 218296 2252
rect 216954 1320 217010 1329
rect 216954 1255 217010 1264
rect 215392 1148 215444 1154
rect 215392 1090 215444 1096
rect 218256 1018 218284 2246
rect 219176 1193 219204 2746
rect 220556 2446 220584 2790
rect 224144 2650 224172 8842
rect 224696 8401 224724 9454
rect 224682 8392 224738 8401
rect 224682 8327 224738 8336
rect 224972 6866 225000 11222
rect 225052 10804 225104 10810
rect 225052 10746 225104 10752
rect 225064 10690 225092 10746
rect 225064 10662 225184 10690
rect 225156 10606 225184 10662
rect 225144 10600 225196 10606
rect 225144 10542 225196 10548
rect 224960 6860 225012 6866
rect 224960 6802 225012 6808
rect 225432 6730 225460 11222
rect 225800 10198 225828 11222
rect 225788 10192 225840 10198
rect 225788 10134 225840 10140
rect 226444 7206 226472 11222
rect 226892 11144 226944 11150
rect 226892 11086 226944 11092
rect 226904 10878 226932 11086
rect 226892 10872 226944 10878
rect 226892 10814 226944 10820
rect 226432 7200 226484 7206
rect 226432 7142 226484 7148
rect 225420 6724 225472 6730
rect 225420 6666 225472 6672
rect 226996 5778 227024 11222
rect 227364 10130 227392 11222
rect 227352 10124 227404 10130
rect 227352 10066 227404 10072
rect 228100 5846 228128 11222
rect 228272 9512 228324 9518
rect 228272 9454 228324 9460
rect 228088 5840 228140 5846
rect 228088 5782 228140 5788
rect 226984 5772 227036 5778
rect 226984 5714 227036 5720
rect 226064 2848 226116 2854
rect 228284 2825 228312 9454
rect 228468 7954 228496 11222
rect 229100 9580 229152 9586
rect 229100 9522 229152 9528
rect 229112 9382 229140 9522
rect 229100 9376 229152 9382
rect 229100 9318 229152 9324
rect 229112 9110 229140 9318
rect 229100 9104 229152 9110
rect 229100 9046 229152 9052
rect 229204 8974 229232 11222
rect 229284 11076 229336 11082
rect 229284 11018 229336 11024
rect 229192 8968 229244 8974
rect 229192 8910 229244 8916
rect 228456 7948 228508 7954
rect 228456 7890 228508 7896
rect 226064 2790 226116 2796
rect 228270 2816 228326 2825
rect 224132 2644 224184 2650
rect 224132 2586 224184 2592
rect 224144 2446 224172 2586
rect 220544 2440 220596 2446
rect 220544 2382 220596 2388
rect 224132 2440 224184 2446
rect 224132 2382 224184 2388
rect 219624 1352 219676 1358
rect 219624 1294 219676 1300
rect 219162 1184 219218 1193
rect 219162 1119 219218 1128
rect 218244 1012 218296 1018
rect 218244 954 218296 960
rect 219532 944 219584 950
rect 219532 886 219584 892
rect 219544 678 219572 886
rect 219636 882 219664 1294
rect 219716 1148 219768 1154
rect 219716 1090 219768 1096
rect 219624 876 219676 882
rect 219624 818 219676 824
rect 219532 672 219584 678
rect 219532 614 219584 620
rect 213734 504 213790 513
rect 213734 439 213790 448
rect 210240 264 210292 270
rect 210240 206 210292 212
rect 207940 196 207992 202
rect 207940 138 207992 144
rect 199496 64 199816 88
rect 205088 128 205140 134
rect 205088 70 205140 76
rect 219728 66 219756 1090
rect 220556 1086 220584 2382
rect 226076 2378 226104 2790
rect 229296 2774 229324 11018
rect 229652 11008 229704 11014
rect 229652 10950 229704 10956
rect 229664 9926 229692 10950
rect 229744 10872 229796 10878
rect 229744 10814 229796 10820
rect 229756 10538 229784 10814
rect 229744 10532 229796 10538
rect 229744 10474 229796 10480
rect 229652 9920 229704 9926
rect 229652 9862 229704 9868
rect 229848 6322 229876 11222
rect 230400 8514 230428 11222
rect 230860 10402 230888 11222
rect 230848 10396 230900 10402
rect 230848 10338 230900 10344
rect 230400 8486 230520 8514
rect 230492 6662 230520 8486
rect 230480 6656 230532 6662
rect 230480 6598 230532 6604
rect 229836 6316 229888 6322
rect 229836 6258 229888 6264
rect 231412 6186 231440 11222
rect 231872 6390 231900 11222
rect 232044 9512 232096 9518
rect 232044 9454 232096 9460
rect 231860 6384 231912 6390
rect 231860 6326 231912 6332
rect 231400 6180 231452 6186
rect 231400 6122 231452 6128
rect 228270 2751 228326 2760
rect 229204 2746 229324 2774
rect 229204 2650 229232 2746
rect 229192 2644 229244 2650
rect 229192 2586 229244 2592
rect 231860 2644 231912 2650
rect 231860 2586 231912 2592
rect 229204 2446 229232 2586
rect 231872 2446 231900 2586
rect 229192 2440 229244 2446
rect 229192 2382 229244 2388
rect 231860 2440 231912 2446
rect 231860 2382 231912 2388
rect 226064 2372 226116 2378
rect 226064 2314 226116 2320
rect 220820 2304 220872 2310
rect 220820 2246 220872 2252
rect 223396 2304 223448 2310
rect 223396 2246 223448 2252
rect 225972 2304 226024 2310
rect 225972 2246 226024 2252
rect 220832 1902 220860 2246
rect 220820 1896 220872 1902
rect 220820 1838 220872 1844
rect 223408 1154 223436 2246
rect 225984 1834 226012 2246
rect 225972 1828 226024 1834
rect 225972 1770 226024 1776
rect 226076 1358 226104 2314
rect 228548 2304 228600 2310
rect 228548 2246 228600 2252
rect 229100 2304 229152 2310
rect 229100 2246 229152 2252
rect 226064 1352 226116 1358
rect 226064 1294 226116 1300
rect 228456 1352 228508 1358
rect 228456 1294 228508 1300
rect 224316 1216 224368 1222
rect 224316 1158 224368 1164
rect 226432 1216 226484 1222
rect 226432 1158 226484 1164
rect 223396 1148 223448 1154
rect 223396 1090 223448 1096
rect 220544 1080 220596 1086
rect 220544 1022 220596 1028
rect 222108 1080 222160 1086
rect 222108 1022 222160 1028
rect 222120 814 222148 1022
rect 224328 814 224356 1158
rect 226444 814 226472 1158
rect 228468 814 228496 1294
rect 228560 1018 228588 2246
rect 229112 1086 229140 2246
rect 232056 2009 232084 9454
rect 232332 9450 232360 11222
rect 232320 9444 232372 9450
rect 232320 9386 232372 9392
rect 232872 9172 232924 9178
rect 232872 9114 232924 9120
rect 232884 2650 232912 9114
rect 233436 6361 233464 11222
rect 233422 6352 233478 6361
rect 233422 6287 233478 6296
rect 233620 5166 233648 11222
rect 233896 8430 233924 11222
rect 234436 9580 234488 9586
rect 234436 9522 234488 9528
rect 233884 8424 233936 8430
rect 233884 8366 233936 8372
rect 233608 5160 233660 5166
rect 233608 5102 233660 5108
rect 234448 2650 234476 9522
rect 234724 4214 234752 11222
rect 235000 7750 235028 11222
rect 235736 10946 235764 11222
rect 235724 10940 235776 10946
rect 235724 10882 235776 10888
rect 236000 9512 236052 9518
rect 236000 9454 236052 9460
rect 234988 7744 235040 7750
rect 234988 7686 235040 7692
rect 234712 4208 234764 4214
rect 234712 4150 234764 4156
rect 236012 3398 236040 9454
rect 236288 6254 236316 11222
rect 236644 11076 236696 11082
rect 236644 11018 236696 11024
rect 236656 10946 236684 11018
rect 236644 10940 236696 10946
rect 236644 10882 236696 10888
rect 236828 9512 236880 9518
rect 236828 9454 236880 9460
rect 236840 8974 236868 9454
rect 236828 8968 236880 8974
rect 236828 8910 236880 8916
rect 236276 6248 236328 6254
rect 236276 6190 236328 6196
rect 236932 5302 236960 11222
rect 237392 8566 237420 11222
rect 237380 8560 237432 8566
rect 237380 8502 237432 8508
rect 237012 7540 237064 7546
rect 237012 7482 237064 7488
rect 236920 5296 236972 5302
rect 236920 5238 236972 5244
rect 236000 3392 236052 3398
rect 236000 3334 236052 3340
rect 237024 2650 237052 7482
rect 237944 5098 237972 11222
rect 238312 6225 238340 11222
rect 238852 10804 238904 10810
rect 238852 10746 238904 10752
rect 238864 10538 238892 10746
rect 238956 10606 238984 11222
rect 239404 11076 239456 11082
rect 239404 11018 239456 11024
rect 239220 11008 239272 11014
rect 239416 10962 239444 11018
rect 239272 10956 239444 10962
rect 239220 10950 239444 10956
rect 239232 10934 239444 10950
rect 239404 10872 239456 10878
rect 239404 10814 239456 10820
rect 239416 10606 239444 10814
rect 238944 10600 238996 10606
rect 238944 10542 238996 10548
rect 239404 10600 239456 10606
rect 239404 10542 239456 10548
rect 238852 10532 238904 10538
rect 238852 10474 238904 10480
rect 239036 10396 239088 10402
rect 239036 10338 239088 10344
rect 238298 6216 238354 6225
rect 238298 6151 238354 6160
rect 237932 5092 237984 5098
rect 237932 5034 237984 5040
rect 232872 2644 232924 2650
rect 232872 2586 232924 2592
rect 234436 2644 234488 2650
rect 234436 2586 234488 2592
rect 237012 2644 237064 2650
rect 237012 2586 237064 2592
rect 234448 2446 234476 2586
rect 237024 2446 237052 2586
rect 239048 2446 239076 10338
rect 239508 7818 239536 11222
rect 239956 9580 240008 9586
rect 239956 9522 240008 9528
rect 239680 9512 239732 9518
rect 239680 9454 239732 9460
rect 239692 9042 239720 9454
rect 239968 9042 239996 9522
rect 239680 9036 239732 9042
rect 239680 8978 239732 8984
rect 239956 9036 240008 9042
rect 239956 8978 240008 8984
rect 239496 7812 239548 7818
rect 239496 7754 239548 7760
rect 240152 4729 240180 11222
rect 240428 10470 240456 11222
rect 240416 10464 240468 10470
rect 240416 10406 240468 10412
rect 241164 5370 241192 11222
rect 241520 10464 241572 10470
rect 241520 10406 241572 10412
rect 241532 9382 241560 10406
rect 241520 9376 241572 9382
rect 241520 9318 241572 9324
rect 241624 6118 241652 11222
rect 242164 8560 242216 8566
rect 242164 8502 242216 8508
rect 241612 6112 241664 6118
rect 241612 6054 241664 6060
rect 241152 5364 241204 5370
rect 241152 5306 241204 5312
rect 240138 4720 240194 4729
rect 240138 4655 240194 4664
rect 242176 2650 242204 8502
rect 242912 6089 242940 11222
rect 242898 6080 242954 6089
rect 242898 6015 242954 6024
rect 243372 4826 243400 11222
rect 244004 9580 244056 9586
rect 244004 9522 244056 9528
rect 243728 9512 243780 9518
rect 243728 9454 243780 9460
rect 243360 4820 243412 4826
rect 243360 4762 243412 4768
rect 243740 3534 243768 9454
rect 244016 9382 244044 9522
rect 244004 9376 244056 9382
rect 244004 9318 244056 9324
rect 244476 4554 244504 11222
rect 244464 4548 244516 4554
rect 244464 4490 244516 4496
rect 244832 4548 244884 4554
rect 244832 4490 244884 4496
rect 243728 3528 243780 3534
rect 243728 3470 243780 3476
rect 244844 2650 244872 4490
rect 245028 4457 245056 11222
rect 245396 10606 245424 11222
rect 245384 10600 245436 10606
rect 245384 10542 245436 10548
rect 246132 8022 246160 11222
rect 246120 8016 246172 8022
rect 246120 7958 246172 7964
rect 246684 4690 246712 11222
rect 246960 10538 246988 11222
rect 246948 10532 247000 10538
rect 246948 10474 247000 10480
rect 247224 10532 247276 10538
rect 247224 10474 247276 10480
rect 246672 4684 246724 4690
rect 246672 4626 246724 4632
rect 245014 4448 245070 4457
rect 245014 4383 245070 4392
rect 247236 2650 247264 10474
rect 247696 4758 247724 11222
rect 248512 11144 248564 11150
rect 248512 11086 248564 11092
rect 248524 5409 248552 11086
rect 248616 9654 248644 11222
rect 248696 10940 248748 10946
rect 248696 10882 248748 10888
rect 249064 10940 249116 10946
rect 249064 10882 249116 10888
rect 248708 10810 248736 10882
rect 248696 10804 248748 10810
rect 248696 10746 248748 10752
rect 249076 10402 249104 10882
rect 249064 10396 249116 10402
rect 249064 10338 249116 10344
rect 248604 9648 248656 9654
rect 248604 9590 248656 9596
rect 248510 5400 248566 5409
rect 248510 5335 248566 5344
rect 247684 4752 247736 4758
rect 247684 4694 247736 4700
rect 249352 4282 249380 11222
rect 249524 7200 249576 7206
rect 249524 7142 249576 7148
rect 249340 4276 249392 4282
rect 249340 4218 249392 4224
rect 242164 2644 242216 2650
rect 242164 2586 242216 2592
rect 244832 2644 244884 2650
rect 244832 2586 244884 2592
rect 247224 2644 247276 2650
rect 247224 2586 247276 2592
rect 242176 2446 242204 2586
rect 244844 2446 244872 2586
rect 247236 2446 247264 2586
rect 234436 2440 234488 2446
rect 234436 2382 234488 2388
rect 237012 2440 237064 2446
rect 237012 2382 237064 2388
rect 239036 2440 239088 2446
rect 239036 2382 239088 2388
rect 242164 2440 242216 2446
rect 242164 2382 242216 2388
rect 244832 2440 244884 2446
rect 244832 2382 244884 2388
rect 247224 2440 247276 2446
rect 247224 2382 247276 2388
rect 233240 2372 233292 2378
rect 233240 2314 233292 2320
rect 243912 2372 243964 2378
rect 243912 2314 243964 2320
rect 232042 2000 232098 2009
rect 232042 1935 232098 1944
rect 233252 1358 233280 2314
rect 233700 2304 233752 2310
rect 233700 2246 233752 2252
rect 236276 2304 236328 2310
rect 236276 2246 236328 2252
rect 241428 2304 241480 2310
rect 241428 2246 241480 2252
rect 242900 2304 242952 2310
rect 242900 2246 242952 2252
rect 233240 1352 233292 1358
rect 233240 1294 233292 1300
rect 230572 1148 230624 1154
rect 230572 1090 230624 1096
rect 229100 1080 229152 1086
rect 229100 1022 229152 1028
rect 228548 1012 228600 1018
rect 228548 954 228600 960
rect 230584 814 230612 1090
rect 233712 1086 233740 2246
rect 234988 1352 235040 1358
rect 234988 1294 235040 1300
rect 233700 1080 233752 1086
rect 233700 1022 233752 1028
rect 231676 1012 231728 1018
rect 231676 954 231728 960
rect 231688 814 231716 954
rect 235000 814 235028 1294
rect 236288 1222 236316 2246
rect 236276 1216 236328 1222
rect 236276 1158 236328 1164
rect 238484 1216 238536 1222
rect 238484 1158 238536 1164
rect 237288 1148 237340 1154
rect 237288 1090 237340 1096
rect 237300 814 237328 1090
rect 238496 814 238524 1158
rect 241440 1086 241468 2246
rect 242912 1086 242940 2246
rect 243924 1222 243952 2314
rect 244096 2304 244148 2310
rect 244016 2264 244096 2292
rect 244016 1358 244044 2264
rect 244096 2246 244148 2252
rect 247040 2304 247092 2310
rect 247040 2246 247092 2252
rect 244004 1352 244056 1358
rect 244004 1294 244056 1300
rect 244096 1284 244148 1290
rect 244372 1284 244424 1290
rect 244148 1244 244372 1272
rect 244096 1226 244148 1232
rect 244372 1226 244424 1232
rect 243912 1216 243964 1222
rect 244648 1216 244700 1222
rect 243912 1158 243964 1164
rect 244384 1164 244648 1170
rect 244384 1158 244700 1164
rect 244384 1142 244688 1158
rect 245752 1148 245804 1154
rect 244384 1086 244412 1142
rect 245752 1090 245804 1096
rect 241428 1080 241480 1086
rect 241428 1022 241480 1028
rect 241520 1080 241572 1086
rect 242900 1080 242952 1086
rect 241520 1022 241572 1028
rect 239404 1012 239456 1018
rect 239404 954 239456 960
rect 239128 944 239180 950
rect 239416 898 239444 954
rect 239180 892 239444 898
rect 239128 886 239444 892
rect 239956 944 240008 950
rect 239956 886 240008 892
rect 239140 870 239444 886
rect 222108 808 222160 814
rect 222108 750 222160 756
rect 224316 808 224368 814
rect 224316 750 224368 756
rect 226432 808 226484 814
rect 226432 750 226484 756
rect 228456 808 228508 814
rect 228456 750 228508 756
rect 230572 808 230624 814
rect 230572 750 230624 756
rect 231676 808 231728 814
rect 231676 750 231728 756
rect 234988 808 235040 814
rect 234988 750 235040 756
rect 237288 808 237340 814
rect 237288 750 237340 756
rect 238484 808 238536 814
rect 238484 750 238536 756
rect 239968 746 239996 886
rect 241532 746 241560 1022
rect 241624 1006 242020 1034
rect 242900 1022 242952 1028
rect 242992 1080 243044 1086
rect 242992 1022 243044 1028
rect 244372 1080 244424 1086
rect 244372 1022 244424 1028
rect 241624 950 241652 1006
rect 241612 944 241664 950
rect 241612 886 241664 892
rect 241704 944 241756 950
rect 241704 886 241756 892
rect 241716 814 241744 886
rect 241992 882 242020 1006
rect 241980 876 242032 882
rect 241980 818 242032 824
rect 243004 814 243032 1022
rect 245764 950 245792 1090
rect 247052 1086 247080 2246
rect 249536 1426 249564 7142
rect 249892 4480 249944 4486
rect 249892 4422 249944 4428
rect 249904 2650 249932 4422
rect 249996 2990 250024 11222
rect 250272 9110 250300 11222
rect 251272 11144 251324 11150
rect 251272 11086 251324 11092
rect 251180 10736 251232 10742
rect 251180 10678 251232 10684
rect 250812 10600 250864 10606
rect 250812 10542 250864 10548
rect 250260 9104 250312 9110
rect 250260 9046 250312 9052
rect 250824 7478 250852 10542
rect 251192 9042 251220 10678
rect 251180 9036 251232 9042
rect 251180 8978 251232 8984
rect 250812 7472 250864 7478
rect 250812 7414 250864 7420
rect 251284 4078 251312 11086
rect 251456 7744 251508 7750
rect 251456 7686 251508 7692
rect 251468 7410 251496 7686
rect 251456 7404 251508 7410
rect 251456 7346 251508 7352
rect 251364 6724 251416 6730
rect 251364 6666 251416 6672
rect 251272 4072 251324 4078
rect 251272 4014 251324 4020
rect 249984 2984 250036 2990
rect 249984 2926 250036 2932
rect 249892 2644 249944 2650
rect 249892 2586 249944 2592
rect 249904 2446 249932 2586
rect 249892 2440 249944 2446
rect 249892 2382 249944 2388
rect 251376 1737 251404 6666
rect 251468 1873 251496 7346
rect 251560 4321 251588 11222
rect 251928 10470 251956 11222
rect 251916 10464 251968 10470
rect 251916 10406 251968 10412
rect 251916 10328 251968 10334
rect 251916 10270 251968 10276
rect 251546 4312 251602 4321
rect 251546 4247 251602 4256
rect 251928 2446 251956 10270
rect 252468 7744 252520 7750
rect 252468 7686 252520 7692
rect 252480 7410 252508 7686
rect 252468 7404 252520 7410
rect 252468 7346 252520 7352
rect 252008 7336 252060 7342
rect 252008 7278 252060 7284
rect 252020 6934 252048 7278
rect 252008 6928 252060 6934
rect 252008 6870 252060 6876
rect 251916 2440 251968 2446
rect 251916 2382 251968 2388
rect 251454 1864 251510 1873
rect 251454 1799 251510 1808
rect 251362 1728 251418 1737
rect 251362 1663 251418 1672
rect 252480 1630 252508 7346
rect 252560 6656 252612 6662
rect 252560 6598 252612 6604
rect 252572 5370 252600 6598
rect 252652 5636 252704 5642
rect 252652 5578 252704 5584
rect 252560 5364 252612 5370
rect 252560 5306 252612 5312
rect 252664 3126 252692 5578
rect 252756 4593 252784 11222
rect 252742 4584 252798 4593
rect 252742 4519 252798 4528
rect 253124 4010 253152 11222
rect 254044 8974 254072 11222
rect 254032 8968 254084 8974
rect 254032 8910 254084 8916
rect 253940 7404 253992 7410
rect 253940 7346 253992 7352
rect 253952 6662 253980 7346
rect 253940 6656 253992 6662
rect 253940 6598 253992 6604
rect 253112 4004 253164 4010
rect 253112 3946 253164 3952
rect 252652 3120 252704 3126
rect 252652 3062 252704 3068
rect 253952 2514 253980 6598
rect 254228 3194 254256 11290
rect 255320 11280 255372 11286
rect 255320 11222 255372 11228
rect 255872 11280 255924 11286
rect 255872 11222 255924 11228
rect 256424 11280 256476 11286
rect 256424 11222 256476 11228
rect 255228 11076 255280 11082
rect 255228 11018 255280 11024
rect 254952 11008 255004 11014
rect 254952 10950 255004 10956
rect 254584 6656 254636 6662
rect 254584 6598 254636 6604
rect 254216 3188 254268 3194
rect 254216 3130 254268 3136
rect 254596 2553 254624 6598
rect 254582 2544 254638 2553
rect 253940 2508 253992 2514
rect 254582 2479 254638 2488
rect 253940 2450 253992 2456
rect 253848 2304 253900 2310
rect 253848 2246 253900 2252
rect 252468 1624 252520 1630
rect 252468 1566 252520 1572
rect 249524 1420 249576 1426
rect 249524 1362 249576 1368
rect 247592 1284 247644 1290
rect 247592 1226 247644 1232
rect 247040 1080 247092 1086
rect 247040 1022 247092 1028
rect 247604 950 247632 1226
rect 253860 1154 253888 2246
rect 254964 1426 254992 10950
rect 255240 7410 255268 11018
rect 255332 10742 255360 11222
rect 255688 11144 255740 11150
rect 255688 11086 255740 11092
rect 255320 10736 255372 10742
rect 255320 10678 255372 10684
rect 255700 9382 255728 11086
rect 255688 9376 255740 9382
rect 255688 9318 255740 9324
rect 255228 7404 255280 7410
rect 255228 7346 255280 7352
rect 255780 7336 255832 7342
rect 255780 7278 255832 7284
rect 255792 2417 255820 7278
rect 255884 4622 255912 11222
rect 256332 6792 256384 6798
rect 256332 6734 256384 6740
rect 256344 6118 256372 6734
rect 256332 6112 256384 6118
rect 256332 6054 256384 6060
rect 255872 4616 255924 4622
rect 255872 4558 255924 4564
rect 256344 2689 256372 6054
rect 256436 3942 256464 11222
rect 258552 10878 258580 11358
rect 258540 10872 258592 10878
rect 258540 10814 258592 10820
rect 256976 10464 257028 10470
rect 256976 10406 257028 10412
rect 256988 7546 257016 10406
rect 258644 10334 258672 11426
rect 258736 10538 258764 11494
rect 258816 11144 258868 11150
rect 258816 11086 258868 11092
rect 258828 10606 258856 11086
rect 262036 11008 262088 11014
rect 262036 10950 262088 10956
rect 260840 10804 260892 10810
rect 260840 10746 260892 10752
rect 258816 10600 258868 10606
rect 258816 10542 258868 10548
rect 258724 10532 258776 10538
rect 258724 10474 258776 10480
rect 258632 10328 258684 10334
rect 258632 10270 258684 10276
rect 260196 9376 260248 9382
rect 260196 9318 260248 9324
rect 258356 7744 258408 7750
rect 258356 7686 258408 7692
rect 256976 7540 257028 7546
rect 256976 7482 257028 7488
rect 256988 7410 257016 7482
rect 256976 7404 257028 7410
rect 256976 7346 257028 7352
rect 258368 6866 258396 7686
rect 258356 6860 258408 6866
rect 258356 6802 258408 6808
rect 257528 6792 257580 6798
rect 257528 6734 257580 6740
rect 259000 6792 259052 6798
rect 259000 6734 259052 6740
rect 259920 6792 259972 6798
rect 259920 6734 259972 6740
rect 257160 6724 257212 6730
rect 257160 6666 257212 6672
rect 257172 6458 257200 6666
rect 257160 6452 257212 6458
rect 257160 6394 257212 6400
rect 257540 6118 257568 6734
rect 259012 6118 259040 6734
rect 259932 6118 259960 6734
rect 257528 6112 257580 6118
rect 257528 6054 257580 6060
rect 259000 6112 259052 6118
rect 259000 6054 259052 6060
rect 259920 6112 259972 6118
rect 259920 6054 259972 6060
rect 256424 3936 256476 3942
rect 256424 3878 256476 3884
rect 256330 2680 256386 2689
rect 256330 2615 256386 2624
rect 255778 2408 255834 2417
rect 255778 2343 255834 2352
rect 255044 2304 255096 2310
rect 255044 2246 255096 2252
rect 255412 2304 255464 2310
rect 257540 2281 257568 6054
rect 257620 3460 257672 3466
rect 257620 3402 257672 3408
rect 257632 2650 257660 3402
rect 257620 2644 257672 2650
rect 257620 2586 257672 2592
rect 257632 2446 257660 2586
rect 257620 2440 257672 2446
rect 257620 2382 257672 2388
rect 258080 2304 258132 2310
rect 255412 2246 255464 2252
rect 257526 2272 257582 2281
rect 254952 1420 255004 1426
rect 254952 1362 255004 1368
rect 254768 1216 254820 1222
rect 254768 1158 254820 1164
rect 253848 1148 253900 1154
rect 253848 1090 253900 1096
rect 253940 1148 253992 1154
rect 253940 1090 253992 1096
rect 248052 1080 248104 1086
rect 253952 1034 253980 1090
rect 248052 1022 248104 1028
rect 245752 944 245804 950
rect 245752 886 245804 892
rect 246028 944 246080 950
rect 246028 886 246080 892
rect 247592 944 247644 950
rect 247592 886 247644 892
rect 241704 808 241756 814
rect 241704 750 241756 756
rect 242992 808 243044 814
rect 242992 750 243044 756
rect 239956 740 240008 746
rect 239956 682 240008 688
rect 241520 740 241572 746
rect 241520 682 241572 688
rect 246040 678 246068 886
rect 248064 814 248092 1022
rect 253768 1006 253980 1034
rect 253768 950 253796 1006
rect 250812 944 250864 950
rect 250812 886 250864 892
rect 253756 944 253808 950
rect 253756 886 253808 892
rect 248052 808 248104 814
rect 248052 750 248104 756
rect 250824 678 250852 886
rect 254124 876 254176 882
rect 254124 818 254176 824
rect 246028 672 246080 678
rect 246028 614 246080 620
rect 250812 672 250864 678
rect 250812 614 250864 620
rect 254136 513 254164 818
rect 254780 678 254808 1158
rect 255056 1086 255084 2246
rect 255424 1290 255452 2246
rect 258080 2246 258132 2252
rect 257526 2207 257582 2216
rect 258092 1358 258120 2246
rect 259012 2145 259040 6054
rect 258998 2136 259054 2145
rect 258998 2071 259054 2080
rect 259932 1562 259960 6054
rect 260208 2650 260236 9318
rect 260852 7410 260880 10746
rect 262048 7546 262076 10950
rect 267096 10940 267148 10946
rect 267096 10882 267148 10888
rect 262404 9920 262456 9926
rect 262404 9862 262456 9868
rect 262036 7540 262088 7546
rect 262036 7482 262088 7488
rect 262048 7410 262076 7482
rect 260840 7404 260892 7410
rect 260840 7346 260892 7352
rect 262036 7404 262088 7410
rect 262036 7346 262088 7352
rect 262220 6996 262272 7002
rect 262220 6938 262272 6944
rect 262232 6458 262260 6938
rect 262220 6452 262272 6458
rect 262220 6394 262272 6400
rect 260840 6316 260892 6322
rect 260840 6258 260892 6264
rect 262312 6316 262364 6322
rect 262312 6258 262364 6264
rect 260852 6118 260880 6258
rect 262220 6248 262272 6254
rect 262220 6190 262272 6196
rect 260840 6112 260892 6118
rect 260840 6054 260892 6060
rect 260196 2644 260248 2650
rect 260196 2586 260248 2592
rect 260208 2446 260236 2586
rect 260852 2582 260880 6054
rect 260840 2576 260892 2582
rect 260840 2518 260892 2524
rect 262232 2446 262260 6190
rect 262324 5574 262352 6258
rect 262416 6254 262444 9862
rect 265348 9104 265400 9110
rect 265348 9046 265400 9052
rect 264980 7336 265032 7342
rect 264980 7278 265032 7284
rect 264336 6316 264388 6322
rect 264336 6258 264388 6264
rect 262404 6248 262456 6254
rect 262404 6190 262456 6196
rect 264348 6118 264376 6258
rect 264336 6112 264388 6118
rect 264336 6054 264388 6060
rect 263140 5704 263192 5710
rect 263140 5646 263192 5652
rect 263152 5574 263180 5646
rect 262312 5568 262364 5574
rect 262312 5510 262364 5516
rect 263140 5568 263192 5574
rect 263140 5510 263192 5516
rect 260196 2440 260248 2446
rect 260196 2382 260248 2388
rect 262220 2440 262272 2446
rect 262220 2382 262272 2388
rect 260840 2304 260892 2310
rect 260840 2246 260892 2252
rect 259920 1556 259972 1562
rect 259920 1498 259972 1504
rect 258080 1352 258132 1358
rect 258080 1294 258132 1300
rect 258908 1352 258960 1358
rect 258908 1294 258960 1300
rect 255412 1284 255464 1290
rect 255412 1226 255464 1232
rect 256884 1284 256936 1290
rect 256884 1226 256936 1232
rect 254952 1080 255004 1086
rect 254952 1022 255004 1028
rect 255044 1080 255096 1086
rect 255044 1022 255096 1028
rect 254768 672 254820 678
rect 254768 614 254820 620
rect 254964 513 254992 1022
rect 256896 814 256924 1226
rect 258920 814 258948 1294
rect 256884 808 256936 814
rect 256884 750 256936 756
rect 258908 808 258960 814
rect 258908 750 258960 756
rect 252558 504 252614 513
rect 252558 439 252614 448
rect 254122 504 254178 513
rect 254122 439 254178 448
rect 254950 504 255006 513
rect 254950 439 255006 448
rect 259366 504 259422 513
rect 260852 474 260880 2246
rect 262324 1494 262352 5510
rect 263152 2106 263180 5510
rect 263416 2508 263468 2514
rect 263416 2450 263468 2456
rect 263140 2100 263192 2106
rect 263140 2042 263192 2048
rect 262404 1624 262456 1630
rect 262404 1566 262456 1572
rect 262312 1488 262364 1494
rect 262312 1430 262364 1436
rect 261208 1420 261260 1426
rect 261208 1362 261260 1368
rect 261220 1086 261248 1362
rect 261208 1080 261260 1086
rect 261208 1022 261260 1028
rect 261300 1080 261352 1086
rect 261300 1022 261352 1028
rect 261312 814 261340 1022
rect 262416 1018 262444 1566
rect 263428 1358 263456 2450
rect 263600 2304 263652 2310
rect 263600 2246 263652 2252
rect 263416 1352 263468 1358
rect 263416 1294 263468 1300
rect 262404 1012 262456 1018
rect 262404 954 262456 960
rect 262496 1012 262548 1018
rect 262496 954 262548 960
rect 262508 814 262536 954
rect 261300 808 261352 814
rect 261300 750 261352 756
rect 262496 808 262548 814
rect 262496 750 262548 756
rect 263416 808 263468 814
rect 263416 750 263468 756
rect 259366 439 259368 448
rect 252572 270 252600 439
rect 259420 439 259422 448
rect 260840 468 260892 474
rect 259368 410 259420 416
rect 260840 410 260892 416
rect 250628 264 250680 270
rect 250364 212 250628 218
rect 250364 206 250680 212
rect 252560 264 252612 270
rect 252560 206 252612 212
rect 263428 218 263456 750
rect 263612 218 263640 2246
rect 264348 2038 264376 6054
rect 264336 2032 264388 2038
rect 264336 1974 264388 1980
rect 264992 1630 265020 7278
rect 265360 2650 265388 9046
rect 267108 7546 267136 10882
rect 272156 10872 272208 10878
rect 272156 10814 272208 10820
rect 267648 8016 267700 8022
rect 267648 7958 267700 7964
rect 270958 7984 271014 7993
rect 267096 7540 267148 7546
rect 267096 7482 267148 7488
rect 267108 7410 267136 7482
rect 267096 7404 267148 7410
rect 267096 7346 267148 7352
rect 267660 6798 267688 7958
rect 270958 7919 271014 7928
rect 268384 7880 268436 7886
rect 268384 7822 268436 7828
rect 268396 6866 268424 7822
rect 270972 7410 271000 7919
rect 272168 7546 272196 10814
rect 275652 9036 275704 9042
rect 275652 8978 275704 8984
rect 272156 7540 272208 7546
rect 272156 7482 272208 7488
rect 272168 7410 272196 7482
rect 270960 7404 271012 7410
rect 270960 7346 271012 7352
rect 272156 7404 272208 7410
rect 272156 7346 272208 7352
rect 268384 6860 268436 6866
rect 268384 6802 268436 6808
rect 267648 6792 267700 6798
rect 267648 6734 267700 6740
rect 265992 6316 266044 6322
rect 265992 6258 266044 6264
rect 266004 5574 266032 6258
rect 268384 5704 268436 5710
rect 268384 5646 268436 5652
rect 269672 5704 269724 5710
rect 269672 5646 269724 5652
rect 265992 5568 266044 5574
rect 265992 5510 266044 5516
rect 266004 3738 266032 5510
rect 268396 5030 268424 5646
rect 269684 5030 269712 5646
rect 270592 5228 270644 5234
rect 270592 5170 270644 5176
rect 270604 5030 270632 5170
rect 271696 5160 271748 5166
rect 271696 5102 271748 5108
rect 268384 5024 268436 5030
rect 268384 4966 268436 4972
rect 269672 5024 269724 5030
rect 269672 4966 269724 4972
rect 270592 5024 270644 5030
rect 270592 4966 270644 4972
rect 265992 3732 266044 3738
rect 265992 3674 266044 3680
rect 265348 2644 265400 2650
rect 265348 2586 265400 2592
rect 265360 2446 265388 2586
rect 265348 2440 265400 2446
rect 265348 2382 265400 2388
rect 267188 2304 267240 2310
rect 267188 2246 267240 2252
rect 267924 2304 267976 2310
rect 267924 2246 267976 2252
rect 268016 2304 268068 2310
rect 268016 2246 268068 2252
rect 264980 1624 265032 1630
rect 264980 1566 265032 1572
rect 267200 1154 267228 2246
rect 267832 1420 267884 1426
rect 267832 1362 267884 1368
rect 267844 1290 267872 1362
rect 267936 1290 267964 2246
rect 267832 1284 267884 1290
rect 267832 1226 267884 1232
rect 267924 1284 267976 1290
rect 267924 1226 267976 1232
rect 268028 1222 268056 2246
rect 268396 1970 268424 4966
rect 268384 1964 268436 1970
rect 268384 1906 268436 1912
rect 269684 1902 269712 4966
rect 270500 3732 270552 3738
rect 270500 3674 270552 3680
rect 270512 2650 270540 3674
rect 270500 2644 270552 2650
rect 270500 2586 270552 2592
rect 270512 2446 270540 2586
rect 270500 2440 270552 2446
rect 270500 2382 270552 2388
rect 269856 2304 269908 2310
rect 269856 2246 269908 2252
rect 269672 1896 269724 1902
rect 269672 1838 269724 1844
rect 269868 1426 269896 2246
rect 270604 1834 270632 4966
rect 271708 4690 271736 5102
rect 271696 4684 271748 4690
rect 271696 4626 271748 4632
rect 273076 3528 273128 3534
rect 273076 3470 273128 3476
rect 273088 2650 273116 3470
rect 275664 2650 275692 8978
rect 276020 8356 276072 8362
rect 276020 8298 276072 8304
rect 276032 7954 276060 8298
rect 277136 8090 277164 11630
rect 311256 11416 311308 11422
rect 311256 11358 311308 11364
rect 282276 10736 282328 10742
rect 282276 10678 282328 10684
rect 282288 8090 282316 10678
rect 287428 10668 287480 10674
rect 287428 10610 287480 10616
rect 287440 8090 287468 10610
rect 292580 10600 292632 10606
rect 292580 10542 292632 10548
rect 292592 8090 292620 10542
rect 297732 10532 297784 10538
rect 297732 10474 297784 10480
rect 277124 8084 277176 8090
rect 277124 8026 277176 8032
rect 282276 8084 282328 8090
rect 282276 8026 282328 8032
rect 287152 8084 287204 8090
rect 287152 8026 287204 8032
rect 287428 8084 287480 8090
rect 287428 8026 287480 8032
rect 292580 8084 292632 8090
rect 292580 8026 292632 8032
rect 293868 8084 293920 8090
rect 293868 8026 293920 8032
rect 276020 7948 276072 7954
rect 276020 7890 276072 7896
rect 277136 7886 277164 8026
rect 282288 7886 282316 8026
rect 287164 7886 287192 8026
rect 292592 7886 292620 8026
rect 277124 7880 277176 7886
rect 277124 7822 277176 7828
rect 282276 7880 282328 7886
rect 282276 7822 282328 7828
rect 287152 7880 287204 7886
rect 287152 7822 287204 7828
rect 292580 7880 292632 7886
rect 292580 7822 292632 7828
rect 280344 7812 280396 7818
rect 280344 7754 280396 7760
rect 286140 7812 286192 7818
rect 286140 7754 286192 7760
rect 291200 7812 291252 7818
rect 291200 7754 291252 7760
rect 273076 2644 273128 2650
rect 273076 2586 273128 2592
rect 275652 2644 275704 2650
rect 275652 2586 275704 2592
rect 273088 2446 273116 2586
rect 275664 2446 275692 2586
rect 273076 2440 273128 2446
rect 273076 2382 273128 2388
rect 275652 2440 275704 2446
rect 275652 2382 275704 2388
rect 276020 2304 276072 2310
rect 276020 2246 276072 2252
rect 278228 2304 278280 2310
rect 278228 2246 278280 2252
rect 278780 2304 278832 2310
rect 278780 2246 278832 2252
rect 270592 1828 270644 1834
rect 270592 1770 270644 1776
rect 273996 1556 274048 1562
rect 273996 1498 274048 1504
rect 271604 1488 271656 1494
rect 271604 1430 271656 1436
rect 273352 1488 273404 1494
rect 273352 1430 273404 1436
rect 269856 1420 269908 1426
rect 269856 1362 269908 1368
rect 268016 1216 268068 1222
rect 268016 1158 268068 1164
rect 268660 1216 268712 1222
rect 268660 1158 268712 1164
rect 267188 1148 267240 1154
rect 267188 1090 267240 1096
rect 267740 1148 267792 1154
rect 267740 1090 267792 1096
rect 265440 944 265492 950
rect 265440 886 265492 892
rect 265452 678 265480 886
rect 265624 876 265676 882
rect 265900 876 265952 882
rect 265676 836 265900 864
rect 265624 818 265676 824
rect 265900 818 265952 824
rect 267752 746 267780 1090
rect 267832 944 267884 950
rect 267884 892 268240 898
rect 267832 886 268240 892
rect 267844 882 268240 886
rect 267844 876 268252 882
rect 267844 870 268200 876
rect 268200 818 268252 824
rect 268672 746 268700 1158
rect 271616 1086 271644 1430
rect 273364 1222 273392 1430
rect 273260 1216 273312 1222
rect 273166 1184 273222 1193
rect 273260 1158 273312 1164
rect 273352 1216 273404 1222
rect 273352 1158 273404 1164
rect 273166 1119 273222 1128
rect 271604 1080 271656 1086
rect 271604 1022 271656 1028
rect 271696 1080 271748 1086
rect 271696 1022 271748 1028
rect 271708 814 271736 1022
rect 273180 950 273208 1119
rect 273272 1068 273300 1158
rect 273272 1040 273392 1068
rect 273364 950 273392 1040
rect 273168 944 273220 950
rect 273168 886 273220 892
rect 273352 944 273404 950
rect 273352 886 273404 892
rect 271696 808 271748 814
rect 271696 750 271748 756
rect 274008 746 274036 1498
rect 274272 1420 274324 1426
rect 274272 1362 274324 1368
rect 274088 1012 274140 1018
rect 274088 954 274140 960
rect 267740 740 267792 746
rect 267740 682 267792 688
rect 268660 740 268712 746
rect 268660 682 268712 688
rect 273996 740 274048 746
rect 273996 682 274048 688
rect 265440 672 265492 678
rect 265440 614 265492 620
rect 274100 626 274128 954
rect 274284 882 274312 1362
rect 276032 1222 276060 2246
rect 278240 1630 278268 2246
rect 278228 1624 278280 1630
rect 278228 1566 278280 1572
rect 276020 1216 276072 1222
rect 276020 1158 276072 1164
rect 278044 1216 278096 1222
rect 278044 1158 278096 1164
rect 276480 1012 276532 1018
rect 276480 954 276532 960
rect 274272 876 274324 882
rect 274824 876 274876 882
rect 274272 818 274324 824
rect 274376 836 274824 864
rect 274376 762 274404 836
rect 274824 818 274876 824
rect 276492 814 276520 954
rect 278056 950 278084 1158
rect 278792 1034 278820 2246
rect 278962 1184 279018 1193
rect 278962 1119 279018 1128
rect 278608 1006 278820 1034
rect 278608 950 278636 1006
rect 278044 944 278096 950
rect 278044 886 278096 892
rect 278596 944 278648 950
rect 278596 886 278648 892
rect 278688 944 278740 950
rect 278688 886 278740 892
rect 274284 734 274404 762
rect 276480 808 276532 814
rect 276480 750 276532 756
rect 278596 808 278648 814
rect 278700 796 278728 886
rect 278976 882 279004 1119
rect 280356 882 280384 7754
rect 285956 5228 286008 5234
rect 285956 5170 286008 5176
rect 283380 5092 283432 5098
rect 283380 5034 283432 5040
rect 280804 4820 280856 4826
rect 280804 4762 280856 4768
rect 280816 2650 280844 4762
rect 283392 2650 283420 5034
rect 285968 2650 285996 5170
rect 286152 3505 286180 7754
rect 291212 7313 291240 7754
rect 291198 7304 291254 7313
rect 291198 7239 291254 7248
rect 291108 5296 291160 5302
rect 291108 5238 291160 5244
rect 288532 5160 288584 5166
rect 288532 5102 288584 5108
rect 286138 3496 286194 3505
rect 286138 3431 286194 3440
rect 288544 2650 288572 5102
rect 291120 2650 291148 5238
rect 293684 4752 293736 4758
rect 293684 4694 293736 4700
rect 293696 2650 293724 4694
rect 293880 4690 293908 8026
rect 297744 7886 297772 10474
rect 302424 10464 302476 10470
rect 302424 10406 302476 10412
rect 302436 8634 302464 10406
rect 307484 10396 307536 10402
rect 307484 10338 307536 10344
rect 306380 9716 306432 9722
rect 306380 9658 306432 9664
rect 302424 8628 302476 8634
rect 302424 8570 302476 8576
rect 302436 8498 302464 8570
rect 306392 8498 306420 9658
rect 307496 8634 307524 10338
rect 307484 8628 307536 8634
rect 307484 8570 307536 8576
rect 307496 8498 307524 8570
rect 311268 8498 311296 11358
rect 330764 11300 331084 11972
rect 330764 11244 330776 11300
rect 330832 11244 330856 11300
rect 330912 11244 330936 11300
rect 330992 11244 331016 11300
rect 331072 11244 331084 11300
rect 330764 11220 331084 11244
rect 330764 11164 330776 11220
rect 330832 11164 330856 11220
rect 330912 11164 330936 11220
rect 330992 11164 331016 11220
rect 331072 11164 331084 11220
rect 330764 11140 331084 11164
rect 330764 11084 330776 11140
rect 330832 11084 330856 11140
rect 330912 11084 330936 11140
rect 330992 11084 331016 11140
rect 331072 11084 331084 11140
rect 330764 11060 331084 11084
rect 330764 11004 330776 11060
rect 330832 11004 330856 11060
rect 330912 11004 330936 11060
rect 330992 11004 331016 11060
rect 331072 11004 331084 11060
rect 312452 10328 312504 10334
rect 312452 10270 312504 10276
rect 312464 8634 312492 10270
rect 316316 10260 316368 10266
rect 316316 10202 316368 10208
rect 317512 10260 317564 10266
rect 317512 10202 317564 10208
rect 312452 8628 312504 8634
rect 312452 8570 312504 8576
rect 312912 8628 312964 8634
rect 312912 8570 312964 8576
rect 312464 8498 312492 8570
rect 302424 8492 302476 8498
rect 302424 8434 302476 8440
rect 306380 8492 306432 8498
rect 306380 8434 306432 8440
rect 307484 8492 307536 8498
rect 307484 8434 307536 8440
rect 311256 8492 311308 8498
rect 311256 8434 311308 8440
rect 312452 8492 312504 8498
rect 312452 8434 312504 8440
rect 301228 8424 301280 8430
rect 301228 8366 301280 8372
rect 297732 7880 297784 7886
rect 297732 7822 297784 7828
rect 296168 7812 296220 7818
rect 296168 7754 296220 7760
rect 293868 4684 293920 4690
rect 293868 4626 293920 4632
rect 296180 3602 296208 7754
rect 298836 4072 298888 4078
rect 298836 4014 298888 4020
rect 296168 3596 296220 3602
rect 296168 3538 296220 3544
rect 296260 3392 296312 3398
rect 296260 3334 296312 3340
rect 296272 2650 296300 3334
rect 298848 2650 298876 4014
rect 301240 3670 301268 8366
rect 309140 4684 309192 4690
rect 309140 4626 309192 4632
rect 301412 4140 301464 4146
rect 301412 4082 301464 4088
rect 301228 3664 301280 3670
rect 301228 3606 301280 3612
rect 301424 2650 301452 4082
rect 306564 3664 306616 3670
rect 306564 3606 306616 3612
rect 303988 3596 304040 3602
rect 303988 3538 304040 3544
rect 304000 2650 304028 3538
rect 306576 2650 306604 3606
rect 309152 2650 309180 4626
rect 312924 4554 312952 8570
rect 316328 8498 316356 10202
rect 317524 8498 317552 10202
rect 322480 10192 322532 10198
rect 322480 10134 322532 10140
rect 321284 10056 321336 10062
rect 321284 9998 321336 10004
rect 321296 8974 321324 9998
rect 322492 8974 322520 10134
rect 326344 9988 326396 9994
rect 326344 9930 326396 9936
rect 326356 8974 326384 9930
rect 330764 9274 331084 11004
rect 330764 9222 330770 9274
rect 330822 9222 330834 9274
rect 330886 9222 330898 9274
rect 330950 9222 330962 9274
rect 331014 9222 331026 9274
rect 331078 9222 331084 9274
rect 330764 8988 331084 9222
rect 321284 8968 321336 8974
rect 321284 8910 321336 8916
rect 322480 8968 322532 8974
rect 322480 8910 322532 8916
rect 326344 8968 326396 8974
rect 326344 8910 326396 8916
rect 327540 8968 327592 8974
rect 327540 8910 327592 8916
rect 330764 8932 330776 8988
rect 330832 8932 330856 8988
rect 330912 8932 330936 8988
rect 330992 8932 331016 8988
rect 331072 8932 331084 8988
rect 327552 8838 327580 8910
rect 330764 8908 331084 8932
rect 330764 8852 330776 8908
rect 330832 8852 330856 8908
rect 330912 8852 330936 8908
rect 330992 8852 331016 8908
rect 331072 8852 331084 8908
rect 327540 8832 327592 8838
rect 327540 8774 327592 8780
rect 330764 8828 331084 8852
rect 316316 8492 316368 8498
rect 316316 8434 316368 8440
rect 317512 8492 317564 8498
rect 317512 8434 317564 8440
rect 327552 6866 327580 8774
rect 330764 8772 330776 8828
rect 330832 8772 330856 8828
rect 330912 8772 330936 8828
rect 330992 8772 331016 8828
rect 331072 8772 331084 8828
rect 330764 8748 331084 8772
rect 330764 8692 330776 8748
rect 330832 8692 330856 8748
rect 330912 8692 330936 8748
rect 330992 8692 331016 8748
rect 331072 8692 331084 8748
rect 330764 8186 331084 8692
rect 330764 8134 330770 8186
rect 330822 8134 330834 8186
rect 330886 8134 330898 8186
rect 330950 8134 330962 8186
rect 331014 8134 331026 8186
rect 331078 8134 331084 8186
rect 330764 7098 331084 8134
rect 330764 7046 330770 7098
rect 330822 7084 330834 7098
rect 330886 7084 330898 7098
rect 330950 7084 330962 7098
rect 331014 7084 331026 7098
rect 330832 7046 330834 7084
rect 331014 7046 331016 7084
rect 331078 7046 331084 7098
rect 330764 7028 330776 7046
rect 330832 7028 330856 7046
rect 330912 7028 330936 7046
rect 330992 7028 331016 7046
rect 331072 7028 331084 7046
rect 330764 7004 331084 7028
rect 330764 6948 330776 7004
rect 330832 6948 330856 7004
rect 330912 6948 330936 7004
rect 330992 6948 331016 7004
rect 331072 6948 331084 7004
rect 330764 6924 331084 6948
rect 330764 6868 330776 6924
rect 330832 6868 330856 6924
rect 330912 6868 330936 6924
rect 330992 6868 331016 6924
rect 331072 6868 331084 6924
rect 327540 6860 327592 6866
rect 327540 6802 327592 6808
rect 330764 6844 331084 6868
rect 330764 6788 330776 6844
rect 330832 6788 330856 6844
rect 330912 6788 330936 6844
rect 330992 6788 331016 6844
rect 331072 6788 331084 6844
rect 330764 6010 331084 6788
rect 330764 5958 330770 6010
rect 330822 5958 330834 6010
rect 330886 5958 330898 6010
rect 330950 5958 330962 6010
rect 331014 5958 331026 6010
rect 331078 5958 331084 6010
rect 330764 5180 331084 5958
rect 330764 5124 330776 5180
rect 330832 5124 330856 5180
rect 330912 5124 330936 5180
rect 330992 5124 331016 5180
rect 331072 5124 331084 5180
rect 330764 5100 331084 5124
rect 330764 5044 330776 5100
rect 330832 5044 330856 5100
rect 330912 5044 330936 5100
rect 330992 5044 331016 5100
rect 331072 5044 331084 5100
rect 330764 5020 331084 5044
rect 330764 4964 330776 5020
rect 330832 4964 330856 5020
rect 330912 4964 330936 5020
rect 330992 4964 331016 5020
rect 331072 4964 331084 5020
rect 330764 4940 331084 4964
rect 330764 4922 330776 4940
rect 330832 4922 330856 4940
rect 330912 4922 330936 4940
rect 330992 4922 331016 4940
rect 331072 4922 331084 4940
rect 330764 4870 330770 4922
rect 330832 4884 330834 4922
rect 331014 4884 331016 4922
rect 330822 4870 330834 4884
rect 330886 4870 330898 4884
rect 330950 4870 330962 4884
rect 331014 4870 331026 4884
rect 331078 4870 331084 4922
rect 322020 4616 322072 4622
rect 322020 4558 322072 4564
rect 312912 4548 312964 4554
rect 312912 4490 312964 4496
rect 319260 4004 319312 4010
rect 319260 3946 319312 3952
rect 319272 2650 319300 3946
rect 322032 2650 322060 4558
rect 330764 3834 331084 4870
rect 330764 3782 330770 3834
rect 330822 3782 330834 3834
rect 330886 3782 330898 3834
rect 330950 3782 330962 3834
rect 331014 3782 331026 3834
rect 331078 3782 331084 3834
rect 330764 3276 331084 3782
rect 330764 3220 330776 3276
rect 330832 3220 330856 3276
rect 330912 3220 330936 3276
rect 330992 3220 331016 3276
rect 331072 3220 331084 3276
rect 330764 3196 331084 3220
rect 330764 3140 330776 3196
rect 330832 3140 330856 3196
rect 330912 3140 330936 3196
rect 330992 3140 331016 3196
rect 331072 3140 331084 3196
rect 330764 3116 331084 3140
rect 330764 3060 330776 3116
rect 330832 3060 330856 3116
rect 330912 3060 330936 3116
rect 330992 3060 331016 3116
rect 331072 3060 331084 3116
rect 330764 3036 331084 3060
rect 330764 2980 330776 3036
rect 330832 2980 330856 3036
rect 330912 2980 330936 3036
rect 330992 2980 331016 3036
rect 331072 2980 331084 3036
rect 330764 2746 331084 2980
rect 330764 2694 330770 2746
rect 330822 2694 330834 2746
rect 330886 2694 330898 2746
rect 330950 2694 330962 2746
rect 331014 2694 331026 2746
rect 331078 2694 331084 2746
rect 280804 2644 280856 2650
rect 280804 2586 280856 2592
rect 283380 2644 283432 2650
rect 283380 2586 283432 2592
rect 285956 2644 286008 2650
rect 285956 2586 286008 2592
rect 288532 2644 288584 2650
rect 288532 2586 288584 2592
rect 291108 2644 291160 2650
rect 291108 2586 291160 2592
rect 293684 2644 293736 2650
rect 293684 2586 293736 2592
rect 296260 2644 296312 2650
rect 296260 2586 296312 2592
rect 298836 2644 298888 2650
rect 298836 2586 298888 2592
rect 301412 2644 301464 2650
rect 301412 2586 301464 2592
rect 303988 2644 304040 2650
rect 303988 2586 304040 2592
rect 306564 2644 306616 2650
rect 306564 2586 306616 2592
rect 309140 2644 309192 2650
rect 309140 2586 309192 2592
rect 319260 2644 319312 2650
rect 319260 2586 319312 2592
rect 322020 2644 322072 2650
rect 322020 2586 322072 2592
rect 280816 2446 280844 2586
rect 282460 2576 282512 2582
rect 282460 2518 282512 2524
rect 280804 2440 280856 2446
rect 280804 2382 280856 2388
rect 282368 1692 282420 1698
rect 282368 1634 282420 1640
rect 282276 1556 282328 1562
rect 282276 1498 282328 1504
rect 282288 1465 282316 1498
rect 282274 1456 282330 1465
rect 282274 1391 282330 1400
rect 282380 1018 282408 1634
rect 282472 1086 282500 2518
rect 283392 2446 283420 2586
rect 285968 2446 285996 2586
rect 288544 2446 288572 2586
rect 291120 2446 291148 2586
rect 291200 2576 291252 2582
rect 291200 2518 291252 2524
rect 283380 2440 283432 2446
rect 283380 2382 283432 2388
rect 285956 2440 286008 2446
rect 285956 2382 286008 2388
rect 288532 2440 288584 2446
rect 288532 2382 288584 2388
rect 291108 2440 291160 2446
rect 291108 2382 291160 2388
rect 282644 2304 282696 2310
rect 282644 2246 282696 2252
rect 282736 2304 282788 2310
rect 282736 2246 282788 2252
rect 285680 2304 285732 2310
rect 285680 2246 285732 2252
rect 289912 2304 289964 2310
rect 289912 2246 289964 2252
rect 282552 1556 282604 1562
rect 282552 1498 282604 1504
rect 282564 1222 282592 1498
rect 282656 1426 282684 2246
rect 282644 1420 282696 1426
rect 282644 1362 282696 1368
rect 282552 1216 282604 1222
rect 282552 1158 282604 1164
rect 282748 1154 282776 2246
rect 283104 1624 283156 1630
rect 282840 1550 283052 1578
rect 283104 1566 283156 1572
rect 282840 1290 282868 1550
rect 282920 1488 282972 1494
rect 282920 1430 282972 1436
rect 282828 1284 282880 1290
rect 282828 1226 282880 1232
rect 282736 1148 282788 1154
rect 282736 1090 282788 1096
rect 282460 1080 282512 1086
rect 282460 1022 282512 1028
rect 282368 1012 282420 1018
rect 282368 954 282420 960
rect 282828 1012 282880 1018
rect 282828 954 282880 960
rect 280896 944 280948 950
rect 280896 886 280948 892
rect 278964 876 279016 882
rect 278964 818 279016 824
rect 280344 876 280396 882
rect 280344 818 280396 824
rect 278648 768 278728 796
rect 278596 750 278648 756
rect 274284 626 274312 734
rect 274100 598 274312 626
rect 280908 610 280936 886
rect 282840 814 282868 954
rect 282932 882 282960 1430
rect 283024 1290 283052 1550
rect 283012 1284 283064 1290
rect 283012 1226 283064 1232
rect 283116 1086 283144 1566
rect 285692 1562 285720 2246
rect 285680 1556 285732 1562
rect 285680 1498 285732 1504
rect 283194 1456 283250 1465
rect 289924 1426 289952 2246
rect 291212 1698 291240 2518
rect 291752 2508 291804 2514
rect 291752 2450 291804 2456
rect 291200 1692 291252 1698
rect 291200 1634 291252 1640
rect 283194 1391 283196 1400
rect 283248 1391 283250 1400
rect 289912 1420 289964 1426
rect 283196 1362 283248 1368
rect 289912 1362 289964 1368
rect 291014 1184 291070 1193
rect 287244 1148 287296 1154
rect 291014 1119 291070 1128
rect 287244 1090 287296 1096
rect 283104 1080 283156 1086
rect 283104 1022 283156 1028
rect 283012 944 283064 950
rect 283196 944 283248 950
rect 283064 904 283196 932
rect 283012 886 283064 892
rect 283196 886 283248 892
rect 282920 876 282972 882
rect 282920 818 282972 824
rect 287256 814 287284 1090
rect 291028 1086 291056 1119
rect 287796 1080 287848 1086
rect 287796 1022 287848 1028
rect 291016 1080 291068 1086
rect 291016 1022 291068 1028
rect 291108 1080 291160 1086
rect 291108 1022 291160 1028
rect 287808 882 287836 1022
rect 289728 944 289780 950
rect 289556 892 289728 898
rect 289556 886 289780 892
rect 289556 882 289768 886
rect 287796 876 287848 882
rect 287796 818 287848 824
rect 289544 876 289768 882
rect 289596 870 289768 876
rect 289544 818 289596 824
rect 291120 814 291148 1022
rect 291764 882 291792 2450
rect 293696 2446 293724 2586
rect 296272 2446 296300 2586
rect 298192 2508 298244 2514
rect 298192 2450 298244 2456
rect 293684 2440 293736 2446
rect 293684 2382 293736 2388
rect 296260 2440 296312 2446
rect 296260 2382 296312 2388
rect 295248 2304 295300 2310
rect 295248 2246 295300 2252
rect 293500 1556 293552 1562
rect 293500 1498 293552 1504
rect 292210 1320 292266 1329
rect 292210 1255 292266 1264
rect 292224 1154 292252 1255
rect 292302 1184 292358 1193
rect 292212 1148 292264 1154
rect 293512 1154 293540 1498
rect 295260 1494 295288 2246
rect 295248 1488 295300 1494
rect 295248 1430 295300 1436
rect 298204 1426 298232 2450
rect 298848 2446 298876 2586
rect 301424 2446 301452 2586
rect 303528 2576 303580 2582
rect 303528 2518 303580 2524
rect 298836 2440 298888 2446
rect 298836 2382 298888 2388
rect 301412 2440 301464 2446
rect 301412 2382 301464 2388
rect 302700 2372 302752 2378
rect 302700 2314 302752 2320
rect 300860 2304 300912 2310
rect 300860 2246 300912 2252
rect 300872 1562 300900 2246
rect 302332 1964 302384 1970
rect 302332 1906 302384 1912
rect 300860 1556 300912 1562
rect 300860 1498 300912 1504
rect 295800 1420 295852 1426
rect 295800 1362 295852 1368
rect 298192 1420 298244 1426
rect 298192 1362 298244 1368
rect 300216 1420 300268 1426
rect 300216 1362 300268 1368
rect 292302 1119 292304 1128
rect 292212 1090 292264 1096
rect 292356 1119 292358 1128
rect 293500 1148 293552 1154
rect 292304 1090 292356 1096
rect 293500 1090 293552 1096
rect 293868 1012 293920 1018
rect 293868 954 293920 960
rect 291752 876 291804 882
rect 291752 818 291804 824
rect 293880 814 293908 954
rect 295812 950 295840 1362
rect 297546 1320 297602 1329
rect 297546 1255 297602 1264
rect 297560 1018 297588 1255
rect 300228 1018 300256 1362
rect 297548 1012 297600 1018
rect 297548 954 297600 960
rect 300216 1012 300268 1018
rect 300216 954 300268 960
rect 300400 1012 300452 1018
rect 300400 954 300452 960
rect 295800 944 295852 950
rect 295800 886 295852 892
rect 300412 814 300440 954
rect 302344 882 302372 1906
rect 302516 1488 302568 1494
rect 302516 1430 302568 1436
rect 302528 1154 302556 1430
rect 302516 1148 302568 1154
rect 302516 1090 302568 1096
rect 302712 1086 302740 2314
rect 303540 1426 303568 2518
rect 304000 2446 304028 2586
rect 306380 2508 306432 2514
rect 306380 2450 306432 2456
rect 303988 2440 304040 2446
rect 303988 2382 304040 2388
rect 306392 1494 306420 2450
rect 306576 2446 306604 2586
rect 309152 2446 309180 2586
rect 322032 2446 322060 2586
rect 306564 2440 306616 2446
rect 306564 2382 306616 2388
rect 309140 2440 309192 2446
rect 309140 2382 309192 2388
rect 314292 2440 314344 2446
rect 314292 2382 314344 2388
rect 319444 2440 319496 2446
rect 319444 2382 319496 2388
rect 322020 2440 322072 2446
rect 322020 2382 322072 2388
rect 329748 2440 329800 2446
rect 329748 2382 329800 2388
rect 309232 2372 309284 2378
rect 309232 2314 309284 2320
rect 306380 1488 306432 1494
rect 306380 1430 306432 1436
rect 303528 1420 303580 1426
rect 303528 1362 303580 1368
rect 306564 1420 306616 1426
rect 306564 1362 306616 1368
rect 304816 1148 304868 1154
rect 304816 1090 304868 1096
rect 302700 1080 302752 1086
rect 302700 1022 302752 1028
rect 302792 1012 302844 1018
rect 302792 954 302844 960
rect 302332 876 302384 882
rect 302332 818 302384 824
rect 282828 808 282880 814
rect 282828 750 282880 756
rect 287244 808 287296 814
rect 287244 750 287296 756
rect 291108 808 291160 814
rect 291108 750 291160 756
rect 293868 808 293920 814
rect 293868 750 293920 756
rect 300400 808 300452 814
rect 300400 750 300452 756
rect 302608 808 302660 814
rect 302804 796 302832 954
rect 304828 814 304856 1090
rect 306576 882 306604 1362
rect 306932 1080 306984 1086
rect 306932 1022 306984 1028
rect 306564 876 306616 882
rect 306564 818 306616 824
rect 306944 814 306972 1022
rect 308128 944 308180 950
rect 308128 886 308180 892
rect 307208 876 307260 882
rect 307392 876 307444 882
rect 307260 836 307392 864
rect 307208 818 307260 824
rect 307392 818 307444 824
rect 308140 814 308168 886
rect 302660 768 302832 796
rect 304816 808 304868 814
rect 302608 750 302660 756
rect 304816 750 304868 756
rect 306932 808 306984 814
rect 306932 750 306984 756
rect 308128 808 308180 814
rect 308128 750 308180 756
rect 280896 604 280948 610
rect 280896 546 280948 552
rect 293868 536 293920 542
rect 293866 504 293868 513
rect 293920 504 293922 513
rect 293866 439 293922 448
rect 298558 504 298614 513
rect 298558 439 298614 448
rect 300398 504 300454 513
rect 300398 439 300454 448
rect 309046 504 309102 513
rect 309046 439 309102 448
rect 250364 202 250668 206
rect 250352 196 250668 202
rect 250404 190 250668 196
rect 263428 190 263640 218
rect 250352 138 250404 144
rect 298572 134 298600 439
rect 300412 134 300440 439
rect 309060 354 309088 439
rect 309244 354 309272 2314
rect 314304 2310 314332 2382
rect 316684 2372 316736 2378
rect 316684 2314 316736 2320
rect 314292 2304 314344 2310
rect 314292 2246 314344 2252
rect 314304 1698 314332 2246
rect 314292 1692 314344 1698
rect 314292 1634 314344 1640
rect 316696 1494 316724 2314
rect 319456 2310 319484 2382
rect 329760 2310 329788 2382
rect 318708 2304 318760 2310
rect 318708 2246 318760 2252
rect 319444 2304 319496 2310
rect 319444 2246 319496 2252
rect 321284 2304 321336 2310
rect 321284 2246 321336 2252
rect 324596 2304 324648 2310
rect 324596 2246 324648 2252
rect 326436 2304 326488 2310
rect 326436 2246 326488 2252
rect 329012 2304 329064 2310
rect 329012 2246 329064 2252
rect 329748 2304 329800 2310
rect 329748 2246 329800 2252
rect 313372 1488 313424 1494
rect 313372 1430 313424 1436
rect 316684 1488 316736 1494
rect 316684 1430 316736 1436
rect 311898 1320 311954 1329
rect 311898 1255 311954 1264
rect 311070 1184 311126 1193
rect 311912 1154 311940 1255
rect 311990 1184 312046 1193
rect 311070 1119 311126 1128
rect 311900 1148 311952 1154
rect 311084 814 311112 1119
rect 311990 1119 311992 1128
rect 311900 1090 311952 1096
rect 312044 1119 312046 1128
rect 311992 1090 312044 1096
rect 313384 882 313412 1430
rect 318720 1426 318748 2246
rect 319456 1494 319484 2246
rect 321296 1970 321324 2246
rect 321284 1964 321336 1970
rect 321284 1906 321336 1912
rect 324608 1562 324636 2246
rect 324596 1556 324648 1562
rect 324596 1498 324648 1504
rect 319444 1488 319496 1494
rect 319444 1430 319496 1436
rect 318708 1420 318760 1426
rect 318708 1362 318760 1368
rect 318062 1320 318118 1329
rect 318062 1255 318118 1264
rect 316512 1142 316908 1170
rect 316512 1018 316540 1142
rect 316880 1018 316908 1142
rect 315304 1012 315356 1018
rect 315304 954 315356 960
rect 316500 1012 316552 1018
rect 316500 954 316552 960
rect 316868 1012 316920 1018
rect 316868 954 316920 960
rect 313372 876 313424 882
rect 313372 818 313424 824
rect 311072 808 311124 814
rect 311072 750 311124 756
rect 315316 513 315344 954
rect 316960 944 317012 950
rect 316960 886 317012 892
rect 316972 814 317000 886
rect 315672 808 315724 814
rect 315948 808 316000 814
rect 315724 768 315948 796
rect 315672 750 315724 756
rect 315948 750 316000 756
rect 316960 808 317012 814
rect 316960 750 317012 756
rect 315302 504 315358 513
rect 315302 439 315358 448
rect 309060 326 309272 354
rect 318076 270 318104 1255
rect 318246 504 318302 513
rect 318246 439 318302 448
rect 318064 264 318116 270
rect 318064 206 318116 212
rect 318260 202 318288 439
rect 326448 202 326476 2246
rect 329024 270 329052 2246
rect 329760 1970 329788 2246
rect 329748 1964 329800 1970
rect 329748 1906 329800 1912
rect 330764 964 331084 2694
rect 331424 11960 331744 11972
rect 331424 11904 331436 11960
rect 331492 11904 331516 11960
rect 331572 11904 331596 11960
rect 331652 11904 331676 11960
rect 331732 11904 331744 11960
rect 331424 11880 331744 11904
rect 331424 11824 331436 11880
rect 331492 11824 331516 11880
rect 331572 11824 331596 11880
rect 331652 11824 331676 11880
rect 331732 11824 331744 11880
rect 331424 11800 331744 11824
rect 331424 11744 331436 11800
rect 331492 11744 331516 11800
rect 331572 11744 331596 11800
rect 331652 11744 331676 11800
rect 331732 11744 331744 11800
rect 331424 11720 331744 11744
rect 331424 11664 331436 11720
rect 331492 11664 331516 11720
rect 331572 11664 331596 11720
rect 331652 11664 331676 11720
rect 331732 11664 331744 11720
rect 331424 9818 331744 11664
rect 359740 11688 359792 11694
rect 359740 11630 359792 11636
rect 354404 11552 354456 11558
rect 354404 11494 354456 11500
rect 346768 11348 346820 11354
rect 346768 11290 346820 11296
rect 347596 11348 347648 11354
rect 347596 11290 347648 11296
rect 336280 11212 336332 11218
rect 336280 11154 336332 11160
rect 342720 11212 342772 11218
rect 342720 11154 342772 11160
rect 332508 10124 332560 10130
rect 332508 10066 332560 10072
rect 331424 9766 331430 9818
rect 331482 9766 331494 9818
rect 331546 9766 331558 9818
rect 331610 9766 331622 9818
rect 331674 9766 331686 9818
rect 331738 9766 331744 9818
rect 331424 9648 331744 9766
rect 331424 9592 331436 9648
rect 331492 9592 331516 9648
rect 331572 9592 331596 9648
rect 331652 9592 331676 9648
rect 331732 9592 331744 9648
rect 331424 9568 331744 9592
rect 331424 9512 331436 9568
rect 331492 9512 331516 9568
rect 331572 9512 331596 9568
rect 331652 9512 331676 9568
rect 331732 9512 331744 9568
rect 331424 9488 331744 9512
rect 331424 9432 331436 9488
rect 331492 9432 331516 9488
rect 331572 9432 331596 9488
rect 331652 9432 331676 9488
rect 331732 9432 331744 9488
rect 331424 9408 331744 9432
rect 331424 9352 331436 9408
rect 331492 9352 331516 9408
rect 331572 9352 331596 9408
rect 331652 9352 331676 9408
rect 331732 9352 331744 9408
rect 331424 8730 331744 9352
rect 332520 8974 332548 10066
rect 336292 8974 336320 11154
rect 337476 10056 337528 10062
rect 337476 9998 337528 10004
rect 337488 8974 337516 9998
rect 340144 9988 340196 9994
rect 340144 9930 340196 9936
rect 340156 9654 340184 9930
rect 342732 9654 342760 11154
rect 340144 9648 340196 9654
rect 340144 9590 340196 9596
rect 342720 9648 342772 9654
rect 342720 9590 342772 9596
rect 346780 9586 346808 11290
rect 347608 9586 347636 11290
rect 354416 9654 354444 11494
rect 358636 11484 358688 11490
rect 358636 11426 358688 11432
rect 355784 11348 355836 11354
rect 355784 11290 355836 11296
rect 355416 11212 355468 11218
rect 355416 11154 355468 11160
rect 354496 11076 354548 11082
rect 354496 11018 354548 11024
rect 354508 10810 354536 11018
rect 355428 10946 355456 11154
rect 355796 11150 355824 11290
rect 355784 11144 355836 11150
rect 355784 11086 355836 11092
rect 355416 10940 355468 10946
rect 355416 10882 355468 10888
rect 354496 10804 354548 10810
rect 354496 10746 354548 10752
rect 354404 9648 354456 9654
rect 354404 9590 354456 9596
rect 354588 9648 354640 9654
rect 354588 9590 354640 9596
rect 346768 9580 346820 9586
rect 346768 9522 346820 9528
rect 347596 9580 347648 9586
rect 347596 9522 347648 9528
rect 350080 9580 350132 9586
rect 350080 9522 350132 9528
rect 338948 9512 339000 9518
rect 338948 9454 339000 9460
rect 344100 9512 344152 9518
rect 344100 9454 344152 9460
rect 349344 9512 349396 9518
rect 349344 9454 349396 9460
rect 338960 9178 338988 9454
rect 338948 9172 339000 9178
rect 338948 9114 339000 9120
rect 332508 8968 332560 8974
rect 332508 8910 332560 8916
rect 336280 8968 336332 8974
rect 336280 8910 336332 8916
rect 337476 8968 337528 8974
rect 337476 8910 337528 8916
rect 331424 8678 331430 8730
rect 331482 8678 331494 8730
rect 331546 8678 331558 8730
rect 331610 8678 331622 8730
rect 331674 8678 331686 8730
rect 331738 8678 331744 8730
rect 331424 7744 331744 8678
rect 331424 7688 331436 7744
rect 331492 7688 331516 7744
rect 331572 7688 331596 7744
rect 331652 7688 331676 7744
rect 331732 7688 331744 7744
rect 331424 7664 331744 7688
rect 331424 7642 331436 7664
rect 331492 7642 331516 7664
rect 331572 7642 331596 7664
rect 331652 7642 331676 7664
rect 331732 7642 331744 7664
rect 331424 7590 331430 7642
rect 331492 7608 331494 7642
rect 331674 7608 331676 7642
rect 331482 7590 331494 7608
rect 331546 7590 331558 7608
rect 331610 7590 331622 7608
rect 331674 7590 331686 7608
rect 331738 7590 331744 7642
rect 331424 7584 331744 7590
rect 331424 7528 331436 7584
rect 331492 7528 331516 7584
rect 331572 7528 331596 7584
rect 331652 7528 331676 7584
rect 331732 7528 331744 7584
rect 331424 7504 331744 7528
rect 331424 7448 331436 7504
rect 331492 7448 331516 7504
rect 331572 7448 331596 7504
rect 331652 7448 331676 7504
rect 331732 7448 331744 7504
rect 344112 7478 344140 9454
rect 349356 8566 349384 9454
rect 350092 9382 350120 9522
rect 351920 9512 351972 9518
rect 351920 9454 351972 9460
rect 350080 9376 350132 9382
rect 350080 9318 350132 9324
rect 350092 8566 350120 9318
rect 351932 8634 351960 9454
rect 354600 9450 354628 9590
rect 358648 9586 358676 11426
rect 359752 10849 359780 11630
rect 359924 11620 359976 11626
rect 359924 11562 359976 11568
rect 359936 11529 359964 11562
rect 446680 11552 446732 11558
rect 359922 11520 359978 11529
rect 359922 11455 359978 11464
rect 363142 11520 363198 11529
rect 363142 11455 363144 11464
rect 363196 11455 363198 11464
rect 446600 11500 446680 11506
rect 446600 11494 446732 11500
rect 446600 11478 446720 11494
rect 363144 11426 363196 11432
rect 445852 11416 445904 11422
rect 445772 11364 445852 11370
rect 445772 11358 445904 11364
rect 441804 11348 441856 11354
rect 441804 11290 441856 11296
rect 442908 11348 442960 11354
rect 442908 11290 442960 11296
rect 445772 11342 445892 11358
rect 360752 11280 360804 11286
rect 360752 11222 360804 11228
rect 360936 11280 360988 11286
rect 360936 11222 360988 11228
rect 361304 11280 361356 11286
rect 361304 11222 361356 11228
rect 362040 11280 362092 11286
rect 362040 11222 362092 11228
rect 362408 11280 362460 11286
rect 362408 11222 362460 11228
rect 363696 11280 363748 11286
rect 363696 11222 363748 11228
rect 364248 11280 364300 11286
rect 364248 11222 364300 11228
rect 365260 11280 365312 11286
rect 365260 11222 365312 11228
rect 365812 11280 365864 11286
rect 365812 11222 365864 11228
rect 366364 11280 366416 11286
rect 366364 11222 366416 11228
rect 366732 11280 366784 11286
rect 366732 11222 366784 11228
rect 367468 11280 367520 11286
rect 367468 11222 367520 11228
rect 368020 11280 368072 11286
rect 368020 11222 368072 11228
rect 368664 11280 368716 11286
rect 368664 11222 368716 11228
rect 369768 11280 369820 11286
rect 369768 11222 369820 11228
rect 370136 11280 370188 11286
rect 370136 11222 370188 11228
rect 370688 11280 370740 11286
rect 370688 11222 370740 11228
rect 371056 11280 371108 11286
rect 371056 11222 371108 11228
rect 371792 11280 371844 11286
rect 371792 11222 371844 11228
rect 372160 11280 372212 11286
rect 372160 11222 372212 11228
rect 372896 11280 372948 11286
rect 372896 11222 372948 11228
rect 373264 11280 373316 11286
rect 373264 11222 373316 11228
rect 374000 11280 374052 11286
rect 374000 11222 374052 11228
rect 374368 11280 374420 11286
rect 374368 11222 374420 11228
rect 375104 11280 375156 11286
rect 375104 11222 375156 11228
rect 375472 11280 375524 11286
rect 375472 11222 375524 11228
rect 376208 11280 376260 11286
rect 376208 11222 376260 11228
rect 377036 11280 377088 11286
rect 377036 11222 377088 11228
rect 377312 11280 377364 11286
rect 377312 11222 377364 11228
rect 377588 11280 377640 11286
rect 377588 11222 377640 11228
rect 378416 11280 378468 11286
rect 378416 11222 378468 11228
rect 378692 11280 378744 11286
rect 378692 11222 378744 11228
rect 379428 11280 379480 11286
rect 379428 11222 379480 11228
rect 380348 11280 380400 11286
rect 380348 11222 380400 11228
rect 381544 11280 381596 11286
rect 381544 11222 381596 11228
rect 382096 11280 382148 11286
rect 382096 11222 382148 11228
rect 382464 11280 382516 11286
rect 382464 11222 382516 11228
rect 383200 11280 383252 11286
rect 383200 11222 383252 11228
rect 384672 11280 384724 11286
rect 384672 11222 384724 11228
rect 385224 11280 385276 11286
rect 385224 11222 385276 11228
rect 385960 11280 386012 11286
rect 385960 11222 386012 11228
rect 386512 11280 386564 11286
rect 386512 11222 386564 11228
rect 387984 11280 388036 11286
rect 387984 11222 388036 11228
rect 389824 11280 389876 11286
rect 389824 11222 389876 11228
rect 390652 11280 390704 11286
rect 390652 11222 390704 11228
rect 391388 11280 391440 11286
rect 391388 11222 391440 11228
rect 391940 11280 391992 11286
rect 391940 11222 391992 11228
rect 392492 11280 392544 11286
rect 392492 11222 392544 11228
rect 392860 11280 392912 11286
rect 392860 11222 392912 11228
rect 393504 11280 393556 11286
rect 393504 11222 393556 11228
rect 394056 11280 394108 11286
rect 394056 11222 394108 11228
rect 394700 11280 394752 11286
rect 394700 11222 394752 11228
rect 395160 11280 395212 11286
rect 395160 11222 395212 11228
rect 395528 11280 395580 11286
rect 395528 11222 395580 11228
rect 396264 11280 396316 11286
rect 396264 11222 396316 11228
rect 397920 11280 397972 11286
rect 397920 11222 397972 11228
rect 398472 11280 398524 11286
rect 398472 11222 398524 11228
rect 400680 11280 400732 11286
rect 400680 11222 400732 11228
rect 400956 11280 401008 11286
rect 400956 11222 401008 11228
rect 402336 11280 402388 11286
rect 402336 11222 402388 11228
rect 403900 11280 403952 11286
rect 403900 11222 403952 11228
rect 438860 11280 438912 11286
rect 438860 11222 438912 11228
rect 440148 11280 440200 11286
rect 440148 11222 440200 11228
rect 440424 11280 440476 11286
rect 440424 11222 440476 11228
rect 440700 11280 440752 11286
rect 440700 11222 440752 11228
rect 360304 10934 360700 10962
rect 360304 10878 360332 10934
rect 360292 10872 360344 10878
rect 359738 10840 359794 10849
rect 359556 10804 359608 10810
rect 360292 10814 360344 10820
rect 360566 10840 360622 10849
rect 359738 10775 359794 10784
rect 360566 10775 360622 10784
rect 359556 10746 359608 10752
rect 359568 10577 359596 10746
rect 360108 10736 360160 10742
rect 360108 10678 360160 10684
rect 360198 10704 360254 10713
rect 359554 10568 359610 10577
rect 359554 10503 359610 10512
rect 360120 10441 360148 10678
rect 360580 10674 360608 10775
rect 360672 10742 360700 10934
rect 360660 10736 360712 10742
rect 360660 10678 360712 10684
rect 360198 10639 360254 10648
rect 360568 10668 360620 10674
rect 360212 10606 360240 10639
rect 360568 10610 360620 10616
rect 360200 10600 360252 10606
rect 360200 10542 360252 10548
rect 360106 10432 360162 10441
rect 360106 10367 360162 10376
rect 355324 9580 355376 9586
rect 355324 9522 355376 9528
rect 357900 9580 357952 9586
rect 357900 9522 357952 9528
rect 358636 9580 358688 9586
rect 358636 9522 358688 9528
rect 354588 9444 354640 9450
rect 354588 9386 354640 9392
rect 355336 9382 355364 9522
rect 357072 9512 357124 9518
rect 357072 9454 357124 9460
rect 355324 9376 355376 9382
rect 355324 9318 355376 9324
rect 355336 8974 355364 9318
rect 355324 8968 355376 8974
rect 355324 8910 355376 8916
rect 351920 8628 351972 8634
rect 351920 8570 351972 8576
rect 349344 8560 349396 8566
rect 349344 8502 349396 8508
rect 350080 8560 350132 8566
rect 350080 8502 350132 8508
rect 349068 7744 349120 7750
rect 349068 7686 349120 7692
rect 331424 6554 331744 7448
rect 344100 7472 344152 7478
rect 344100 7414 344152 7420
rect 331424 6502 331430 6554
rect 331482 6502 331494 6554
rect 331546 6502 331558 6554
rect 331610 6502 331622 6554
rect 331674 6502 331686 6554
rect 331738 6502 331744 6554
rect 331424 5840 331744 6502
rect 331424 5784 331436 5840
rect 331492 5784 331516 5840
rect 331572 5784 331596 5840
rect 331652 5784 331676 5840
rect 331732 5784 331744 5840
rect 331424 5760 331744 5784
rect 331424 5704 331436 5760
rect 331492 5704 331516 5760
rect 331572 5704 331596 5760
rect 331652 5704 331676 5760
rect 331732 5704 331744 5760
rect 331424 5680 331744 5704
rect 331424 5624 331436 5680
rect 331492 5624 331516 5680
rect 331572 5624 331596 5680
rect 331652 5624 331676 5680
rect 331732 5624 331744 5680
rect 331424 5600 331744 5624
rect 331424 5544 331436 5600
rect 331492 5544 331516 5600
rect 331572 5544 331596 5600
rect 331652 5544 331676 5600
rect 331732 5544 331744 5600
rect 331424 5466 331744 5544
rect 331424 5414 331430 5466
rect 331482 5414 331494 5466
rect 331546 5414 331558 5466
rect 331610 5414 331622 5466
rect 331674 5414 331686 5466
rect 331738 5414 331744 5466
rect 331424 4378 331744 5414
rect 334900 4548 334952 4554
rect 334900 4490 334952 4496
rect 331424 4326 331430 4378
rect 331482 4326 331494 4378
rect 331546 4326 331558 4378
rect 331610 4326 331622 4378
rect 331674 4326 331686 4378
rect 331738 4326 331744 4378
rect 331424 3936 331744 4326
rect 331424 3880 331436 3936
rect 331492 3880 331516 3936
rect 331572 3880 331596 3936
rect 331652 3880 331676 3936
rect 331732 3880 331744 3936
rect 331424 3856 331744 3880
rect 331424 3800 331436 3856
rect 331492 3800 331516 3856
rect 331572 3800 331596 3856
rect 331652 3800 331676 3856
rect 331732 3800 331744 3856
rect 331424 3776 331744 3800
rect 331424 3720 331436 3776
rect 331492 3720 331516 3776
rect 331572 3720 331596 3776
rect 331652 3720 331676 3776
rect 331732 3720 331744 3776
rect 331424 3696 331744 3720
rect 331424 3640 331436 3696
rect 331492 3640 331516 3696
rect 331572 3640 331596 3696
rect 331652 3640 331676 3696
rect 331732 3640 331744 3696
rect 331424 3290 331744 3640
rect 331424 3238 331430 3290
rect 331482 3238 331494 3290
rect 331546 3238 331558 3290
rect 331610 3238 331622 3290
rect 331674 3238 331686 3290
rect 331738 3238 331744 3290
rect 331220 2304 331272 2310
rect 331220 2246 331272 2252
rect 331232 1018 331260 2246
rect 331424 2202 331744 3238
rect 334912 2582 334940 4490
rect 349080 2582 349108 7686
rect 357084 4486 357112 9454
rect 357912 9382 357940 9522
rect 360200 9512 360252 9518
rect 360200 9454 360252 9460
rect 357900 9376 357952 9382
rect 357900 9318 357952 9324
rect 357440 9172 357492 9178
rect 357440 9114 357492 9120
rect 357072 4480 357124 4486
rect 357072 4422 357124 4428
rect 355508 3936 355560 3942
rect 355508 3878 355560 3884
rect 351920 3188 351972 3194
rect 351920 3130 351972 3136
rect 334900 2576 334952 2582
rect 334900 2518 334952 2524
rect 349068 2576 349120 2582
rect 349068 2518 349120 2524
rect 351932 2514 351960 3130
rect 355520 2582 355548 3878
rect 357452 3738 357480 9114
rect 357912 8634 357940 9318
rect 357900 8628 357952 8634
rect 357900 8570 357952 8576
rect 358820 7540 358872 7546
rect 358820 7482 358872 7488
rect 358832 6730 358860 7482
rect 358820 6724 358872 6730
rect 358820 6666 358872 6672
rect 357440 3732 357492 3738
rect 357440 3674 357492 3680
rect 355416 2576 355468 2582
rect 352930 2544 352986 2553
rect 351920 2508 351972 2514
rect 355416 2518 355468 2524
rect 355508 2576 355560 2582
rect 355508 2518 355560 2524
rect 352930 2479 352932 2488
rect 351920 2450 351972 2456
rect 352984 2479 352986 2488
rect 352932 2450 352984 2456
rect 332324 2440 332376 2446
rect 332324 2382 332376 2388
rect 337476 2440 337528 2446
rect 337476 2382 337528 2388
rect 340052 2440 340104 2446
rect 340052 2382 340104 2388
rect 342628 2440 342680 2446
rect 342628 2382 342680 2388
rect 345204 2440 345256 2446
rect 345204 2382 345256 2388
rect 350354 2408 350410 2417
rect 332336 2310 332364 2382
rect 337488 2310 337516 2382
rect 340064 2310 340092 2382
rect 342640 2310 342668 2382
rect 345216 2310 345244 2382
rect 350354 2343 350356 2352
rect 350408 2343 350410 2352
rect 350356 2314 350408 2320
rect 332324 2304 332376 2310
rect 332324 2246 332376 2252
rect 334164 2304 334216 2310
rect 334164 2246 334216 2252
rect 336740 2304 336792 2310
rect 336740 2246 336792 2252
rect 337476 2304 337528 2310
rect 337476 2246 337528 2252
rect 339316 2304 339368 2310
rect 339316 2246 339368 2252
rect 340052 2304 340104 2310
rect 340052 2246 340104 2252
rect 341892 2304 341944 2310
rect 341892 2246 341944 2252
rect 342628 2304 342680 2310
rect 342628 2246 342680 2252
rect 344468 2304 344520 2310
rect 344468 2246 344520 2252
rect 345204 2304 345256 2310
rect 345204 2246 345256 2252
rect 347044 2304 347096 2310
rect 347044 2246 347096 2252
rect 352196 2304 352248 2310
rect 352196 2246 352248 2252
rect 331424 2150 331430 2202
rect 331482 2150 331494 2202
rect 331546 2150 331558 2202
rect 331610 2150 331622 2202
rect 331674 2150 331686 2202
rect 331738 2150 331744 2202
rect 330764 908 330776 964
rect 330832 908 330856 964
rect 330912 908 330936 964
rect 330992 908 331016 964
rect 331072 908 331084 964
rect 331220 1012 331272 1018
rect 331220 954 331272 960
rect 330764 884 331084 908
rect 330764 828 330776 884
rect 330832 828 330856 884
rect 330912 828 330936 884
rect 330992 828 331016 884
rect 331072 828 331084 884
rect 330764 804 331084 828
rect 330764 748 330776 804
rect 330832 748 330856 804
rect 330912 748 330936 804
rect 330992 748 331016 804
rect 331072 748 331084 804
rect 330764 724 331084 748
rect 330764 668 330776 724
rect 330832 668 330856 724
rect 330912 668 330936 724
rect 330992 668 331016 724
rect 331072 668 331084 724
rect 329012 264 329064 270
rect 329012 206 329064 212
rect 318248 196 318300 202
rect 318248 138 318300 144
rect 326436 196 326488 202
rect 326436 138 326488 144
rect 298560 128 298612 134
rect 298560 70 298612 76
rect 300400 128 300452 134
rect 300400 70 300452 76
rect 199496 8 199508 64
rect 199564 8 199588 64
rect 199644 8 199668 64
rect 199724 8 199748 64
rect 199804 8 199816 64
rect 199496 -4 199816 8
rect 219716 60 219768 66
rect 219716 2 219768 8
rect 317880 60 317932 66
rect 318064 60 318116 66
rect 317932 20 318064 48
rect 317880 2 317932 8
rect 318064 2 318116 8
rect 330764 -4 331084 668
rect 331424 304 331744 2150
rect 332336 1426 332364 2246
rect 332324 1420 332376 1426
rect 332324 1362 332376 1368
rect 334176 1086 334204 2246
rect 336752 1154 336780 2246
rect 337488 1766 337516 2246
rect 337476 1760 337528 1766
rect 337476 1702 337528 1708
rect 336740 1148 336792 1154
rect 336740 1090 336792 1096
rect 334164 1080 334216 1086
rect 334164 1022 334216 1028
rect 339328 882 339356 2246
rect 340064 2106 340092 2246
rect 340052 2100 340104 2106
rect 340052 2042 340104 2048
rect 341904 950 341932 2246
rect 342640 2038 342668 2246
rect 342628 2032 342680 2038
rect 342628 1974 342680 1980
rect 341892 944 341944 950
rect 341892 886 341944 892
rect 339316 876 339368 882
rect 339316 818 339368 824
rect 331424 248 331436 304
rect 331492 248 331516 304
rect 331572 248 331596 304
rect 331652 248 331676 304
rect 331732 248 331744 304
rect 331424 224 331744 248
rect 331424 168 331436 224
rect 331492 168 331516 224
rect 331572 168 331596 224
rect 331652 168 331676 224
rect 331732 168 331744 224
rect 331424 144 331744 168
rect 331424 88 331436 144
rect 331492 88 331516 144
rect 331572 88 331596 144
rect 331652 88 331676 144
rect 331732 88 331744 144
rect 331424 64 331744 88
rect 344480 66 344508 2246
rect 345216 1630 345244 2246
rect 345204 1624 345256 1630
rect 345204 1566 345256 1572
rect 347056 134 347084 2246
rect 352208 1834 352236 2246
rect 352196 1828 352248 1834
rect 352196 1770 352248 1776
rect 355428 814 355456 2518
rect 357992 2372 358044 2378
rect 357992 2314 358044 2320
rect 357348 2304 357400 2310
rect 357348 2246 357400 2252
rect 357360 950 357388 2246
rect 358004 1086 358032 2314
rect 358084 2304 358136 2310
rect 358084 2246 358136 2252
rect 359924 2304 359976 2310
rect 359924 2246 359976 2252
rect 358096 1902 358124 2246
rect 358084 1896 358136 1902
rect 358084 1838 358136 1844
rect 359832 1828 359884 1834
rect 359832 1770 359884 1776
rect 357992 1080 358044 1086
rect 357992 1022 358044 1028
rect 357348 944 357400 950
rect 357348 886 357400 892
rect 359844 882 359872 1770
rect 359936 1018 359964 2246
rect 360212 1358 360240 9454
rect 360764 5370 360792 11222
rect 360948 6934 360976 11222
rect 361316 10577 361344 11222
rect 361396 11008 361448 11014
rect 361396 10950 361448 10956
rect 361408 10810 361436 10950
rect 361396 10804 361448 10810
rect 361396 10746 361448 10752
rect 361302 10568 361358 10577
rect 361302 10503 361358 10512
rect 361488 8288 361540 8294
rect 361488 8230 361540 8236
rect 360936 6928 360988 6934
rect 360936 6870 360988 6876
rect 360752 5364 360804 5370
rect 360752 5306 360804 5312
rect 360660 5024 360712 5030
rect 360660 4966 360712 4972
rect 360672 2650 360700 4966
rect 361500 4554 361528 8230
rect 362052 7274 362080 11222
rect 362420 11082 362448 11222
rect 362592 11144 362644 11150
rect 362592 11086 362644 11092
rect 362408 11076 362460 11082
rect 362408 11018 362460 11024
rect 362604 10946 362632 11086
rect 363420 11008 363472 11014
rect 363420 10950 363472 10956
rect 362592 10940 362644 10946
rect 362592 10882 362644 10888
rect 363328 10872 363380 10878
rect 363328 10814 363380 10820
rect 363340 10713 363368 10814
rect 363326 10704 363382 10713
rect 363326 10639 363382 10648
rect 363432 10606 363460 10950
rect 363708 10810 363736 11222
rect 363696 10804 363748 10810
rect 363696 10746 363748 10752
rect 364156 10804 364208 10810
rect 364156 10746 364208 10752
rect 363420 10600 363472 10606
rect 363420 10542 363472 10548
rect 362132 9512 362184 9518
rect 362132 9454 362184 9460
rect 363696 9512 363748 9518
rect 363696 9454 363748 9460
rect 362144 8906 362172 9454
rect 362132 8900 362184 8906
rect 362132 8842 362184 8848
rect 362316 7472 362368 7478
rect 362316 7414 362368 7420
rect 362040 7268 362092 7274
rect 362040 7210 362092 7216
rect 361580 6724 361632 6730
rect 361580 6666 361632 6672
rect 361488 4548 361540 4554
rect 361488 4490 361540 4496
rect 360660 2644 360712 2650
rect 360660 2586 360712 2592
rect 360672 2446 360700 2586
rect 360660 2440 360712 2446
rect 360660 2382 360712 2388
rect 361592 1698 361620 6666
rect 362328 6458 362356 7414
rect 362316 6452 362368 6458
rect 362316 6394 362368 6400
rect 363708 3466 363736 9454
rect 364168 8974 364196 10746
rect 364156 8968 364208 8974
rect 364156 8910 364208 8916
rect 364260 8022 364288 11222
rect 364524 11212 364576 11218
rect 364524 11154 364576 11160
rect 364536 10742 364564 11154
rect 364984 10940 365036 10946
rect 364984 10882 365036 10888
rect 364524 10736 364576 10742
rect 364524 10678 364576 10684
rect 364996 8566 365024 10882
rect 364984 8560 365036 8566
rect 364984 8502 365036 8508
rect 364248 8016 364300 8022
rect 364248 7958 364300 7964
rect 364708 7948 364760 7954
rect 364708 7890 364760 7896
rect 363696 3460 363748 3466
rect 363696 3402 363748 3408
rect 364720 3398 364748 7890
rect 364984 7404 365036 7410
rect 364984 7346 365036 7352
rect 364996 6254 365024 7346
rect 365272 7002 365300 11222
rect 365824 10674 365852 11222
rect 365812 10668 365864 10674
rect 365812 10610 365864 10616
rect 365812 8968 365864 8974
rect 365812 8910 365864 8916
rect 365720 8016 365772 8022
rect 365720 7958 365772 7964
rect 365260 6996 365312 7002
rect 365260 6938 365312 6944
rect 365628 6656 365680 6662
rect 365628 6598 365680 6604
rect 364984 6248 365036 6254
rect 364984 6190 365036 6196
rect 364708 3392 364760 3398
rect 364708 3334 364760 3340
rect 365076 2644 365128 2650
rect 365076 2586 365128 2592
rect 365260 2644 365312 2650
rect 365260 2586 365312 2592
rect 361580 1692 361632 1698
rect 361580 1634 361632 1640
rect 360200 1352 360252 1358
rect 360200 1294 360252 1300
rect 365088 1154 365116 2586
rect 365272 2446 365300 2586
rect 365260 2440 365312 2446
rect 365260 2382 365312 2388
rect 365640 1970 365668 6598
rect 365732 5846 365760 7958
rect 365720 5840 365772 5846
rect 365720 5782 365772 5788
rect 365824 3534 365852 8910
rect 366272 8424 366324 8430
rect 366272 8366 366324 8372
rect 366284 7886 366312 8366
rect 366272 7880 366324 7886
rect 366272 7822 366324 7828
rect 366376 7818 366404 11222
rect 366744 10441 366772 11222
rect 367100 10600 367152 10606
rect 367100 10542 367152 10548
rect 366730 10432 366786 10441
rect 366730 10367 366786 10376
rect 367112 9382 367140 10542
rect 367284 9648 367336 9654
rect 367284 9590 367336 9596
rect 367296 9382 367324 9590
rect 367100 9376 367152 9382
rect 367100 9318 367152 9324
rect 367284 9376 367336 9382
rect 367284 9318 367336 9324
rect 367296 8566 367324 9318
rect 367284 8560 367336 8566
rect 367284 8502 367336 8508
rect 367480 8430 367508 11222
rect 368032 11014 368060 11222
rect 368020 11008 368072 11014
rect 368020 10950 368072 10956
rect 368572 9920 368624 9926
rect 368572 9862 368624 9868
rect 368584 9654 368612 9862
rect 368572 9648 368624 9654
rect 368572 9590 368624 9596
rect 367468 8424 367520 8430
rect 367468 8366 367520 8372
rect 367100 7948 367152 7954
rect 367100 7890 367152 7896
rect 366364 7812 366416 7818
rect 366364 7754 366416 7760
rect 367112 6322 367140 7890
rect 368480 7812 368532 7818
rect 368480 7754 368532 7760
rect 367928 6452 367980 6458
rect 367928 6394 367980 6400
rect 367100 6316 367152 6322
rect 367100 6258 367152 6264
rect 365812 3528 365864 3534
rect 365812 3470 365864 3476
rect 367100 2304 367152 2310
rect 367100 2246 367152 2252
rect 365628 1964 365680 1970
rect 365628 1906 365680 1912
rect 365076 1148 365128 1154
rect 365076 1090 365128 1096
rect 367112 1086 367140 2246
rect 367940 1494 367968 6394
rect 368492 6390 368520 7754
rect 368676 7546 368704 11222
rect 368940 11212 368992 11218
rect 368940 11154 368992 11160
rect 368952 10878 368980 11154
rect 368940 10872 368992 10878
rect 368940 10814 368992 10820
rect 368848 9580 368900 9586
rect 368848 9522 368900 9528
rect 368860 9382 368888 9522
rect 368848 9376 368900 9382
rect 368848 9318 368900 9324
rect 368664 7540 368716 7546
rect 368664 7482 368716 7488
rect 369780 7478 369808 11222
rect 370148 10538 370176 11222
rect 370136 10532 370188 10538
rect 370136 10474 370188 10480
rect 369768 7472 369820 7478
rect 369768 7414 369820 7420
rect 370700 7410 370728 11222
rect 371068 10470 371096 11222
rect 371056 10464 371108 10470
rect 371056 10406 371108 10412
rect 371332 9580 371384 9586
rect 371332 9522 371384 9528
rect 371056 9512 371108 9518
rect 371056 9454 371108 9460
rect 371068 9110 371096 9454
rect 371056 9104 371108 9110
rect 371056 9046 371108 9052
rect 371344 8838 371372 9522
rect 371332 8832 371384 8838
rect 371332 8774 371384 8780
rect 371804 8022 371832 11222
rect 372172 10402 372200 11222
rect 372160 10396 372212 10402
rect 372160 10338 372212 10344
rect 372712 9512 372764 9518
rect 372712 9454 372764 9460
rect 371792 8016 371844 8022
rect 371792 7958 371844 7964
rect 372528 8016 372580 8022
rect 372528 7958 372580 7964
rect 370780 7540 370832 7546
rect 370780 7482 370832 7488
rect 370688 7404 370740 7410
rect 370688 7346 370740 7352
rect 368480 6384 368532 6390
rect 368480 6326 368532 6332
rect 369952 6384 370004 6390
rect 369952 6326 370004 6332
rect 369860 6180 369912 6186
rect 369860 6122 369912 6128
rect 369872 2650 369900 6122
rect 369860 2644 369912 2650
rect 369860 2586 369912 2592
rect 369964 2514 369992 6326
rect 370792 5778 370820 7482
rect 372540 5914 372568 7958
rect 372528 5908 372580 5914
rect 372528 5850 372580 5856
rect 370780 5772 370832 5778
rect 370780 5714 370832 5720
rect 372620 3732 372672 3738
rect 372620 3674 372672 3680
rect 369952 2508 370004 2514
rect 369952 2450 370004 2456
rect 368388 2440 368440 2446
rect 368388 2382 368440 2388
rect 370964 2440 371016 2446
rect 370964 2382 371016 2388
rect 368400 2310 368428 2382
rect 370976 2310 371004 2382
rect 368388 2304 368440 2310
rect 368388 2246 368440 2252
rect 370964 2304 371016 2310
rect 370964 2246 371016 2252
rect 368400 1698 368428 2246
rect 368388 1692 368440 1698
rect 368388 1634 368440 1640
rect 370976 1494 371004 2246
rect 372632 1562 372660 3674
rect 372620 1556 372672 1562
rect 372620 1498 372672 1504
rect 367928 1488 367980 1494
rect 367928 1430 367980 1436
rect 370964 1488 371016 1494
rect 370964 1430 371016 1436
rect 372724 1358 372752 9454
rect 372908 7954 372936 11222
rect 373276 10334 373304 11222
rect 373264 10328 373316 10334
rect 373264 10270 373316 10276
rect 373540 9512 373592 9518
rect 373540 9454 373592 9460
rect 373552 9382 373580 9454
rect 373644 9450 373856 9466
rect 373632 9444 373868 9450
rect 373684 9438 373816 9444
rect 373632 9386 373684 9392
rect 373816 9386 373868 9392
rect 373540 9376 373592 9382
rect 373540 9318 373592 9324
rect 372896 7948 372948 7954
rect 372896 7890 372948 7896
rect 374012 7818 374040 11222
rect 374380 10266 374408 11222
rect 374460 10804 374512 10810
rect 374460 10746 374512 10752
rect 374472 10606 374500 10746
rect 374460 10600 374512 10606
rect 374460 10542 374512 10548
rect 374368 10260 374420 10266
rect 374368 10202 374420 10208
rect 374276 9580 374328 9586
rect 374276 9522 374328 9528
rect 374288 9382 374316 9522
rect 374276 9376 374328 9382
rect 374276 9318 374328 9324
rect 374288 9110 374316 9318
rect 374276 9104 374328 9110
rect 374276 9046 374328 9052
rect 374000 7812 374052 7818
rect 374000 7754 374052 7760
rect 374276 7812 374328 7818
rect 374276 7754 374328 7760
rect 373448 7472 373500 7478
rect 373448 7414 373500 7420
rect 372804 6792 372856 6798
rect 372804 6734 372856 6740
rect 372816 1766 372844 6734
rect 373460 5642 373488 7414
rect 373448 5636 373500 5642
rect 373448 5578 373500 5584
rect 374288 4078 374316 7754
rect 375116 7546 375144 11222
rect 375484 10198 375512 11222
rect 375472 10192 375524 10198
rect 375472 10134 375524 10140
rect 375932 9512 375984 9518
rect 375932 9454 375984 9460
rect 375944 9178 375972 9454
rect 375932 9172 375984 9178
rect 375932 9114 375984 9120
rect 376220 8022 376248 11222
rect 376852 10396 376904 10402
rect 376852 10338 376904 10344
rect 376760 9580 376812 9586
rect 376760 9522 376812 9528
rect 376772 9382 376800 9522
rect 376760 9376 376812 9382
rect 376760 9318 376812 9324
rect 376772 9178 376800 9318
rect 376760 9172 376812 9178
rect 376760 9114 376812 9120
rect 376864 8634 376892 10338
rect 376852 8628 376904 8634
rect 376852 8570 376904 8576
rect 376208 8016 376260 8022
rect 376208 7958 376260 7964
rect 375564 7948 375616 7954
rect 375564 7890 375616 7896
rect 375104 7540 375156 7546
rect 375104 7482 375156 7488
rect 375380 7540 375432 7546
rect 375380 7482 375432 7488
rect 375392 4146 375420 7482
rect 375380 4140 375432 4146
rect 375380 4082 375432 4088
rect 374276 4072 374328 4078
rect 374276 4014 374328 4020
rect 373540 2644 373592 2650
rect 373540 2586 373592 2592
rect 373448 2576 373500 2582
rect 373448 2518 373500 2524
rect 372804 1760 372856 1766
rect 372804 1702 372856 1708
rect 372712 1352 372764 1358
rect 372712 1294 372764 1300
rect 362592 1080 362644 1086
rect 362592 1022 362644 1028
rect 367100 1080 367152 1086
rect 367100 1022 367152 1028
rect 359924 1012 359976 1018
rect 359924 954 359976 960
rect 359832 876 359884 882
rect 359832 818 359884 824
rect 362604 814 362632 1022
rect 373460 814 373488 2518
rect 373552 1086 373580 2586
rect 375576 1426 375604 7890
rect 377048 6866 377076 11222
rect 377324 7478 377352 11222
rect 377600 10130 377628 11222
rect 378140 10464 378192 10470
rect 378140 10406 378192 10412
rect 377588 10124 377640 10130
rect 377588 10066 377640 10072
rect 378152 8566 378180 10406
rect 378324 9512 378376 9518
rect 378324 9454 378376 9460
rect 378336 8974 378364 9454
rect 378324 8968 378376 8974
rect 378324 8910 378376 8916
rect 378140 8560 378192 8566
rect 378140 8502 378192 8508
rect 378428 8090 378456 11222
rect 378704 10062 378732 11222
rect 378692 10056 378744 10062
rect 378692 9998 378744 10004
rect 379440 9994 379468 11222
rect 380360 10810 380388 11222
rect 380348 10804 380400 10810
rect 380348 10746 380400 10752
rect 381556 10742 381584 11222
rect 381544 10736 381596 10742
rect 381544 10678 381596 10684
rect 379980 10600 380032 10606
rect 379980 10542 380032 10548
rect 379428 9988 379480 9994
rect 379428 9930 379480 9936
rect 379244 9648 379296 9654
rect 379244 9590 379296 9596
rect 379152 9580 379204 9586
rect 379152 9522 379204 9528
rect 379164 9382 379192 9522
rect 379256 9382 379284 9590
rect 379992 9518 380020 10542
rect 382108 9722 382136 11222
rect 382476 10674 382504 11222
rect 382464 10668 382516 10674
rect 382464 10610 382516 10616
rect 383212 10402 383240 11222
rect 383568 11008 383620 11014
rect 383568 10950 383620 10956
rect 383200 10396 383252 10402
rect 383200 10338 383252 10344
rect 382188 10328 382240 10334
rect 382188 10270 382240 10276
rect 382096 9716 382148 9722
rect 382096 9658 382148 9664
rect 382200 9654 382228 10270
rect 382924 10260 382976 10266
rect 382924 10202 382976 10208
rect 382188 9648 382240 9654
rect 382188 9590 382240 9596
rect 379980 9512 380032 9518
rect 379980 9454 380032 9460
rect 380808 9512 380860 9518
rect 380808 9454 380860 9460
rect 379152 9376 379204 9382
rect 379152 9318 379204 9324
rect 379244 9376 379296 9382
rect 379244 9318 379296 9324
rect 379164 8634 379192 9318
rect 380820 9042 380848 9454
rect 380808 9036 380860 9042
rect 380808 8978 380860 8984
rect 382936 8838 382964 10202
rect 383016 9512 383068 9518
rect 383016 9454 383068 9460
rect 382924 8832 382976 8838
rect 382924 8774 382976 8780
rect 379152 8628 379204 8634
rect 379152 8570 379204 8576
rect 378416 8084 378468 8090
rect 378416 8026 378468 8032
rect 382280 8016 382332 8022
rect 382280 7958 382332 7964
rect 377312 7472 377364 7478
rect 377312 7414 377364 7420
rect 377036 6860 377088 6866
rect 377036 6802 377088 6808
rect 378140 6316 378192 6322
rect 378140 6258 378192 6264
rect 378152 2774 378180 6258
rect 381544 6248 381596 6254
rect 381544 6190 381596 6196
rect 378692 4072 378744 4078
rect 378692 4014 378744 4020
rect 378060 2746 378180 2774
rect 378060 2650 378088 2746
rect 376116 2644 376168 2650
rect 376116 2586 376168 2592
rect 378048 2644 378100 2650
rect 378048 2586 378100 2592
rect 378140 2644 378192 2650
rect 378140 2586 378192 2592
rect 376128 2446 376156 2586
rect 378152 2446 378180 2586
rect 376116 2440 376168 2446
rect 376116 2382 376168 2388
rect 378140 2440 378192 2446
rect 378140 2382 378192 2388
rect 376392 2304 376444 2310
rect 376392 2246 376444 2252
rect 377956 2304 378008 2310
rect 377956 2246 378008 2252
rect 375564 1420 375616 1426
rect 375564 1362 375616 1368
rect 376404 1154 376432 2246
rect 377968 2106 377996 2246
rect 377956 2100 378008 2106
rect 377956 2042 378008 2048
rect 378704 1834 378732 4014
rect 380900 2576 380952 2582
rect 380900 2518 380952 2524
rect 381084 2576 381136 2582
rect 381084 2518 381136 2524
rect 378692 1828 378744 1834
rect 378692 1770 378744 1776
rect 376392 1148 376444 1154
rect 376392 1090 376444 1096
rect 373540 1080 373592 1086
rect 373540 1022 373592 1028
rect 380912 814 380940 2518
rect 381096 2310 381124 2518
rect 381268 2440 381320 2446
rect 381268 2382 381320 2388
rect 381280 2310 381308 2382
rect 381084 2304 381136 2310
rect 381084 2246 381136 2252
rect 381268 2304 381320 2310
rect 381268 2246 381320 2252
rect 381280 1562 381308 2246
rect 381556 1766 381584 6190
rect 382292 1970 382320 7958
rect 382280 1964 382332 1970
rect 382280 1906 382332 1912
rect 381544 1760 381596 1766
rect 381544 1702 381596 1708
rect 381268 1556 381320 1562
rect 381268 1498 381320 1504
rect 383028 1222 383056 9454
rect 383580 8906 383608 10950
rect 384684 9382 384712 11222
rect 385236 10470 385264 11222
rect 385868 11144 385920 11150
rect 385868 11086 385920 11092
rect 385776 11076 385828 11082
rect 385776 11018 385828 11024
rect 385224 10464 385276 10470
rect 385224 10406 385276 10412
rect 385788 9450 385816 11018
rect 385776 9444 385828 9450
rect 385776 9386 385828 9392
rect 384672 9376 384724 9382
rect 384672 9318 384724 9324
rect 385880 9110 385908 11086
rect 385972 10334 386000 11222
rect 385960 10328 386012 10334
rect 385960 10270 386012 10276
rect 386524 10266 386552 11222
rect 387064 11144 387116 11150
rect 387064 11086 387116 11092
rect 386512 10260 386564 10266
rect 386512 10202 386564 10208
rect 385868 9104 385920 9110
rect 385868 9046 385920 9052
rect 383568 8900 383620 8906
rect 383568 8842 383620 8848
rect 387076 8634 387104 11086
rect 387996 9178 388024 11222
rect 388996 11212 389048 11218
rect 388996 11154 389048 11160
rect 389008 9654 389036 11154
rect 388996 9648 389048 9654
rect 388996 9590 389048 9596
rect 387984 9172 388036 9178
rect 387984 9114 388036 9120
rect 387064 8628 387116 8634
rect 387064 8570 387116 8576
rect 389180 5364 389232 5370
rect 389180 5306 389232 5312
rect 383200 2644 383252 2650
rect 383200 2586 383252 2592
rect 383292 2644 383344 2650
rect 383292 2586 383344 2592
rect 383844 2644 383896 2650
rect 383844 2586 383896 2592
rect 383212 2310 383240 2586
rect 383108 2304 383160 2310
rect 383108 2246 383160 2252
rect 383200 2304 383252 2310
rect 383200 2246 383252 2252
rect 383120 2038 383148 2246
rect 383304 2106 383332 2586
rect 383752 2304 383804 2310
rect 383752 2246 383804 2252
rect 383292 2100 383344 2106
rect 383292 2042 383344 2048
rect 383108 2032 383160 2038
rect 383108 1974 383160 1980
rect 383764 1970 383792 2246
rect 383752 1964 383804 1970
rect 383752 1906 383804 1912
rect 383016 1216 383068 1222
rect 383016 1158 383068 1164
rect 383856 814 383884 2586
rect 385040 2576 385092 2582
rect 385040 2518 385092 2524
rect 383936 2440 383988 2446
rect 383936 2382 383988 2388
rect 383948 2310 383976 2382
rect 383936 2304 383988 2310
rect 383936 2246 383988 2252
rect 383948 2106 383976 2246
rect 383936 2100 383988 2106
rect 383936 2042 383988 2048
rect 385052 814 385080 2518
rect 386420 2440 386472 2446
rect 386420 2382 386472 2388
rect 388996 2440 389048 2446
rect 388996 2382 389048 2388
rect 386432 2310 386460 2382
rect 389008 2310 389036 2382
rect 386420 2304 386472 2310
rect 386420 2246 386472 2252
rect 388996 2304 389048 2310
rect 388996 2246 389048 2252
rect 386432 1426 386460 2246
rect 387800 2032 387852 2038
rect 387800 1974 387852 1980
rect 386420 1420 386472 1426
rect 386420 1362 386472 1368
rect 387812 814 387840 1974
rect 389008 1834 389036 2246
rect 388996 1828 389048 1834
rect 388996 1770 389048 1776
rect 389192 1630 389220 5306
rect 389836 4826 389864 11222
rect 390560 11008 390612 11014
rect 390560 10950 390612 10956
rect 390572 5234 390600 10950
rect 390560 5228 390612 5234
rect 390560 5170 390612 5176
rect 390664 5098 390692 11222
rect 391400 5166 391428 11222
rect 391952 5302 391980 11222
rect 392124 8084 392176 8090
rect 392124 8026 392176 8032
rect 391940 5296 391992 5302
rect 391940 5238 391992 5244
rect 391388 5160 391440 5166
rect 391388 5102 391440 5108
rect 390652 5092 390704 5098
rect 390652 5034 390704 5040
rect 389824 4820 389876 4826
rect 389824 4762 389876 4768
rect 390560 4820 390612 4826
rect 390560 4762 390612 4768
rect 390572 2417 390600 4762
rect 392136 3602 392164 8026
rect 392504 4758 392532 11222
rect 392872 7886 392900 11222
rect 392860 7880 392912 7886
rect 392860 7822 392912 7828
rect 393516 7818 393544 11222
rect 393504 7812 393556 7818
rect 393504 7754 393556 7760
rect 393964 7812 394016 7818
rect 393964 7754 394016 7760
rect 392492 4752 392544 4758
rect 392492 4694 392544 4700
rect 392124 3596 392176 3602
rect 392124 3538 392176 3544
rect 390652 2644 390704 2650
rect 390652 2586 390704 2592
rect 390558 2408 390614 2417
rect 390558 2343 390614 2352
rect 389180 1624 389232 1630
rect 389180 1566 389232 1572
rect 390664 814 390692 2586
rect 391940 2576 391992 2582
rect 391940 2518 391992 2524
rect 392032 2576 392084 2582
rect 392032 2518 392084 2524
rect 393320 2576 393372 2582
rect 393976 2553 394004 7754
rect 394068 7546 394096 11222
rect 394712 8090 394740 11222
rect 394700 8084 394752 8090
rect 394700 8026 394752 8032
rect 394056 7540 394108 7546
rect 394056 7482 394108 7488
rect 395172 3670 395200 11222
rect 395540 4690 395568 11222
rect 396080 11008 396132 11014
rect 396080 10950 396132 10956
rect 396092 6730 396120 10950
rect 396080 6724 396132 6730
rect 396080 6666 396132 6672
rect 395528 4684 395580 4690
rect 395528 4626 395580 4632
rect 395160 3664 395212 3670
rect 395160 3606 395212 3612
rect 395436 3528 395488 3534
rect 395436 3470 395488 3476
rect 394056 2644 394108 2650
rect 394056 2586 394108 2592
rect 393320 2518 393372 2524
rect 393962 2544 394018 2553
rect 391572 2440 391624 2446
rect 391572 2382 391624 2388
rect 391584 2310 391612 2382
rect 391572 2304 391624 2310
rect 391572 2246 391624 2252
rect 391584 2038 391612 2246
rect 391572 2032 391624 2038
rect 391572 1974 391624 1980
rect 391952 814 391980 2518
rect 392044 1970 392072 2518
rect 393332 2446 393360 2518
rect 393962 2479 394018 2488
rect 393320 2440 393372 2446
rect 393320 2382 393372 2388
rect 392032 1964 392084 1970
rect 392032 1906 392084 1912
rect 394068 814 394096 2586
rect 395252 2576 395304 2582
rect 395252 2518 395304 2524
rect 394148 2440 394200 2446
rect 394148 2382 394200 2388
rect 394160 1766 394188 2382
rect 394148 1760 394200 1766
rect 394148 1702 394200 1708
rect 395264 814 395292 2518
rect 395448 1494 395476 3470
rect 396276 3194 396304 11222
rect 397460 11008 397512 11014
rect 397460 10950 397512 10956
rect 397472 4010 397500 10950
rect 397932 6458 397960 11222
rect 397920 6452 397972 6458
rect 397920 6394 397972 6400
rect 398484 4622 398512 11222
rect 399300 11144 399352 11150
rect 399300 11086 399352 11092
rect 399852 11144 399904 11150
rect 399852 11086 399904 11092
rect 398840 6452 398892 6458
rect 398840 6394 398892 6400
rect 398472 4616 398524 4622
rect 398472 4558 398524 4564
rect 397460 4004 397512 4010
rect 397460 3946 397512 3952
rect 397368 3460 397420 3466
rect 397368 3402 397420 3408
rect 396264 3188 396316 3194
rect 396264 3130 396316 3136
rect 396724 2440 396776 2446
rect 396724 2382 396776 2388
rect 396736 1630 396764 2382
rect 397380 2106 397408 3402
rect 398748 2644 398800 2650
rect 398748 2586 398800 2592
rect 397644 2576 397696 2582
rect 397644 2518 397696 2524
rect 397368 2100 397420 2106
rect 397368 2042 397420 2048
rect 396724 1624 396776 1630
rect 396724 1566 396776 1572
rect 395436 1488 395488 1494
rect 395436 1430 395488 1436
rect 397656 814 397684 2518
rect 398760 2446 398788 2586
rect 398748 2440 398800 2446
rect 398748 2382 398800 2388
rect 398852 2310 398880 6394
rect 399312 3738 399340 11086
rect 399864 6390 399892 11086
rect 400312 11008 400364 11014
rect 400312 10950 400364 10956
rect 400324 6662 400352 10950
rect 400692 7954 400720 11222
rect 400968 8294 400996 11222
rect 401968 11008 402020 11014
rect 401968 10950 402020 10956
rect 400956 8288 401008 8294
rect 400956 8230 401008 8236
rect 400680 7948 400732 7954
rect 400680 7890 400732 7896
rect 401980 6798 402008 10950
rect 402348 8022 402376 11222
rect 403072 11008 403124 11014
rect 403072 10950 403124 10956
rect 403624 11008 403676 11014
rect 403624 10950 403676 10956
rect 402336 8016 402388 8022
rect 402336 7958 402388 7964
rect 401968 6792 402020 6798
rect 401968 6734 402020 6740
rect 400312 6656 400364 6662
rect 400312 6598 400364 6604
rect 399852 6384 399904 6390
rect 399852 6326 399904 6332
rect 400312 6384 400364 6390
rect 400312 6326 400364 6332
rect 399300 3732 399352 3738
rect 399300 3674 399352 3680
rect 400220 2576 400272 2582
rect 400220 2518 400272 2524
rect 398840 2304 398892 2310
rect 398840 2246 398892 2252
rect 400232 814 400260 2518
rect 400324 2514 400352 6326
rect 400404 5160 400456 5166
rect 400404 5102 400456 5108
rect 400312 2508 400364 2514
rect 400312 2450 400364 2456
rect 400416 1698 400444 5102
rect 403084 4078 403112 10950
rect 403636 5370 403664 10950
rect 403912 7750 403940 11222
rect 430212 8288 430264 8294
rect 430212 8230 430264 8236
rect 426164 8016 426216 8022
rect 426164 7958 426216 7964
rect 419908 7880 419960 7886
rect 419908 7822 419960 7828
rect 403900 7744 403952 7750
rect 403900 7686 403952 7692
rect 414756 7744 414808 7750
rect 414756 7686 414808 7692
rect 408500 6656 408552 6662
rect 408500 6598 408552 6604
rect 403624 5364 403676 5370
rect 403624 5306 403676 5312
rect 403992 5228 404044 5234
rect 403992 5170 404044 5176
rect 403072 4072 403124 4078
rect 403072 4014 403124 4020
rect 404004 2378 404032 5170
rect 404360 5092 404412 5098
rect 404360 5034 404412 5040
rect 404372 2582 404400 5034
rect 408512 2650 408540 6598
rect 408500 2644 408552 2650
rect 408500 2586 408552 2592
rect 414768 2582 414796 7686
rect 417056 5296 417108 5302
rect 417056 5238 417108 5244
rect 404360 2576 404412 2582
rect 404360 2518 404412 2524
rect 414756 2576 414808 2582
rect 414756 2518 414808 2524
rect 404372 2446 404400 2518
rect 404360 2440 404412 2446
rect 404360 2382 404412 2388
rect 403992 2372 404044 2378
rect 403992 2314 404044 2320
rect 402428 2304 402480 2310
rect 402428 2246 402480 2252
rect 405924 2304 405976 2310
rect 405924 2246 405976 2252
rect 406292 2304 406344 2310
rect 406292 2246 406344 2252
rect 407028 2304 407080 2310
rect 407028 2246 407080 2252
rect 408868 2304 408920 2310
rect 408868 2246 408920 2252
rect 409604 2304 409656 2310
rect 409604 2246 409656 2252
rect 411444 2304 411496 2310
rect 411444 2246 411496 2252
rect 414020 2304 414072 2310
rect 414020 2246 414072 2252
rect 416504 2304 416556 2310
rect 416504 2246 416556 2252
rect 400404 1692 400456 1698
rect 400404 1634 400456 1640
rect 402440 814 402468 2246
rect 355416 808 355468 814
rect 355416 750 355468 756
rect 362592 808 362644 814
rect 362592 750 362644 756
rect 373448 808 373500 814
rect 373448 750 373500 756
rect 380900 808 380952 814
rect 380900 750 380952 756
rect 383844 808 383896 814
rect 383844 750 383896 756
rect 385040 808 385092 814
rect 385040 750 385092 756
rect 387800 808 387852 814
rect 387800 750 387852 756
rect 390652 808 390704 814
rect 390652 750 390704 756
rect 391940 808 391992 814
rect 391940 750 391992 756
rect 394056 808 394108 814
rect 394056 750 394108 756
rect 395252 808 395304 814
rect 395252 750 395304 756
rect 397644 808 397696 814
rect 397644 750 397696 756
rect 400220 808 400272 814
rect 400220 750 400272 756
rect 402428 808 402480 814
rect 402428 750 402480 756
rect 405936 746 405964 2246
rect 406304 814 406332 2246
rect 407040 1494 407068 2246
rect 407028 1488 407080 1494
rect 407028 1430 407080 1436
rect 408880 814 408908 2246
rect 409616 2106 409644 2246
rect 409604 2100 409656 2106
rect 409604 2042 409656 2048
rect 411456 814 411484 2246
rect 414032 814 414060 2246
rect 416516 814 416544 2246
rect 417068 1562 417096 5238
rect 419920 2582 419948 7822
rect 420920 3664 420972 3670
rect 420920 3606 420972 3612
rect 419908 2576 419960 2582
rect 419908 2518 419960 2524
rect 417332 2440 417384 2446
rect 417332 2382 417384 2388
rect 417344 2310 417372 2382
rect 417332 2304 417384 2310
rect 417332 2246 417384 2252
rect 419172 2304 419224 2310
rect 419172 2246 419224 2252
rect 417344 1970 417372 2246
rect 417332 1964 417384 1970
rect 417332 1906 417384 1912
rect 417056 1556 417108 1562
rect 417056 1498 417108 1504
rect 419184 814 419212 2246
rect 420932 2038 420960 3606
rect 426176 2582 426204 7958
rect 426992 5364 427044 5370
rect 426992 5306 427044 5312
rect 426164 2576 426216 2582
rect 426164 2518 426216 2524
rect 422484 2440 422536 2446
rect 422484 2382 422536 2388
rect 422496 2310 422524 2382
rect 421748 2304 421800 2310
rect 421748 2246 421800 2252
rect 422484 2304 422536 2310
rect 422484 2246 422536 2252
rect 423588 2304 423640 2310
rect 423588 2246 423640 2252
rect 426072 2304 426124 2310
rect 426072 2246 426124 2252
rect 420920 2032 420972 2038
rect 420920 1974 420972 1980
rect 421760 814 421788 2246
rect 422496 2038 422524 2246
rect 422484 2032 422536 2038
rect 422484 1974 422536 1980
rect 423600 814 423628 2246
rect 426084 814 426112 2246
rect 427004 1426 427032 5306
rect 430224 2582 430252 8230
rect 432052 6724 432104 6730
rect 432052 6666 432104 6672
rect 430212 2576 430264 2582
rect 430212 2518 430264 2524
rect 431776 2576 431828 2582
rect 431776 2518 431828 2524
rect 427636 2440 427688 2446
rect 427636 2382 427688 2388
rect 427648 2310 427676 2382
rect 427636 2304 427688 2310
rect 427636 2246 427688 2252
rect 427728 2304 427780 2310
rect 427728 2246 427780 2252
rect 430488 2304 430540 2310
rect 430488 2246 430540 2252
rect 427648 1698 427676 2246
rect 427636 1692 427688 1698
rect 427636 1634 427688 1640
rect 426992 1420 427044 1426
rect 426992 1362 427044 1368
rect 427740 814 427768 2246
rect 430500 814 430528 2246
rect 431788 814 431816 2518
rect 432064 1834 432092 6666
rect 438872 4826 438900 11222
rect 440160 7818 440188 11222
rect 440332 11076 440384 11082
rect 440332 11018 440384 11024
rect 440240 11008 440292 11014
rect 440240 10950 440292 10956
rect 440148 7812 440200 7818
rect 440148 7754 440200 7760
rect 440252 6458 440280 10950
rect 440240 6452 440292 6458
rect 440240 6394 440292 6400
rect 440344 5098 440372 11018
rect 439136 5092 439188 5098
rect 439136 5034 439188 5040
rect 440332 5092 440384 5098
rect 440332 5034 440384 5040
rect 439148 4826 439176 5034
rect 440148 5024 440200 5030
rect 440148 4966 440200 4972
rect 438860 4820 438912 4826
rect 438860 4762 438912 4768
rect 439136 4820 439188 4826
rect 439136 4762 439188 4768
rect 435364 3596 435416 3602
rect 435364 3538 435416 3544
rect 435376 2582 435404 3538
rect 435364 2576 435416 2582
rect 435364 2518 435416 2524
rect 436836 2576 436888 2582
rect 436836 2518 436888 2524
rect 432788 2440 432840 2446
rect 432788 2382 432840 2388
rect 432800 2310 432828 2382
rect 432788 2304 432840 2310
rect 432788 2246 432840 2252
rect 434628 2304 434680 2310
rect 434628 2246 434680 2252
rect 432052 1828 432104 1834
rect 432052 1770 432104 1776
rect 432800 1562 432828 2246
rect 432788 1556 432840 1562
rect 432788 1498 432840 1504
rect 434640 814 434668 2246
rect 436848 814 436876 2518
rect 440160 1766 440188 4966
rect 440240 4140 440292 4146
rect 440240 4082 440292 4088
rect 440252 2378 440280 4082
rect 440436 3942 440464 11222
rect 440712 6254 440740 11222
rect 441620 11008 441672 11014
rect 441620 10950 441672 10956
rect 440976 6860 441028 6866
rect 440976 6802 441028 6808
rect 440700 6248 440752 6254
rect 440700 6190 440752 6196
rect 440424 3936 440476 3942
rect 440424 3878 440476 3884
rect 440240 2372 440292 2378
rect 440240 2314 440292 2320
rect 440516 2304 440568 2310
rect 440516 2246 440568 2252
rect 440528 1766 440556 2246
rect 440148 1760 440200 1766
rect 440148 1702 440200 1708
rect 440516 1760 440568 1766
rect 440516 1702 440568 1708
rect 440988 1630 441016 6802
rect 441632 6186 441660 10950
rect 441712 10940 441764 10946
rect 441712 10882 441764 10888
rect 441724 6390 441752 10882
rect 441712 6384 441764 6390
rect 441712 6326 441764 6332
rect 441620 6180 441672 6186
rect 441620 6122 441672 6128
rect 441816 5166 441844 11290
rect 442080 11008 442132 11014
rect 442080 10950 442132 10956
rect 442632 11008 442684 11014
rect 442632 10950 442684 10956
rect 441804 5160 441856 5166
rect 441804 5102 441856 5108
rect 442092 3534 442120 10950
rect 442644 6322 442672 10950
rect 442920 8378 442948 11290
rect 443184 11280 443236 11286
rect 443184 11222 443236 11228
rect 443460 11280 443512 11286
rect 443460 11222 443512 11228
rect 444012 11280 444064 11286
rect 444012 11222 444064 11228
rect 444564 11280 444616 11286
rect 444564 11222 444616 11228
rect 444748 11280 444800 11286
rect 444748 11222 444800 11228
rect 445024 11280 445076 11286
rect 445024 11222 445076 11228
rect 445300 11280 445352 11286
rect 445300 11222 445352 11228
rect 443092 11008 443144 11014
rect 443092 10950 443144 10956
rect 442920 8350 443040 8378
rect 442908 6384 442960 6390
rect 442908 6326 442960 6332
rect 442632 6316 442684 6322
rect 442632 6258 442684 6264
rect 442080 3528 442132 3534
rect 442080 3470 442132 3476
rect 442356 2304 442408 2310
rect 442356 2246 442408 2252
rect 440976 1624 441028 1630
rect 440976 1566 441028 1572
rect 442368 1086 442396 2246
rect 442920 1494 442948 6326
rect 443012 5234 443040 8350
rect 443104 5370 443132 10950
rect 443092 5364 443144 5370
rect 443092 5306 443144 5312
rect 443196 5302 443224 11222
rect 443184 5296 443236 5302
rect 443184 5238 443236 5244
rect 443000 5228 443052 5234
rect 443000 5170 443052 5176
rect 443472 3466 443500 11222
rect 444024 6730 444052 11222
rect 444380 10940 444432 10946
rect 444380 10882 444432 10888
rect 444012 6724 444064 6730
rect 444012 6666 444064 6672
rect 443736 5364 443788 5370
rect 443736 5306 443788 5312
rect 443460 3460 443512 3466
rect 443460 3402 443512 3408
rect 443092 2304 443144 2310
rect 443092 2246 443144 2252
rect 443104 1902 443132 2246
rect 443748 2106 443776 5306
rect 444392 3670 444420 10882
rect 444576 5030 444604 11222
rect 444760 6866 444788 11222
rect 444748 6860 444800 6866
rect 444748 6802 444800 6808
rect 445036 6662 445064 11222
rect 445024 6656 445076 6662
rect 445024 6598 445076 6604
rect 444564 5024 444616 5030
rect 444564 4966 444616 4972
rect 445312 4146 445340 11222
rect 445576 8084 445628 8090
rect 445576 8026 445628 8032
rect 445300 4140 445352 4146
rect 445300 4082 445352 4088
rect 444380 3664 444432 3670
rect 444380 3606 444432 3612
rect 444380 2304 444432 2310
rect 444380 2246 444432 2252
rect 443736 2100 443788 2106
rect 443736 2042 443788 2048
rect 443092 1896 443144 1902
rect 443092 1838 443144 1844
rect 442908 1488 442960 1494
rect 442908 1430 442960 1436
rect 442356 1080 442408 1086
rect 442356 1022 442408 1028
rect 444392 950 444420 2246
rect 445588 1698 445616 8026
rect 445668 6180 445720 6186
rect 445668 6122 445720 6128
rect 445680 2514 445708 6122
rect 445772 4826 445800 11342
rect 445852 11280 445904 11286
rect 445852 11222 445904 11228
rect 446128 11280 446180 11286
rect 446128 11222 446180 11228
rect 445864 6390 445892 11222
rect 445852 6384 445904 6390
rect 445852 6326 445904 6332
rect 446140 5370 446168 11222
rect 446128 5364 446180 5370
rect 446128 5306 446180 5312
rect 445760 4820 445812 4826
rect 445760 4762 445812 4768
rect 446600 2650 446628 11478
rect 446680 11348 446732 11354
rect 446680 11290 446732 11296
rect 447784 11348 447836 11354
rect 447784 11290 447836 11296
rect 448060 11348 448112 11354
rect 448060 11290 448112 11296
rect 462692 11300 463012 11972
rect 446692 7750 446720 11290
rect 447140 11008 447192 11014
rect 447140 10950 447192 10956
rect 447692 11008 447744 11014
rect 447692 10950 447744 10956
rect 447048 8288 447100 8294
rect 447048 8230 447100 8236
rect 447060 8090 447088 8230
rect 447048 8084 447100 8090
rect 447048 8026 447100 8032
rect 446680 7744 446732 7750
rect 446680 7686 446732 7692
rect 446588 2644 446640 2650
rect 446588 2586 446640 2592
rect 445668 2508 445720 2514
rect 445668 2450 445720 2456
rect 445760 2304 445812 2310
rect 445760 2246 445812 2252
rect 445576 1692 445628 1698
rect 445576 1634 445628 1640
rect 444380 944 444432 950
rect 444380 886 444432 892
rect 445772 882 445800 2246
rect 447152 1970 447180 10950
rect 447232 10940 447284 10946
rect 447232 10882 447284 10888
rect 447244 7886 447272 10882
rect 447232 7880 447284 7886
rect 447232 7822 447284 7828
rect 447704 2038 447732 10950
rect 447796 8022 447824 11290
rect 448072 8294 448100 11290
rect 462692 11244 462704 11300
rect 462760 11244 462784 11300
rect 462840 11244 462864 11300
rect 462920 11244 462944 11300
rect 463000 11244 463012 11300
rect 462692 11220 463012 11244
rect 462692 11164 462704 11220
rect 462760 11164 462784 11220
rect 462840 11164 462864 11220
rect 462920 11164 462944 11220
rect 463000 11164 463012 11220
rect 462692 11140 463012 11164
rect 462692 11084 462704 11140
rect 462760 11084 462784 11140
rect 462840 11084 462864 11140
rect 462920 11084 462944 11140
rect 463000 11084 463012 11140
rect 462692 11060 463012 11084
rect 462692 11004 462704 11060
rect 462760 11004 462784 11060
rect 462840 11004 462864 11060
rect 462920 11004 462944 11060
rect 463000 11004 463012 11060
rect 448336 10940 448388 10946
rect 448336 10882 448388 10888
rect 448348 8362 448376 10882
rect 462692 9274 463012 11004
rect 462692 9222 462698 9274
rect 462750 9222 462762 9274
rect 462814 9222 462826 9274
rect 462878 9222 462890 9274
rect 462942 9222 462954 9274
rect 463006 9222 463012 9274
rect 462692 8988 463012 9222
rect 462692 8932 462704 8988
rect 462760 8932 462784 8988
rect 462840 8932 462864 8988
rect 462920 8932 462944 8988
rect 463000 8932 463012 8988
rect 462692 8908 463012 8932
rect 462692 8852 462704 8908
rect 462760 8852 462784 8908
rect 462840 8852 462864 8908
rect 462920 8852 462944 8908
rect 463000 8852 463012 8908
rect 462692 8828 463012 8852
rect 462692 8772 462704 8828
rect 462760 8772 462784 8828
rect 462840 8772 462864 8828
rect 462920 8772 462944 8828
rect 463000 8772 463012 8828
rect 462692 8748 463012 8772
rect 462692 8692 462704 8748
rect 462760 8692 462784 8748
rect 462840 8692 462864 8748
rect 462920 8692 462944 8748
rect 463000 8692 463012 8748
rect 448336 8356 448388 8362
rect 448336 8298 448388 8304
rect 448060 8288 448112 8294
rect 448060 8230 448112 8236
rect 462692 8186 463012 8692
rect 462692 8134 462698 8186
rect 462750 8134 462762 8186
rect 462814 8134 462826 8186
rect 462878 8134 462890 8186
rect 462942 8134 462954 8186
rect 463006 8134 463012 8186
rect 447784 8016 447836 8022
rect 447784 7958 447836 7964
rect 462692 7098 463012 8134
rect 462692 7046 462698 7098
rect 462750 7084 462762 7098
rect 462814 7084 462826 7098
rect 462878 7084 462890 7098
rect 462942 7084 462954 7098
rect 462760 7046 462762 7084
rect 462942 7046 462944 7084
rect 463006 7046 463012 7098
rect 462692 7028 462704 7046
rect 462760 7028 462784 7046
rect 462840 7028 462864 7046
rect 462920 7028 462944 7046
rect 463000 7028 463012 7046
rect 462692 7004 463012 7028
rect 462692 6948 462704 7004
rect 462760 6948 462784 7004
rect 462840 6948 462864 7004
rect 462920 6948 462944 7004
rect 463000 6948 463012 7004
rect 462692 6924 463012 6948
rect 462692 6868 462704 6924
rect 462760 6868 462784 6924
rect 462840 6868 462864 6924
rect 462920 6868 462944 6924
rect 463000 6868 463012 6924
rect 462692 6844 463012 6868
rect 462692 6788 462704 6844
rect 462760 6788 462784 6844
rect 462840 6788 462864 6844
rect 462920 6788 462944 6844
rect 463000 6788 463012 6844
rect 459560 6248 459612 6254
rect 459560 6190 459612 6196
rect 456800 5024 456852 5030
rect 456800 4966 456852 4972
rect 450820 4820 450872 4826
rect 450820 4762 450872 4768
rect 450832 2650 450860 4762
rect 455972 3460 456024 3466
rect 455972 3402 456024 3408
rect 450820 2644 450872 2650
rect 450820 2586 450872 2592
rect 450832 2446 450860 2586
rect 455420 2576 455472 2582
rect 455420 2518 455472 2524
rect 450820 2440 450872 2446
rect 450820 2382 450872 2388
rect 448244 2304 448296 2310
rect 448244 2246 448296 2252
rect 448520 2304 448572 2310
rect 448520 2246 448572 2252
rect 451372 2304 451424 2310
rect 451372 2246 451424 2252
rect 453396 2304 453448 2310
rect 453396 2246 453448 2252
rect 447692 2032 447744 2038
rect 447692 1974 447744 1980
rect 447140 1964 447192 1970
rect 447140 1906 447192 1912
rect 448256 1698 448284 2246
rect 448244 1692 448296 1698
rect 448244 1634 448296 1640
rect 448532 1290 448560 2246
rect 448520 1284 448572 1290
rect 448520 1226 448572 1232
rect 451384 1222 451412 2246
rect 451372 1216 451424 1222
rect 451372 1158 451424 1164
rect 453408 1154 453436 2246
rect 453396 1148 453448 1154
rect 453396 1090 453448 1096
rect 455432 882 455460 2518
rect 455984 2446 456012 3402
rect 455972 2440 456024 2446
rect 455972 2382 456024 2388
rect 456812 1562 456840 4966
rect 459572 2514 459600 6190
rect 462692 6010 463012 6788
rect 462692 5958 462698 6010
rect 462750 5958 462762 6010
rect 462814 5958 462826 6010
rect 462878 5958 462890 6010
rect 462942 5958 462954 6010
rect 463006 5958 463012 6010
rect 462692 5180 463012 5958
rect 462692 5124 462704 5180
rect 462760 5124 462784 5180
rect 462840 5124 462864 5180
rect 462920 5124 462944 5180
rect 463000 5124 463012 5180
rect 462692 5100 463012 5124
rect 462692 5044 462704 5100
rect 462760 5044 462784 5100
rect 462840 5044 462864 5100
rect 462920 5044 462944 5100
rect 463000 5044 463012 5100
rect 462692 5020 463012 5044
rect 462692 4964 462704 5020
rect 462760 4964 462784 5020
rect 462840 4964 462864 5020
rect 462920 4964 462944 5020
rect 463000 4964 463012 5020
rect 462692 4940 463012 4964
rect 462692 4922 462704 4940
rect 462760 4922 462784 4940
rect 462840 4922 462864 4940
rect 462920 4922 462944 4940
rect 463000 4922 463012 4940
rect 462692 4870 462698 4922
rect 462760 4884 462762 4922
rect 462942 4884 462944 4922
rect 462750 4870 462762 4884
rect 462814 4870 462826 4884
rect 462878 4870 462890 4884
rect 462942 4870 462954 4884
rect 463006 4870 463012 4922
rect 462692 3834 463012 4870
rect 462692 3782 462698 3834
rect 462750 3782 462762 3834
rect 462814 3782 462826 3834
rect 462878 3782 462890 3834
rect 462942 3782 462954 3834
rect 463006 3782 463012 3834
rect 462692 3276 463012 3782
rect 462692 3220 462704 3276
rect 462760 3220 462784 3276
rect 462840 3220 462864 3276
rect 462920 3220 462944 3276
rect 463000 3220 463012 3276
rect 462692 3196 463012 3220
rect 462692 3140 462704 3196
rect 462760 3140 462784 3196
rect 462840 3140 462864 3196
rect 462920 3140 462944 3196
rect 463000 3140 463012 3196
rect 462692 3116 463012 3140
rect 462692 3060 462704 3116
rect 462760 3060 462784 3116
rect 462840 3060 462864 3116
rect 462920 3060 462944 3116
rect 463000 3060 463012 3116
rect 462692 3036 463012 3060
rect 462692 2980 462704 3036
rect 462760 2980 462784 3036
rect 462840 2980 462864 3036
rect 462920 2980 462944 3036
rect 463000 2980 463012 3036
rect 462692 2746 463012 2980
rect 462692 2694 462698 2746
rect 462750 2694 462762 2746
rect 462814 2694 462826 2746
rect 462878 2694 462890 2746
rect 462942 2694 462954 2746
rect 463006 2694 463012 2746
rect 459560 2508 459612 2514
rect 459560 2450 459612 2456
rect 460388 2304 460440 2310
rect 460388 2246 460440 2252
rect 462320 2304 462372 2310
rect 462320 2246 462372 2252
rect 456800 1556 456852 1562
rect 456800 1498 456852 1504
rect 460400 1358 460428 2246
rect 460388 1352 460440 1358
rect 460388 1294 460440 1300
rect 462332 1290 462360 2246
rect 462320 1284 462372 1290
rect 462320 1226 462372 1232
rect 462692 964 463012 2694
rect 462692 908 462704 964
rect 462760 908 462784 964
rect 462840 908 462864 964
rect 462920 908 462944 964
rect 463000 908 463012 964
rect 462692 884 463012 908
rect 445760 876 445812 882
rect 445760 818 445812 824
rect 455420 876 455472 882
rect 455420 818 455472 824
rect 462692 828 462704 884
rect 462760 828 462784 884
rect 462840 828 462864 884
rect 462920 828 462944 884
rect 463000 828 463012 884
rect 406292 808 406344 814
rect 406292 750 406344 756
rect 408868 808 408920 814
rect 408868 750 408920 756
rect 411444 808 411496 814
rect 411444 750 411496 756
rect 414020 808 414072 814
rect 414020 750 414072 756
rect 416504 808 416556 814
rect 416504 750 416556 756
rect 419172 808 419224 814
rect 419172 750 419224 756
rect 421748 808 421800 814
rect 421748 750 421800 756
rect 423588 808 423640 814
rect 423588 750 423640 756
rect 426072 808 426124 814
rect 426072 750 426124 756
rect 427728 808 427780 814
rect 427728 750 427780 756
rect 430488 808 430540 814
rect 430488 750 430540 756
rect 431776 808 431828 814
rect 431776 750 431828 756
rect 434628 808 434680 814
rect 434628 750 434680 756
rect 436836 808 436888 814
rect 436836 750 436888 756
rect 462692 804 463012 828
rect 462692 748 462704 804
rect 462760 748 462784 804
rect 462840 748 462864 804
rect 462920 748 462944 804
rect 463000 748 463012 804
rect 405924 740 405976 746
rect 405924 682 405976 688
rect 462692 724 463012 748
rect 462692 668 462704 724
rect 462760 668 462784 724
rect 462840 668 462864 724
rect 462920 668 462944 724
rect 463000 668 463012 724
rect 347044 128 347096 134
rect 347044 70 347096 76
rect 331424 8 331436 64
rect 331492 8 331516 64
rect 331572 8 331596 64
rect 331652 8 331676 64
rect 331732 8 331744 64
rect 331424 -4 331744 8
rect 344468 60 344520 66
rect 344468 2 344520 8
rect 462692 -4 463012 668
rect 463352 11960 463672 11972
rect 463352 11904 463364 11960
rect 463420 11904 463444 11960
rect 463500 11904 463524 11960
rect 463580 11904 463604 11960
rect 463660 11904 463672 11960
rect 463352 11880 463672 11904
rect 463352 11824 463364 11880
rect 463420 11824 463444 11880
rect 463500 11824 463524 11880
rect 463580 11824 463604 11880
rect 463660 11824 463672 11880
rect 463352 11800 463672 11824
rect 463352 11744 463364 11800
rect 463420 11744 463444 11800
rect 463500 11744 463524 11800
rect 463580 11744 463604 11800
rect 463660 11744 463672 11800
rect 463352 11720 463672 11744
rect 463352 11664 463364 11720
rect 463420 11664 463444 11720
rect 463500 11664 463524 11720
rect 463580 11664 463604 11720
rect 463660 11664 463672 11720
rect 463352 9818 463672 11664
rect 530676 11960 530996 11972
rect 530676 11904 530688 11960
rect 530744 11904 530768 11960
rect 530824 11904 530848 11960
rect 530904 11904 530928 11960
rect 530984 11904 530996 11960
rect 530676 11880 530996 11904
rect 530676 11824 530688 11880
rect 530744 11824 530768 11880
rect 530824 11824 530848 11880
rect 530904 11824 530928 11880
rect 530984 11824 530996 11880
rect 530676 11800 530996 11824
rect 530676 11744 530688 11800
rect 530744 11744 530768 11800
rect 530824 11744 530848 11800
rect 530904 11744 530928 11800
rect 530984 11744 530996 11800
rect 530676 11720 530996 11744
rect 530676 11664 530688 11720
rect 530744 11664 530768 11720
rect 530824 11664 530848 11720
rect 530904 11664 530928 11720
rect 530984 11664 530996 11720
rect 483664 11416 483716 11422
rect 483584 11364 483664 11370
rect 483584 11358 483716 11364
rect 481824 11348 481876 11354
rect 481824 11290 481876 11296
rect 482836 11348 482888 11354
rect 482836 11290 482888 11296
rect 483112 11348 483164 11354
rect 483112 11290 483164 11296
rect 483584 11342 483704 11358
rect 484492 11348 484544 11354
rect 480720 11280 480772 11286
rect 480720 11222 480772 11228
rect 481272 11280 481324 11286
rect 481272 11222 481324 11228
rect 478880 11008 478932 11014
rect 478880 10950 478932 10956
rect 480352 11008 480404 11014
rect 480352 10950 480404 10956
rect 463352 9766 463358 9818
rect 463410 9766 463422 9818
rect 463474 9766 463486 9818
rect 463538 9766 463550 9818
rect 463602 9766 463614 9818
rect 463666 9766 463672 9818
rect 463352 9648 463672 9766
rect 463352 9592 463364 9648
rect 463420 9592 463444 9648
rect 463500 9592 463524 9648
rect 463580 9592 463604 9648
rect 463660 9592 463672 9648
rect 463352 9568 463672 9592
rect 463352 9512 463364 9568
rect 463420 9512 463444 9568
rect 463500 9512 463524 9568
rect 463580 9512 463604 9568
rect 463660 9512 463672 9568
rect 463352 9488 463672 9512
rect 463352 9432 463364 9488
rect 463420 9432 463444 9488
rect 463500 9432 463524 9488
rect 463580 9432 463604 9488
rect 463660 9432 463672 9488
rect 463352 9408 463672 9432
rect 463352 9352 463364 9408
rect 463420 9352 463444 9408
rect 463500 9352 463524 9408
rect 463580 9352 463604 9408
rect 463660 9352 463672 9408
rect 463352 8730 463672 9352
rect 463352 8678 463358 8730
rect 463410 8678 463422 8730
rect 463474 8678 463486 8730
rect 463538 8678 463550 8730
rect 463602 8678 463614 8730
rect 463666 8678 463672 8730
rect 463352 7744 463672 8678
rect 463352 7688 463364 7744
rect 463420 7688 463444 7744
rect 463500 7688 463524 7744
rect 463580 7688 463604 7744
rect 463660 7688 463672 7744
rect 463352 7664 463672 7688
rect 463352 7642 463364 7664
rect 463420 7642 463444 7664
rect 463500 7642 463524 7664
rect 463580 7642 463604 7664
rect 463660 7642 463672 7664
rect 463352 7590 463358 7642
rect 463420 7608 463422 7642
rect 463602 7608 463604 7642
rect 463410 7590 463422 7608
rect 463474 7590 463486 7608
rect 463538 7590 463550 7608
rect 463602 7590 463614 7608
rect 463666 7590 463672 7642
rect 463352 7584 463672 7590
rect 463352 7528 463364 7584
rect 463420 7528 463444 7584
rect 463500 7528 463524 7584
rect 463580 7528 463604 7584
rect 463660 7528 463672 7584
rect 463352 7504 463672 7528
rect 463352 7448 463364 7504
rect 463420 7448 463444 7504
rect 463500 7448 463524 7504
rect 463580 7448 463604 7504
rect 463660 7448 463672 7504
rect 463352 6554 463672 7448
rect 463352 6502 463358 6554
rect 463410 6502 463422 6554
rect 463474 6502 463486 6554
rect 463538 6502 463550 6554
rect 463602 6502 463614 6554
rect 463666 6502 463672 6554
rect 463352 5840 463672 6502
rect 464528 6316 464580 6322
rect 464528 6258 464580 6264
rect 463352 5784 463364 5840
rect 463420 5784 463444 5840
rect 463500 5784 463524 5840
rect 463580 5784 463604 5840
rect 463660 5784 463672 5840
rect 463352 5760 463672 5784
rect 463352 5704 463364 5760
rect 463420 5704 463444 5760
rect 463500 5704 463524 5760
rect 463580 5704 463604 5760
rect 463660 5704 463672 5760
rect 463352 5680 463672 5704
rect 463352 5624 463364 5680
rect 463420 5624 463444 5680
rect 463500 5624 463524 5680
rect 463580 5624 463604 5680
rect 463660 5624 463672 5680
rect 463352 5600 463672 5624
rect 463352 5544 463364 5600
rect 463420 5544 463444 5600
rect 463500 5544 463524 5600
rect 463580 5544 463604 5600
rect 463660 5544 463672 5600
rect 463352 5466 463672 5544
rect 463352 5414 463358 5466
rect 463410 5414 463422 5466
rect 463474 5414 463486 5466
rect 463538 5414 463550 5466
rect 463602 5414 463614 5466
rect 463666 5414 463672 5466
rect 463352 4378 463672 5414
rect 463352 4326 463358 4378
rect 463410 4326 463422 4378
rect 463474 4326 463486 4378
rect 463538 4326 463550 4378
rect 463602 4326 463614 4378
rect 463666 4326 463672 4378
rect 463352 3936 463672 4326
rect 463352 3880 463364 3936
rect 463420 3880 463444 3936
rect 463500 3880 463524 3936
rect 463580 3880 463604 3936
rect 463660 3880 463672 3936
rect 463352 3856 463672 3880
rect 463352 3800 463364 3856
rect 463420 3800 463444 3856
rect 463500 3800 463524 3856
rect 463580 3800 463604 3856
rect 463660 3800 463672 3856
rect 463352 3776 463672 3800
rect 463352 3720 463364 3776
rect 463420 3720 463444 3776
rect 463500 3720 463524 3776
rect 463580 3720 463604 3776
rect 463660 3720 463672 3776
rect 463352 3696 463672 3720
rect 463352 3640 463364 3696
rect 463420 3640 463444 3696
rect 463500 3640 463524 3696
rect 463580 3640 463604 3696
rect 463660 3640 463672 3696
rect 463352 3290 463672 3640
rect 463352 3238 463358 3290
rect 463410 3238 463422 3290
rect 463474 3238 463486 3290
rect 463538 3238 463550 3290
rect 463602 3238 463614 3290
rect 463666 3238 463672 3290
rect 463352 2202 463672 3238
rect 464540 2650 464568 6258
rect 477500 5364 477552 5370
rect 477500 5306 477552 5312
rect 475292 5160 475344 5166
rect 475292 5102 475344 5108
rect 464528 2644 464580 2650
rect 464528 2586 464580 2592
rect 466092 2576 466144 2582
rect 466368 2576 466420 2582
rect 466144 2524 466368 2530
rect 466092 2518 466420 2524
rect 466104 2502 466408 2518
rect 463700 2440 463752 2446
rect 463700 2382 463752 2388
rect 468852 2440 468904 2446
rect 468852 2382 468904 2388
rect 471428 2440 471480 2446
rect 471428 2382 471480 2388
rect 473912 2440 473964 2446
rect 473912 2382 473964 2388
rect 463712 2310 463740 2382
rect 468864 2310 468892 2382
rect 471440 2310 471468 2382
rect 473924 2310 473952 2382
rect 463700 2304 463752 2310
rect 463700 2246 463752 2252
rect 463792 2304 463844 2310
rect 463792 2246 463844 2252
rect 466460 2304 466512 2310
rect 466460 2246 466512 2252
rect 468852 2304 468904 2310
rect 468852 2246 468904 2252
rect 469220 2304 469272 2310
rect 469220 2246 469272 2252
rect 471428 2304 471480 2310
rect 471428 2246 471480 2252
rect 471888 2304 471940 2310
rect 471888 2246 471940 2252
rect 473912 2304 473964 2310
rect 473912 2246 473964 2252
rect 474004 2304 474056 2310
rect 474004 2246 474056 2252
rect 463352 2150 463358 2202
rect 463410 2150 463422 2202
rect 463474 2150 463486 2202
rect 463538 2150 463550 2202
rect 463602 2150 463614 2202
rect 463666 2150 463672 2202
rect 463352 304 463672 2150
rect 463712 2038 463740 2246
rect 463700 2032 463752 2038
rect 463700 1974 463752 1980
rect 463804 1222 463832 2246
rect 463792 1216 463844 1222
rect 463792 1158 463844 1164
rect 464252 1148 464304 1154
rect 464252 1090 464304 1096
rect 464264 814 464292 1090
rect 466472 1086 466500 2246
rect 468864 1834 468892 2246
rect 468852 1828 468904 1834
rect 468852 1770 468904 1776
rect 469232 1154 469260 2246
rect 471440 1970 471468 2246
rect 471428 1964 471480 1970
rect 471428 1906 471480 1912
rect 470600 1284 470652 1290
rect 470600 1226 470652 1232
rect 469220 1148 469272 1154
rect 469220 1090 469272 1096
rect 466460 1080 466512 1086
rect 466460 1022 466512 1028
rect 470612 882 470640 1226
rect 471900 1018 471928 2246
rect 473924 1630 473952 2246
rect 473912 1624 473964 1630
rect 473912 1566 473964 1572
rect 474016 1290 474044 2246
rect 475304 1766 475332 5102
rect 475384 2372 475436 2378
rect 475384 2314 475436 2320
rect 475396 2106 475424 2314
rect 475936 2304 475988 2310
rect 475936 2246 475988 2252
rect 475384 2100 475436 2106
rect 475384 2042 475436 2048
rect 475292 1760 475344 1766
rect 475292 1702 475344 1708
rect 474004 1284 474056 1290
rect 474004 1226 474056 1232
rect 472900 1216 472952 1222
rect 472900 1158 472952 1164
rect 471888 1012 471940 1018
rect 471888 954 471940 960
rect 470600 876 470652 882
rect 470600 818 470652 824
rect 472912 814 472940 1158
rect 475948 950 475976 2246
rect 477512 1698 477540 5306
rect 478892 5030 478920 10950
rect 480260 10940 480312 10946
rect 480260 10882 480312 10888
rect 480272 6254 480300 10882
rect 480260 6248 480312 6254
rect 480260 6190 480312 6196
rect 478880 5024 478932 5030
rect 478880 4966 478932 4972
rect 480364 3602 480392 10950
rect 480444 7948 480496 7954
rect 480444 7890 480496 7896
rect 480352 3596 480404 3602
rect 480352 3538 480404 3544
rect 480456 2774 480484 7890
rect 480732 5166 480760 11222
rect 481180 11144 481232 11150
rect 481180 11086 481232 11092
rect 480720 5160 480772 5166
rect 480720 5102 480772 5108
rect 480272 2746 480484 2774
rect 478512 2304 478564 2310
rect 478512 2246 478564 2252
rect 477500 1692 477552 1698
rect 477500 1634 477552 1640
rect 478524 1222 478552 2246
rect 480272 1834 480300 2746
rect 481192 1902 481220 11086
rect 481284 6186 481312 11222
rect 481640 10940 481692 10946
rect 481640 10882 481692 10888
rect 481272 6180 481324 6186
rect 481272 6122 481324 6128
rect 481652 5370 481680 10882
rect 481836 9674 481864 11290
rect 482100 11280 482152 11286
rect 482100 11222 482152 11228
rect 482284 11280 482336 11286
rect 482284 11222 482336 11228
rect 481836 9646 481956 9674
rect 481824 8288 481876 8294
rect 481824 8230 481876 8236
rect 481732 8084 481784 8090
rect 481732 8026 481784 8032
rect 481640 5364 481692 5370
rect 481640 5306 481692 5312
rect 481744 5250 481772 8026
rect 481652 5222 481772 5250
rect 481652 2514 481680 5222
rect 481732 5160 481784 5166
rect 481732 5102 481784 5108
rect 481744 2514 481772 5102
rect 481640 2508 481692 2514
rect 481640 2450 481692 2456
rect 481732 2508 481784 2514
rect 481732 2450 481784 2456
rect 481836 2038 481864 8230
rect 481928 4826 481956 9646
rect 482008 8016 482060 8022
rect 482008 7958 482060 7964
rect 482020 5166 482048 7958
rect 482112 6322 482140 11222
rect 482100 6316 482152 6322
rect 482100 6258 482152 6264
rect 482008 5160 482060 5166
rect 482008 5102 482060 5108
rect 481916 4820 481968 4826
rect 481916 4762 481968 4768
rect 482296 3466 482324 11222
rect 482848 9674 482876 11290
rect 483020 10940 483072 10946
rect 483020 10882 483072 10888
rect 482756 9646 482876 9674
rect 482284 3460 482336 3466
rect 482284 3402 482336 3408
rect 482756 2106 482784 9646
rect 483032 2582 483060 10882
rect 483124 8294 483152 11290
rect 483112 8288 483164 8294
rect 483112 8230 483164 8236
rect 483584 2650 483612 11342
rect 484492 11290 484544 11296
rect 486148 11348 486200 11354
rect 486148 11290 486200 11296
rect 486700 11348 486752 11354
rect 486700 11290 486752 11296
rect 486976 11348 487028 11354
rect 486976 11290 487028 11296
rect 488540 11348 488592 11354
rect 488540 11290 488592 11296
rect 488816 11348 488868 11354
rect 488816 11290 488868 11296
rect 530016 11300 530336 11312
rect 483664 11280 483716 11286
rect 483664 11222 483716 11228
rect 484216 11280 484268 11286
rect 484216 11222 484268 11228
rect 483676 7954 483704 11222
rect 484124 11008 484176 11014
rect 484124 10950 484176 10956
rect 483664 7948 483716 7954
rect 483664 7890 483716 7896
rect 483572 2644 483624 2650
rect 483572 2586 483624 2592
rect 483020 2576 483072 2582
rect 483020 2518 483072 2524
rect 483572 2304 483624 2310
rect 483572 2246 483624 2252
rect 482744 2100 482796 2106
rect 482744 2042 482796 2048
rect 481824 2032 481876 2038
rect 481824 1974 481876 1980
rect 481180 1896 481232 1902
rect 481180 1838 481232 1844
rect 480260 1828 480312 1834
rect 480260 1770 480312 1776
rect 481548 1352 481600 1358
rect 481548 1294 481600 1300
rect 478512 1216 478564 1222
rect 478512 1158 478564 1164
rect 478880 1148 478932 1154
rect 478880 1090 478932 1096
rect 475936 944 475988 950
rect 475936 886 475988 892
rect 478892 814 478920 1090
rect 481560 814 481588 1294
rect 483584 1018 483612 2246
rect 484136 1970 484164 10950
rect 484124 1964 484176 1970
rect 484124 1906 484176 1912
rect 484228 1630 484256 11222
rect 484308 10940 484360 10946
rect 484308 10882 484360 10888
rect 484320 2650 484348 10882
rect 484504 8090 484532 11290
rect 485780 11144 485832 11150
rect 485780 11086 485832 11092
rect 484952 11008 485004 11014
rect 484952 10950 485004 10956
rect 485044 11008 485096 11014
rect 485044 10950 485096 10956
rect 484492 8084 484544 8090
rect 484492 8026 484544 8032
rect 484308 2644 484360 2650
rect 484308 2586 484360 2592
rect 484320 2446 484348 2586
rect 484308 2440 484360 2446
rect 484308 2382 484360 2388
rect 484964 2378 484992 10950
rect 485056 8022 485084 10950
rect 485044 8016 485096 8022
rect 485044 7958 485096 7964
rect 485792 3194 485820 11086
rect 486160 8294 486188 11290
rect 486424 11280 486476 11286
rect 486424 11222 486476 11228
rect 486148 8288 486200 8294
rect 486148 8230 486200 8236
rect 486436 7546 486464 11222
rect 486424 7540 486476 7546
rect 486424 7482 486476 7488
rect 486712 7478 486740 11290
rect 486988 8022 487016 11290
rect 487252 11280 487304 11286
rect 487252 11222 487304 11228
rect 487528 11280 487580 11286
rect 487528 11222 487580 11228
rect 487804 11280 487856 11286
rect 487804 11222 487856 11228
rect 488080 11280 488132 11286
rect 488080 11222 488132 11228
rect 488356 11280 488408 11286
rect 488356 11222 488408 11228
rect 486976 8016 487028 8022
rect 486976 7958 487028 7964
rect 487264 7886 487292 11222
rect 487540 8090 487568 11222
rect 487528 8084 487580 8090
rect 487528 8026 487580 8032
rect 487816 7954 487844 11222
rect 487804 7948 487856 7954
rect 487804 7890 487856 7896
rect 487252 7880 487304 7886
rect 487252 7822 487304 7828
rect 488092 7818 488120 11222
rect 488080 7812 488132 7818
rect 488080 7754 488132 7760
rect 488368 7750 488396 11222
rect 488552 8378 488580 11290
rect 488460 8350 488580 8378
rect 488356 7744 488408 7750
rect 488356 7686 488408 7692
rect 486700 7472 486752 7478
rect 486700 7414 486752 7420
rect 488460 4826 488488 8350
rect 488540 8288 488592 8294
rect 488540 8230 488592 8236
rect 488448 4820 488500 4826
rect 488448 4762 488500 4768
rect 488552 3194 488580 8230
rect 485780 3188 485832 3194
rect 485780 3130 485832 3136
rect 488540 3188 488592 3194
rect 488540 3130 488592 3136
rect 485792 2446 485820 3130
rect 488552 2514 488580 3130
rect 488828 2774 488856 11290
rect 530016 11244 530028 11300
rect 530084 11244 530108 11300
rect 530164 11244 530188 11300
rect 530244 11244 530268 11300
rect 530324 11244 530336 11300
rect 530016 11220 530336 11244
rect 530016 11164 530028 11220
rect 530084 11164 530108 11220
rect 530164 11164 530188 11220
rect 530244 11164 530268 11220
rect 530324 11164 530336 11220
rect 530016 11140 530336 11164
rect 530016 11084 530028 11140
rect 530084 11084 530108 11140
rect 530164 11084 530188 11140
rect 530244 11084 530268 11140
rect 530324 11084 530336 11140
rect 530016 11060 530336 11084
rect 530016 11004 530028 11060
rect 530084 11004 530108 11060
rect 530164 11004 530188 11060
rect 530244 11004 530268 11060
rect 530324 11004 530336 11060
rect 530016 8988 530336 11004
rect 530016 8932 530028 8988
rect 530084 8932 530108 8988
rect 530164 8932 530188 8988
rect 530244 8932 530268 8988
rect 530324 8932 530336 8988
rect 530016 8908 530336 8932
rect 530016 8852 530028 8908
rect 530084 8852 530108 8908
rect 530164 8852 530188 8908
rect 530244 8852 530268 8908
rect 530324 8852 530336 8908
rect 530016 8828 530336 8852
rect 530016 8772 530028 8828
rect 530084 8772 530108 8828
rect 530164 8772 530188 8828
rect 530244 8772 530268 8828
rect 530324 8772 530336 8828
rect 530016 8748 530336 8772
rect 530016 8692 530028 8748
rect 530084 8692 530108 8748
rect 530164 8692 530188 8748
rect 530244 8692 530268 8748
rect 530324 8692 530336 8748
rect 501328 8084 501380 8090
rect 501328 8026 501380 8032
rect 496176 8016 496228 8022
rect 496176 7958 496228 7964
rect 491024 7540 491076 7546
rect 491024 7482 491076 7488
rect 491036 3194 491064 7482
rect 493600 7472 493652 7478
rect 493600 7414 493652 7420
rect 493612 3194 493640 7414
rect 496188 3194 496216 7958
rect 498752 7880 498804 7886
rect 498752 7822 498804 7828
rect 498764 3194 498792 7822
rect 501340 3194 501368 8026
rect 503904 7948 503956 7954
rect 503904 7890 503956 7896
rect 503916 3194 503944 7890
rect 506480 7812 506532 7818
rect 506480 7754 506532 7760
rect 506492 3194 506520 7754
rect 509056 7744 509108 7750
rect 509056 7686 509108 7692
rect 509068 3194 509096 7686
rect 530016 7084 530336 8692
rect 530016 7028 530028 7084
rect 530084 7028 530108 7084
rect 530164 7028 530188 7084
rect 530244 7028 530268 7084
rect 530324 7028 530336 7084
rect 530016 7004 530336 7028
rect 530016 6948 530028 7004
rect 530084 6948 530108 7004
rect 530164 6948 530188 7004
rect 530244 6948 530268 7004
rect 530324 6948 530336 7004
rect 530016 6924 530336 6948
rect 530016 6868 530028 6924
rect 530084 6868 530108 6924
rect 530164 6868 530188 6924
rect 530244 6868 530268 6924
rect 530324 6868 530336 6924
rect 530016 6844 530336 6868
rect 530016 6788 530028 6844
rect 530084 6788 530108 6844
rect 530164 6788 530188 6844
rect 530244 6788 530268 6844
rect 530324 6788 530336 6844
rect 530016 5180 530336 6788
rect 530016 5124 530028 5180
rect 530084 5124 530108 5180
rect 530164 5124 530188 5180
rect 530244 5124 530268 5180
rect 530324 5124 530336 5180
rect 530016 5100 530336 5124
rect 530016 5044 530028 5100
rect 530084 5044 530108 5100
rect 530164 5044 530188 5100
rect 530244 5044 530268 5100
rect 530324 5044 530336 5100
rect 530016 5020 530336 5044
rect 530016 4964 530028 5020
rect 530084 4964 530108 5020
rect 530164 4964 530188 5020
rect 530244 4964 530268 5020
rect 530324 4964 530336 5020
rect 530016 4940 530336 4964
rect 530016 4884 530028 4940
rect 530084 4884 530108 4940
rect 530164 4884 530188 4940
rect 530244 4884 530268 4940
rect 530324 4884 530336 4940
rect 511632 4820 511684 4826
rect 511632 4762 511684 4768
rect 511644 3194 511672 4762
rect 530016 3276 530336 4884
rect 530016 3220 530028 3276
rect 530084 3220 530108 3276
rect 530164 3220 530188 3276
rect 530244 3220 530268 3276
rect 530324 3220 530336 3276
rect 530016 3196 530336 3220
rect 491024 3188 491076 3194
rect 491024 3130 491076 3136
rect 493600 3188 493652 3194
rect 493600 3130 493652 3136
rect 496176 3188 496228 3194
rect 496176 3130 496228 3136
rect 498752 3188 498804 3194
rect 498752 3130 498804 3136
rect 501328 3188 501380 3194
rect 501328 3130 501380 3136
rect 503904 3188 503956 3194
rect 503904 3130 503956 3136
rect 506480 3188 506532 3194
rect 506480 3130 506532 3136
rect 509056 3188 509108 3194
rect 509056 3130 509108 3136
rect 511632 3188 511684 3194
rect 511632 3130 511684 3136
rect 530016 3140 530028 3196
rect 530084 3140 530108 3196
rect 530164 3140 530188 3196
rect 530244 3140 530268 3196
rect 530324 3140 530336 3196
rect 488736 2746 488856 2774
rect 488540 2508 488592 2514
rect 488540 2450 488592 2456
rect 488736 2446 488764 2746
rect 491036 2446 491064 3130
rect 493612 2446 493640 3130
rect 496188 2446 496216 3130
rect 498764 2446 498792 3130
rect 501340 2446 501368 3130
rect 503916 2446 503944 3130
rect 506492 2446 506520 3130
rect 509068 2446 509096 3130
rect 511644 2446 511672 3130
rect 530016 3116 530336 3140
rect 530016 3060 530028 3116
rect 530084 3060 530108 3116
rect 530164 3060 530188 3116
rect 530244 3060 530268 3116
rect 530324 3060 530336 3116
rect 530016 3036 530336 3060
rect 530016 2980 530028 3036
rect 530084 2980 530108 3036
rect 530164 2980 530188 3036
rect 530244 2980 530268 3036
rect 530324 2980 530336 3036
rect 514208 2848 514260 2854
rect 514208 2790 514260 2796
rect 514220 2446 514248 2790
rect 485780 2440 485832 2446
rect 485780 2382 485832 2388
rect 488724 2440 488776 2446
rect 488724 2382 488776 2388
rect 491024 2440 491076 2446
rect 491024 2382 491076 2388
rect 493600 2440 493652 2446
rect 493600 2382 493652 2388
rect 496176 2440 496228 2446
rect 496176 2382 496228 2388
rect 498752 2440 498804 2446
rect 498752 2382 498804 2388
rect 501328 2440 501380 2446
rect 501328 2382 501380 2388
rect 503904 2440 503956 2446
rect 503904 2382 503956 2388
rect 506480 2440 506532 2446
rect 506480 2382 506532 2388
rect 509056 2440 509108 2446
rect 509056 2382 509108 2388
rect 511632 2440 511684 2446
rect 511632 2382 511684 2388
rect 514208 2440 514260 2446
rect 514208 2382 514260 2388
rect 484952 2372 485004 2378
rect 484952 2314 485004 2320
rect 486148 2304 486200 2310
rect 486148 2246 486200 2252
rect 488724 2304 488776 2310
rect 488724 2246 488776 2252
rect 491300 2304 491352 2310
rect 491300 2246 491352 2252
rect 493876 2304 493928 2310
rect 493876 2246 493928 2252
rect 496452 2304 496504 2310
rect 496452 2246 496504 2252
rect 498200 2304 498252 2310
rect 498200 2246 498252 2252
rect 500316 2304 500368 2310
rect 500316 2246 500368 2252
rect 502340 2304 502392 2310
rect 502340 2246 502392 2252
rect 505100 2304 505152 2310
rect 505100 2246 505152 2252
rect 509332 2304 509384 2310
rect 509332 2246 509384 2252
rect 510528 2304 510580 2310
rect 510528 2246 510580 2252
rect 484216 1624 484268 1630
rect 484216 1566 484268 1572
rect 485964 1284 486016 1290
rect 485964 1226 486016 1232
rect 483756 1216 483808 1222
rect 483756 1158 483808 1164
rect 483572 1012 483624 1018
rect 483572 954 483624 960
rect 483768 814 483796 1158
rect 485976 814 486004 1226
rect 486160 882 486188 2246
rect 488736 1154 488764 2246
rect 491312 1358 491340 2246
rect 491300 1352 491352 1358
rect 491300 1294 491352 1300
rect 493888 1222 493916 2246
rect 496464 1290 496492 2246
rect 496452 1284 496504 1290
rect 496452 1226 496504 1232
rect 493876 1216 493928 1222
rect 493876 1158 493928 1164
rect 488724 1148 488776 1154
rect 488724 1090 488776 1096
rect 491116 1148 491168 1154
rect 491116 1090 491168 1096
rect 486148 876 486200 882
rect 486148 818 486200 824
rect 464252 808 464304 814
rect 464252 750 464304 756
rect 472900 808 472952 814
rect 472900 750 472952 756
rect 478880 808 478932 814
rect 478880 750 478932 756
rect 481548 808 481600 814
rect 481548 750 481600 756
rect 483756 808 483808 814
rect 483756 750 483808 756
rect 485964 808 486016 814
rect 485964 750 486016 756
rect 491128 746 491156 1090
rect 498212 1086 498240 2246
rect 499212 1284 499264 1290
rect 499212 1226 499264 1232
rect 498292 1216 498344 1222
rect 498292 1158 498344 1164
rect 498200 1080 498252 1086
rect 498200 1022 498252 1028
rect 498304 814 498332 1158
rect 499120 1148 499172 1154
rect 499120 1090 499172 1096
rect 499132 950 499160 1090
rect 499224 1086 499252 1226
rect 499212 1080 499264 1086
rect 499212 1022 499264 1028
rect 500328 1018 500356 2246
rect 502352 1086 502380 2246
rect 505112 1154 505140 2246
rect 505100 1148 505152 1154
rect 505100 1090 505152 1096
rect 502340 1080 502392 1086
rect 502340 1022 502392 1028
rect 500316 1012 500368 1018
rect 500316 954 500368 960
rect 499120 944 499172 950
rect 499120 886 499172 892
rect 509344 882 509372 2246
rect 510540 1222 510568 2246
rect 510528 1216 510580 1222
rect 510528 1158 510580 1164
rect 509332 876 509384 882
rect 509332 818 509384 824
rect 498292 808 498344 814
rect 498292 750 498344 756
rect 491116 740 491168 746
rect 491116 682 491168 688
rect 463352 248 463364 304
rect 463420 248 463444 304
rect 463500 248 463524 304
rect 463580 248 463604 304
rect 463660 248 463672 304
rect 463352 224 463672 248
rect 463352 168 463364 224
rect 463420 168 463444 224
rect 463500 168 463524 224
rect 463580 168 463604 224
rect 463660 168 463672 224
rect 463352 144 463672 168
rect 463352 88 463364 144
rect 463420 88 463444 144
rect 463500 88 463524 144
rect 463580 88 463604 144
rect 463660 88 463672 144
rect 463352 64 463672 88
rect 514220 66 514248 2382
rect 530016 964 530336 2980
rect 530016 908 530028 964
rect 530084 908 530108 964
rect 530164 908 530188 964
rect 530244 908 530268 964
rect 530324 908 530336 964
rect 530016 884 530336 908
rect 530016 828 530028 884
rect 530084 828 530108 884
rect 530164 828 530188 884
rect 530244 828 530268 884
rect 530324 828 530336 884
rect 530016 804 530336 828
rect 530016 748 530028 804
rect 530084 748 530108 804
rect 530164 748 530188 804
rect 530244 748 530268 804
rect 530324 748 530336 804
rect 530016 724 530336 748
rect 530016 668 530028 724
rect 530084 668 530108 724
rect 530164 668 530188 724
rect 530244 668 530268 724
rect 530324 668 530336 724
rect 530016 656 530336 668
rect 530676 9648 530996 11664
rect 530676 9592 530688 9648
rect 530744 9592 530768 9648
rect 530824 9592 530848 9648
rect 530904 9592 530928 9648
rect 530984 9592 530996 9648
rect 530676 9568 530996 9592
rect 530676 9512 530688 9568
rect 530744 9512 530768 9568
rect 530824 9512 530848 9568
rect 530904 9512 530928 9568
rect 530984 9512 530996 9568
rect 530676 9488 530996 9512
rect 530676 9432 530688 9488
rect 530744 9432 530768 9488
rect 530824 9432 530848 9488
rect 530904 9432 530928 9488
rect 530984 9432 530996 9488
rect 530676 9408 530996 9432
rect 530676 9352 530688 9408
rect 530744 9352 530768 9408
rect 530824 9352 530848 9408
rect 530904 9352 530928 9408
rect 530984 9352 530996 9408
rect 530676 7744 530996 9352
rect 530676 7688 530688 7744
rect 530744 7688 530768 7744
rect 530824 7688 530848 7744
rect 530904 7688 530928 7744
rect 530984 7688 530996 7744
rect 530676 7664 530996 7688
rect 530676 7608 530688 7664
rect 530744 7608 530768 7664
rect 530824 7608 530848 7664
rect 530904 7608 530928 7664
rect 530984 7608 530996 7664
rect 530676 7584 530996 7608
rect 530676 7528 530688 7584
rect 530744 7528 530768 7584
rect 530824 7528 530848 7584
rect 530904 7528 530928 7584
rect 530984 7528 530996 7584
rect 530676 7504 530996 7528
rect 530676 7448 530688 7504
rect 530744 7448 530768 7504
rect 530824 7448 530848 7504
rect 530904 7448 530928 7504
rect 530984 7448 530996 7504
rect 530676 5840 530996 7448
rect 530676 5784 530688 5840
rect 530744 5784 530768 5840
rect 530824 5784 530848 5840
rect 530904 5784 530928 5840
rect 530984 5784 530996 5840
rect 530676 5760 530996 5784
rect 530676 5704 530688 5760
rect 530744 5704 530768 5760
rect 530824 5704 530848 5760
rect 530904 5704 530928 5760
rect 530984 5704 530996 5760
rect 530676 5680 530996 5704
rect 530676 5624 530688 5680
rect 530744 5624 530768 5680
rect 530824 5624 530848 5680
rect 530904 5624 530928 5680
rect 530984 5624 530996 5680
rect 530676 5600 530996 5624
rect 530676 5544 530688 5600
rect 530744 5544 530768 5600
rect 530824 5544 530848 5600
rect 530904 5544 530928 5600
rect 530984 5544 530996 5600
rect 530676 3936 530996 5544
rect 530676 3880 530688 3936
rect 530744 3880 530768 3936
rect 530824 3880 530848 3936
rect 530904 3880 530928 3936
rect 530984 3880 530996 3936
rect 530676 3856 530996 3880
rect 530676 3800 530688 3856
rect 530744 3800 530768 3856
rect 530824 3800 530848 3856
rect 530904 3800 530928 3856
rect 530984 3800 530996 3856
rect 530676 3776 530996 3800
rect 530676 3720 530688 3776
rect 530744 3720 530768 3776
rect 530824 3720 530848 3776
rect 530904 3720 530928 3776
rect 530984 3720 530996 3776
rect 530676 3696 530996 3720
rect 530676 3640 530688 3696
rect 530744 3640 530768 3696
rect 530824 3640 530848 3696
rect 530904 3640 530928 3696
rect 530984 3640 530996 3696
rect 530676 304 530996 3640
rect 530676 248 530688 304
rect 530744 248 530768 304
rect 530824 248 530848 304
rect 530904 248 530928 304
rect 530984 248 530996 304
rect 530676 224 530996 248
rect 530676 168 530688 224
rect 530744 168 530768 224
rect 530824 168 530848 224
rect 530904 168 530928 224
rect 530984 168 530996 224
rect 530676 144 530996 168
rect 530676 88 530688 144
rect 530744 88 530768 144
rect 530824 88 530848 144
rect 530904 88 530928 144
rect 530984 88 530996 144
rect 463352 8 463364 64
rect 463420 8 463444 64
rect 463500 8 463524 64
rect 463580 8 463604 64
rect 463660 8 463672 64
rect 463352 -4 463672 8
rect 514208 60 514260 66
rect 514208 2 514260 8
rect 530676 64 530996 88
rect 530676 8 530688 64
rect 530744 8 530768 64
rect 530824 8 530848 64
rect 530904 8 530928 64
rect 530984 8 530996 64
rect 530676 -4 530996 8
<< via2 >>
rect -1064 11904 -1008 11960
rect -984 11904 -928 11960
rect -904 11904 -848 11960
rect -824 11904 -768 11960
rect -1064 11824 -1008 11880
rect -984 11824 -928 11880
rect -904 11824 -848 11880
rect -824 11824 -768 11880
rect -1064 11744 -1008 11800
rect -984 11744 -928 11800
rect -904 11744 -848 11800
rect -824 11744 -768 11800
rect -1064 11664 -1008 11720
rect -984 11664 -928 11720
rect -904 11664 -848 11720
rect -824 11664 -768 11720
rect -1064 9592 -1008 9648
rect -984 9592 -928 9648
rect -904 9592 -848 9648
rect -824 9592 -768 9648
rect -1064 9512 -1008 9568
rect -984 9512 -928 9568
rect -904 9512 -848 9568
rect -824 9512 -768 9568
rect -1064 9432 -1008 9488
rect -984 9432 -928 9488
rect -904 9432 -848 9488
rect -824 9432 -768 9488
rect -1064 9352 -1008 9408
rect -984 9352 -928 9408
rect -904 9352 -848 9408
rect -824 9352 -768 9408
rect -1064 7688 -1008 7744
rect -984 7688 -928 7744
rect -904 7688 -848 7744
rect -824 7688 -768 7744
rect -1064 7608 -1008 7664
rect -984 7608 -928 7664
rect -904 7608 -848 7664
rect -824 7608 -768 7664
rect -1064 7528 -1008 7584
rect -984 7528 -928 7584
rect -904 7528 -848 7584
rect -824 7528 -768 7584
rect -1064 7448 -1008 7504
rect -984 7448 -928 7504
rect -904 7448 -848 7504
rect -824 7448 -768 7504
rect -1064 5784 -1008 5840
rect -984 5784 -928 5840
rect -904 5784 -848 5840
rect -824 5784 -768 5840
rect -1064 5704 -1008 5760
rect -984 5704 -928 5760
rect -904 5704 -848 5760
rect -824 5704 -768 5760
rect -1064 5624 -1008 5680
rect -984 5624 -928 5680
rect -904 5624 -848 5680
rect -824 5624 -768 5680
rect -1064 5544 -1008 5600
rect -984 5544 -928 5600
rect -904 5544 -848 5600
rect -824 5544 -768 5600
rect -1064 3880 -1008 3936
rect -984 3880 -928 3936
rect -904 3880 -848 3936
rect -824 3880 -768 3936
rect -1064 3800 -1008 3856
rect -984 3800 -928 3856
rect -904 3800 -848 3856
rect -824 3800 -768 3856
rect -1064 3720 -1008 3776
rect -984 3720 -928 3776
rect -904 3720 -848 3776
rect -824 3720 -768 3776
rect -1064 3640 -1008 3696
rect -984 3640 -928 3696
rect -904 3640 -848 3696
rect -824 3640 -768 3696
rect -404 11244 -348 11300
rect -324 11244 -268 11300
rect -244 11244 -188 11300
rect -164 11244 -108 11300
rect -404 11164 -348 11220
rect -324 11164 -268 11220
rect -244 11164 -188 11220
rect -164 11164 -108 11220
rect -404 11084 -348 11140
rect -324 11084 -268 11140
rect -244 11084 -188 11140
rect -164 11084 -108 11140
rect -404 11004 -348 11060
rect -324 11004 -268 11060
rect -244 11004 -188 11060
rect -164 11004 -108 11060
rect 66920 11244 66976 11300
rect 67000 11244 67056 11300
rect 67080 11244 67136 11300
rect 67160 11244 67216 11300
rect 66920 11164 66976 11220
rect 67000 11164 67056 11220
rect 67080 11164 67136 11220
rect 67160 11164 67216 11220
rect 66920 11084 66976 11140
rect 67000 11084 67056 11140
rect 67080 11084 67136 11140
rect 67160 11084 67216 11140
rect 66920 11004 66976 11060
rect 67000 11004 67056 11060
rect 67080 11004 67136 11060
rect 67160 11004 67216 11060
rect -404 8932 -348 8988
rect -324 8932 -268 8988
rect -244 8932 -188 8988
rect -164 8932 -108 8988
rect -404 8852 -348 8908
rect -324 8852 -268 8908
rect -244 8852 -188 8908
rect -164 8852 -108 8908
rect -404 8772 -348 8828
rect -324 8772 -268 8828
rect -244 8772 -188 8828
rect -164 8772 -108 8828
rect -404 8692 -348 8748
rect -324 8692 -268 8748
rect -244 8692 -188 8748
rect -164 8692 -108 8748
rect -404 7028 -348 7084
rect -324 7028 -268 7084
rect -244 7028 -188 7084
rect -164 7028 -108 7084
rect -404 6948 -348 7004
rect -324 6948 -268 7004
rect -244 6948 -188 7004
rect -164 6948 -108 7004
rect -404 6868 -348 6924
rect -324 6868 -268 6924
rect -244 6868 -188 6924
rect -164 6868 -108 6924
rect -404 6788 -348 6844
rect -324 6788 -268 6844
rect -244 6788 -188 6844
rect -164 6788 -108 6844
rect -404 5124 -348 5180
rect -324 5124 -268 5180
rect -244 5124 -188 5180
rect -164 5124 -108 5180
rect -404 5044 -348 5100
rect -324 5044 -268 5100
rect -244 5044 -188 5100
rect -164 5044 -108 5100
rect -404 4964 -348 5020
rect -324 4964 -268 5020
rect -244 4964 -188 5020
rect -164 4964 -108 5020
rect -404 4884 -348 4940
rect -324 4884 -268 4940
rect -244 4884 -188 4940
rect -164 4884 -108 4940
rect -404 3220 -348 3276
rect -324 3220 -268 3276
rect -244 3220 -188 3276
rect -164 3220 -108 3276
rect -404 3140 -348 3196
rect -324 3140 -268 3196
rect -244 3140 -188 3196
rect -164 3140 -108 3196
rect -404 3060 -348 3116
rect -324 3060 -268 3116
rect -244 3060 -188 3116
rect -164 3060 -108 3116
rect -404 2980 -348 3036
rect -324 2980 -268 3036
rect -244 2980 -188 3036
rect -164 2980 -108 3036
rect -404 908 -348 964
rect -324 908 -268 964
rect -244 908 -188 964
rect -164 908 -108 964
rect -404 828 -348 884
rect -324 828 -268 884
rect -244 828 -188 884
rect -164 828 -108 884
rect -404 748 -348 804
rect -324 748 -268 804
rect -244 748 -188 804
rect -164 748 -108 804
rect 28354 2372 28410 2408
rect 28354 2352 28356 2372
rect 28356 2352 28408 2372
rect 28408 2352 28410 2372
rect 32770 3440 32826 3496
rect 41234 2508 41290 2544
rect 41234 2488 41236 2508
rect 41236 2488 41288 2508
rect 41288 2488 41290 2508
rect 48962 2624 49018 2680
rect 55954 2760 56010 2816
rect 66920 8932 66976 8988
rect 67000 8932 67056 8988
rect 67080 8932 67136 8988
rect 67160 8932 67216 8988
rect 66920 8852 66976 8908
rect 67000 8852 67056 8908
rect 67080 8852 67136 8908
rect 67160 8852 67216 8908
rect 66920 8772 66976 8828
rect 67000 8772 67056 8828
rect 67080 8772 67136 8828
rect 67160 8772 67216 8828
rect 66920 8692 66976 8748
rect 67000 8692 67056 8748
rect 67080 8692 67136 8748
rect 67160 8692 67216 8748
rect 67580 11904 67636 11960
rect 67660 11904 67716 11960
rect 67740 11904 67796 11960
rect 67820 11904 67876 11960
rect 67580 11824 67636 11880
rect 67660 11824 67716 11880
rect 67740 11824 67796 11880
rect 67820 11824 67876 11880
rect 67580 11744 67636 11800
rect 67660 11744 67716 11800
rect 67740 11744 67796 11800
rect 67820 11744 67876 11800
rect 67580 11664 67636 11720
rect 67660 11664 67716 11720
rect 67740 11664 67796 11720
rect 67820 11664 67876 11720
rect 67580 9592 67636 9648
rect 67660 9592 67716 9648
rect 67740 9592 67796 9648
rect 67820 9592 67876 9648
rect 67580 9512 67636 9568
rect 67660 9512 67716 9568
rect 67740 9512 67796 9568
rect 67820 9512 67876 9568
rect 67580 9432 67636 9488
rect 67660 9432 67716 9488
rect 67740 9432 67796 9488
rect 67820 9432 67876 9488
rect 67580 9352 67636 9408
rect 67660 9352 67716 9408
rect 67740 9352 67796 9408
rect 67820 9352 67876 9408
rect 67270 8472 67326 8528
rect 66920 7046 66966 7084
rect 66966 7046 66976 7084
rect 67000 7046 67030 7084
rect 67030 7046 67042 7084
rect 67042 7046 67056 7084
rect 67080 7046 67094 7084
rect 67094 7046 67106 7084
rect 67106 7046 67136 7084
rect 67160 7046 67170 7084
rect 67170 7046 67216 7084
rect 66920 7028 66976 7046
rect 67000 7028 67056 7046
rect 67080 7028 67136 7046
rect 67160 7028 67216 7046
rect 66920 6948 66976 7004
rect 67000 6948 67056 7004
rect 67080 6948 67136 7004
rect 67160 6948 67216 7004
rect 66920 6868 66976 6924
rect 67000 6868 67056 6924
rect 67080 6868 67136 6924
rect 67160 6868 67216 6924
rect 66920 6788 66976 6844
rect 67000 6788 67056 6844
rect 67080 6788 67136 6844
rect 67160 6788 67216 6844
rect 66920 5124 66976 5180
rect 67000 5124 67056 5180
rect 67080 5124 67136 5180
rect 67160 5124 67216 5180
rect 66920 5044 66976 5100
rect 67000 5044 67056 5100
rect 67080 5044 67136 5100
rect 67160 5044 67216 5100
rect 66920 4964 66976 5020
rect 67000 4964 67056 5020
rect 67080 4964 67136 5020
rect 67160 4964 67216 5020
rect 66920 4922 66976 4940
rect 67000 4922 67056 4940
rect 67080 4922 67136 4940
rect 67160 4922 67216 4940
rect 66920 4884 66966 4922
rect 66966 4884 66976 4922
rect 67000 4884 67030 4922
rect 67030 4884 67042 4922
rect 67042 4884 67056 4922
rect 67080 4884 67094 4922
rect 67094 4884 67106 4922
rect 67106 4884 67136 4922
rect 67160 4884 67170 4922
rect 67170 4884 67216 4922
rect 64418 2080 64474 2136
rect 67580 7688 67636 7744
rect 67660 7688 67716 7744
rect 67740 7688 67796 7744
rect 67820 7688 67876 7744
rect 67580 7642 67636 7664
rect 67660 7642 67716 7664
rect 67740 7642 67796 7664
rect 67820 7642 67876 7664
rect 67580 7608 67626 7642
rect 67626 7608 67636 7642
rect 67660 7608 67690 7642
rect 67690 7608 67702 7642
rect 67702 7608 67716 7642
rect 67740 7608 67754 7642
rect 67754 7608 67766 7642
rect 67766 7608 67796 7642
rect 67820 7608 67830 7642
rect 67830 7608 67876 7642
rect 67580 7528 67636 7584
rect 67660 7528 67716 7584
rect 67740 7528 67796 7584
rect 67820 7528 67876 7584
rect 67580 7448 67636 7504
rect 67660 7448 67716 7504
rect 67740 7448 67796 7504
rect 67820 7448 67876 7504
rect 67580 5784 67636 5840
rect 67660 5784 67716 5840
rect 67740 5784 67796 5840
rect 67820 5784 67876 5840
rect 67580 5704 67636 5760
rect 67660 5704 67716 5760
rect 67740 5704 67796 5760
rect 67820 5704 67876 5760
rect 67580 5624 67636 5680
rect 67660 5624 67716 5680
rect 67740 5624 67796 5680
rect 67820 5624 67876 5680
rect 67580 5544 67636 5600
rect 67660 5544 67716 5600
rect 67740 5544 67796 5600
rect 67820 5544 67876 5600
rect 67580 3880 67636 3936
rect 67660 3880 67716 3936
rect 67740 3880 67796 3936
rect 67820 3880 67876 3936
rect 67580 3800 67636 3856
rect 67660 3800 67716 3856
rect 67740 3800 67796 3856
rect 67820 3800 67876 3856
rect 67580 3720 67636 3776
rect 67660 3720 67716 3776
rect 67740 3720 67796 3776
rect 67820 3720 67876 3776
rect 67580 3640 67636 3696
rect 67660 3640 67716 3696
rect 67740 3640 67796 3696
rect 67820 3640 67876 3696
rect 66920 3220 66976 3276
rect 67000 3220 67056 3276
rect 67080 3220 67136 3276
rect 67160 3220 67216 3276
rect 66920 3140 66976 3196
rect 67000 3140 67056 3196
rect 67080 3140 67136 3196
rect 67160 3140 67216 3196
rect 66920 3060 66976 3116
rect 67000 3060 67056 3116
rect 67080 3060 67136 3116
rect 67160 3060 67216 3116
rect 66920 2980 66976 3036
rect 67000 2980 67056 3036
rect 67080 2980 67136 3036
rect 67160 2980 67216 3036
rect 66920 908 66976 964
rect 67000 908 67056 964
rect 67080 908 67136 964
rect 67160 908 67216 964
rect 66920 828 66976 884
rect 67000 828 67056 884
rect 67080 828 67136 884
rect 67160 828 67216 884
rect -404 668 -348 724
rect -324 668 -268 724
rect -244 668 -188 724
rect -164 668 -108 724
rect 66920 748 66976 804
rect 67000 748 67056 804
rect 67080 748 67136 804
rect 67160 748 67216 804
rect 66920 668 66976 724
rect 67000 668 67056 724
rect 67080 668 67136 724
rect 67160 668 67216 724
rect -1064 248 -1008 304
rect -984 248 -928 304
rect -904 248 -848 304
rect -824 248 -768 304
rect -1064 168 -1008 224
rect -984 168 -928 224
rect -904 168 -848 224
rect -824 168 -768 224
rect -1064 88 -1008 144
rect -984 88 -928 144
rect -904 88 -848 144
rect -824 88 -768 144
rect -1064 8 -1008 64
rect -984 8 -928 64
rect -904 8 -848 64
rect -824 8 -768 64
rect 68098 1128 68154 1184
rect 69846 1128 69902 1184
rect 72146 1672 72202 1728
rect 81714 4664 81770 4720
rect 67580 248 67636 304
rect 67660 248 67716 304
rect 67740 248 67796 304
rect 67820 248 67876 304
rect 67580 168 67636 224
rect 67660 168 67716 224
rect 67740 168 67796 224
rect 67820 168 67876 224
rect 67580 88 67636 144
rect 67660 88 67716 144
rect 67740 88 67796 144
rect 67820 88 67876 144
rect 79874 1536 79930 1592
rect 81346 1148 81402 1184
rect 81346 1128 81348 1148
rect 81348 1128 81400 1148
rect 81400 1128 81402 1148
rect 84014 1128 84070 1184
rect 86866 1264 86922 1320
rect 87326 1400 87382 1456
rect 93490 7928 93546 7984
rect 92386 4528 92442 4584
rect 90178 1128 90234 1184
rect 95330 1808 95386 1864
rect 96618 1400 96674 1456
rect 94778 1264 94834 1320
rect 101862 8064 101918 8120
rect 96710 1128 96766 1184
rect 97538 1264 97594 1320
rect 99010 2216 99066 2272
rect 98826 1400 98882 1456
rect 97906 1128 97962 1184
rect 99378 1944 99434 2000
rect 103058 9152 103114 9208
rect 101126 1400 101182 1456
rect 100758 1264 100814 1320
rect 100942 1264 100998 1320
rect 104438 3440 104494 3496
rect 105082 3476 105084 3496
rect 105084 3476 105136 3496
rect 105136 3476 105138 3496
rect 105082 3440 105138 3476
rect 105634 3460 105690 3496
rect 105634 3440 105636 3460
rect 105636 3440 105688 3460
rect 105688 3440 105690 3460
rect 108302 1400 108358 1456
rect 108854 1264 108910 1320
rect 111890 2216 111946 2272
rect 114190 6568 114246 6624
rect 112994 2796 112996 2816
rect 112996 2796 113048 2816
rect 113048 2796 113050 2816
rect 112994 2760 113050 2796
rect 113178 2760 113234 2816
rect 112350 1944 112406 2000
rect 114558 1400 114614 1456
rect 111890 1128 111946 1184
rect 114742 1264 114798 1320
rect 89166 484 89168 504
rect 89168 484 89220 504
rect 89220 484 89222 504
rect 89166 448 89222 484
rect 94686 448 94742 504
rect 97906 468 97962 504
rect 97906 448 97908 468
rect 97908 448 97960 468
rect 97960 448 97962 468
rect 103610 448 103666 504
rect 108854 448 108910 504
rect 109130 448 109186 504
rect 110694 448 110750 504
rect 115110 1164 115112 1184
rect 115112 1164 115164 1184
rect 115164 1164 115166 1184
rect 115110 1128 115166 1164
rect 114742 468 114798 504
rect 114742 448 114744 468
rect 114744 448 114796 468
rect 114796 448 114798 468
rect 116030 448 116086 504
rect 118606 1944 118662 2000
rect 117962 1264 118018 1320
rect 118514 1128 118570 1184
rect 119342 2760 119398 2816
rect 118790 1128 118846 1184
rect 119526 1400 119582 1456
rect 125506 6316 125562 6352
rect 125506 6296 125508 6316
rect 125508 6296 125560 6316
rect 125560 6296 125562 6316
rect 125690 4664 125746 4720
rect 130934 6160 130990 6216
rect 121090 2760 121146 2816
rect 120170 1128 120226 1184
rect 124494 1944 124550 2000
rect 126242 1944 126298 2000
rect 131210 4548 131266 4584
rect 131210 4528 131212 4548
rect 131212 4528 131264 4548
rect 131264 4528 131266 4548
rect 127070 1400 127126 1456
rect 135534 6024 135590 6080
rect 133510 4664 133566 4720
rect 130474 1400 130530 1456
rect 137834 4392 137890 4448
rect 141330 5344 141386 5400
rect 136638 2352 136694 2408
rect 135258 1400 135314 1456
rect 145930 4528 145986 4584
rect 144826 4256 144882 4312
rect 146850 2372 146906 2408
rect 146850 2352 146852 2372
rect 146852 2352 146904 2372
rect 146904 2352 146906 2372
rect 146390 1400 146446 1456
rect 149058 2488 149114 2544
rect 156694 2624 156750 2680
rect 67580 8 67636 64
rect 67660 8 67716 64
rect 67740 8 67796 64
rect 67820 8 67876 64
rect 150530 1400 150586 1456
rect 154670 1400 154726 1456
rect 156970 1400 157026 1456
rect 157154 1400 157210 1456
rect 158902 2488 158958 2544
rect 158718 1672 158774 1728
rect 164146 2624 164202 2680
rect 168194 1672 168250 1728
rect 169298 2252 169300 2272
rect 169300 2252 169352 2272
rect 169352 2252 169354 2272
rect 169298 2216 169354 2252
rect 168378 1400 168434 1456
rect 168562 1400 168618 1456
rect 175278 8472 175334 8528
rect 172518 8336 172574 8392
rect 176658 8200 176714 8256
rect 184202 8472 184258 8528
rect 182914 7248 182970 7304
rect 171230 2080 171286 2136
rect 173070 1400 173126 1456
rect 174450 2080 174506 2136
rect 178038 1672 178094 1728
rect 178682 1672 178738 1728
rect 176382 1400 176438 1456
rect 183558 1400 183614 1456
rect 183926 1400 183982 1456
rect 186134 1536 186190 1592
rect 199508 11904 199564 11960
rect 199588 11904 199644 11960
rect 199668 11904 199724 11960
rect 199748 11904 199804 11960
rect 198848 11244 198904 11300
rect 198928 11244 198984 11300
rect 199008 11244 199064 11300
rect 199088 11244 199144 11300
rect 198848 11164 198904 11220
rect 198928 11164 198984 11220
rect 199008 11164 199064 11220
rect 199088 11164 199144 11220
rect 198370 9988 198426 10024
rect 198370 9968 198372 9988
rect 198372 9968 198424 9988
rect 198424 9968 198426 9988
rect 197818 9832 197874 9888
rect 187330 1672 187386 1728
rect 190458 1808 190514 1864
rect 191102 1808 191158 1864
rect 189078 1536 189134 1592
rect 191746 1400 191802 1456
rect 195150 1536 195206 1592
rect 195978 3440 196034 3496
rect 196162 3440 196218 3496
rect 195150 1400 195206 1456
rect 198646 10784 198702 10840
rect 198848 11084 198904 11140
rect 198928 11084 198984 11140
rect 199008 11084 199064 11140
rect 199088 11084 199144 11140
rect 199508 11824 199564 11880
rect 199588 11824 199644 11880
rect 199668 11824 199724 11880
rect 199748 11824 199804 11880
rect 199508 11744 199564 11800
rect 199588 11744 199644 11800
rect 199668 11744 199724 11800
rect 199748 11744 199804 11800
rect 199508 11664 199564 11720
rect 199588 11664 199644 11720
rect 199668 11664 199724 11720
rect 199748 11664 199804 11720
rect 199382 11464 199438 11520
rect 198848 11004 198904 11060
rect 198928 11004 198984 11060
rect 199008 11004 199064 11060
rect 199088 11004 199144 11060
rect 198646 10104 198702 10160
rect 199290 10648 199346 10704
rect 199290 10512 199346 10568
rect 202050 11464 202106 11520
rect 200946 10784 201002 10840
rect 201498 10376 201554 10432
rect 199508 9592 199564 9648
rect 199588 9592 199644 9648
rect 199668 9592 199724 9648
rect 199748 9592 199804 9648
rect 199508 9512 199564 9568
rect 199588 9512 199644 9568
rect 199668 9512 199724 9568
rect 199748 9512 199804 9568
rect 199508 9432 199564 9488
rect 199588 9432 199644 9488
rect 199668 9432 199724 9488
rect 199748 9432 199804 9488
rect 199508 9352 199564 9408
rect 199588 9352 199644 9408
rect 199668 9352 199724 9408
rect 199748 9352 199804 9408
rect 198848 8932 198904 8988
rect 198928 8932 198984 8988
rect 199008 8932 199064 8988
rect 199088 8932 199144 8988
rect 198848 8852 198904 8908
rect 198928 8852 198984 8908
rect 199008 8852 199064 8908
rect 199088 8852 199144 8908
rect 198848 8772 198904 8828
rect 198928 8772 198984 8828
rect 199008 8772 199064 8828
rect 199088 8772 199144 8828
rect 198848 8692 198904 8748
rect 198928 8692 198984 8748
rect 199008 8692 199064 8748
rect 199088 8692 199144 8748
rect 198848 7046 198894 7084
rect 198894 7046 198904 7084
rect 198928 7046 198958 7084
rect 198958 7046 198970 7084
rect 198970 7046 198984 7084
rect 199008 7046 199022 7084
rect 199022 7046 199034 7084
rect 199034 7046 199064 7084
rect 199088 7046 199098 7084
rect 199098 7046 199144 7084
rect 198848 7028 198904 7046
rect 198928 7028 198984 7046
rect 199008 7028 199064 7046
rect 199088 7028 199144 7046
rect 198848 6948 198904 7004
rect 198928 6948 198984 7004
rect 199008 6948 199064 7004
rect 199088 6948 199144 7004
rect 198848 6868 198904 6924
rect 198928 6868 198984 6924
rect 199008 6868 199064 6924
rect 199088 6868 199144 6924
rect 198848 6788 198904 6844
rect 198928 6788 198984 6844
rect 199008 6788 199064 6844
rect 199088 6788 199144 6844
rect 198848 5124 198904 5180
rect 198928 5124 198984 5180
rect 199008 5124 199064 5180
rect 199088 5124 199144 5180
rect 198848 5044 198904 5100
rect 198928 5044 198984 5100
rect 199008 5044 199064 5100
rect 199088 5044 199144 5100
rect 198848 4964 198904 5020
rect 198928 4964 198984 5020
rect 199008 4964 199064 5020
rect 199088 4964 199144 5020
rect 198848 4922 198904 4940
rect 198928 4922 198984 4940
rect 199008 4922 199064 4940
rect 199088 4922 199144 4940
rect 198848 4884 198894 4922
rect 198894 4884 198904 4922
rect 198928 4884 198958 4922
rect 198958 4884 198970 4922
rect 198970 4884 198984 4922
rect 199008 4884 199022 4922
rect 199022 4884 199034 4922
rect 199034 4884 199064 4922
rect 199088 4884 199098 4922
rect 199098 4884 199144 4922
rect 198848 3220 198904 3276
rect 198928 3220 198984 3276
rect 199008 3220 199064 3276
rect 199088 3220 199144 3276
rect 198848 3140 198904 3196
rect 198928 3140 198984 3196
rect 199008 3140 199064 3196
rect 199088 3140 199144 3196
rect 198848 3060 198904 3116
rect 198928 3060 198984 3116
rect 199008 3060 199064 3116
rect 199088 3060 199144 3116
rect 198848 2980 198904 3036
rect 198928 2980 198984 3036
rect 199008 2980 199064 3036
rect 199088 2980 199144 3036
rect 198848 908 198904 964
rect 198928 908 198984 964
rect 199008 908 199064 964
rect 199088 908 199144 964
rect 198848 828 198904 884
rect 198928 828 198984 884
rect 199008 828 199064 884
rect 199088 828 199144 884
rect 198848 748 198904 804
rect 198928 748 198984 804
rect 199008 748 199064 804
rect 199088 748 199144 804
rect 198848 668 198904 724
rect 198928 668 198984 724
rect 199008 668 199064 724
rect 199088 668 199144 724
rect 199508 7688 199564 7744
rect 199588 7688 199644 7744
rect 199668 7688 199724 7744
rect 199748 7688 199804 7744
rect 199508 7642 199564 7664
rect 199588 7642 199644 7664
rect 199668 7642 199724 7664
rect 199748 7642 199804 7664
rect 199508 7608 199554 7642
rect 199554 7608 199564 7642
rect 199588 7608 199618 7642
rect 199618 7608 199630 7642
rect 199630 7608 199644 7642
rect 199668 7608 199682 7642
rect 199682 7608 199694 7642
rect 199694 7608 199724 7642
rect 199748 7608 199758 7642
rect 199758 7608 199804 7642
rect 199508 7528 199564 7584
rect 199588 7528 199644 7584
rect 199668 7528 199724 7584
rect 199748 7528 199804 7584
rect 199508 7448 199564 7504
rect 199588 7448 199644 7504
rect 199668 7448 199724 7504
rect 199748 7448 199804 7504
rect 199508 5784 199564 5840
rect 199588 5784 199644 5840
rect 199668 5784 199724 5840
rect 199748 5784 199804 5840
rect 199508 5704 199564 5760
rect 199588 5704 199644 5760
rect 199668 5704 199724 5760
rect 199748 5704 199804 5760
rect 199508 5624 199564 5680
rect 199588 5624 199644 5680
rect 199668 5624 199724 5680
rect 199748 5624 199804 5680
rect 199508 5544 199564 5600
rect 199588 5544 199644 5600
rect 199668 5544 199724 5600
rect 199748 5544 199804 5600
rect 199508 3880 199564 3936
rect 199588 3880 199644 3936
rect 199668 3880 199724 3936
rect 199748 3880 199804 3936
rect 199508 3800 199564 3856
rect 199588 3800 199644 3856
rect 199668 3800 199724 3856
rect 199748 3800 199804 3856
rect 199508 3720 199564 3776
rect 199588 3720 199644 3776
rect 199668 3720 199724 3776
rect 199748 3720 199804 3776
rect 199508 3640 199564 3696
rect 199588 3640 199644 3696
rect 199668 3640 199724 3696
rect 199748 3640 199804 3696
rect 203982 10512 204038 10568
rect 203706 10240 203762 10296
rect 203522 10104 203578 10160
rect 202970 8200 203026 8256
rect 202510 7928 202566 7984
rect 202694 7928 202750 7984
rect 204534 9968 204590 10024
rect 205454 11464 205510 11520
rect 207294 11464 207350 11520
rect 213642 11464 213698 11520
rect 214378 11484 214434 11520
rect 214378 11464 214380 11484
rect 214380 11464 214432 11484
rect 214432 11464 214434 11484
rect 205730 10684 205732 10704
rect 205732 10684 205784 10704
rect 205784 10684 205786 10704
rect 205730 10648 205786 10684
rect 205822 10512 205878 10568
rect 206190 10376 206246 10432
rect 206742 10240 206798 10296
rect 205638 10004 205640 10024
rect 205640 10004 205692 10024
rect 205692 10004 205694 10024
rect 205638 9968 205694 10004
rect 207386 10512 207442 10568
rect 207294 9968 207350 10024
rect 205546 9832 205602 9888
rect 206282 9832 206338 9888
rect 208674 10104 208730 10160
rect 210146 10276 210148 10296
rect 210148 10276 210200 10296
rect 210200 10276 210202 10296
rect 210146 10240 210202 10276
rect 210330 10396 210386 10432
rect 210330 10376 210332 10396
rect 210332 10376 210384 10396
rect 210384 10376 210386 10396
rect 210238 9832 210294 9888
rect 210238 9152 210294 9208
rect 210054 8064 210110 8120
rect 199508 248 199564 304
rect 199588 248 199644 304
rect 199668 248 199724 304
rect 199748 248 199804 304
rect 199508 168 199564 224
rect 199588 168 199644 224
rect 199668 168 199724 224
rect 199748 168 199804 224
rect 199508 88 199564 144
rect 199588 88 199644 144
rect 199668 88 199724 144
rect 199748 88 199804 144
rect 214102 10104 214158 10160
rect 215574 8472 215630 8528
rect 222198 6568 222254 6624
rect 216954 1264 217010 1320
rect 224682 8336 224738 8392
rect 219162 1128 219218 1184
rect 213734 448 213790 504
rect 228270 2760 228326 2816
rect 233422 6296 233478 6352
rect 238298 6160 238354 6216
rect 240138 4664 240194 4720
rect 242898 6024 242954 6080
rect 245014 4392 245070 4448
rect 248510 5344 248566 5400
rect 232042 1944 232098 2000
rect 251546 4256 251602 4312
rect 251454 1808 251510 1864
rect 251362 1672 251418 1728
rect 252742 4528 252798 4584
rect 254582 2488 254638 2544
rect 256330 2624 256386 2680
rect 255778 2352 255834 2408
rect 257526 2216 257582 2272
rect 258998 2080 259054 2136
rect 252558 448 252614 504
rect 254122 448 254178 504
rect 254950 448 255006 504
rect 259366 468 259422 504
rect 259366 448 259368 468
rect 259368 448 259420 468
rect 259420 448 259422 468
rect 270958 7928 271014 7984
rect 273166 1128 273222 1184
rect 278962 1128 279018 1184
rect 291198 7248 291254 7304
rect 286138 3440 286194 3496
rect 330776 11244 330832 11300
rect 330856 11244 330912 11300
rect 330936 11244 330992 11300
rect 331016 11244 331072 11300
rect 330776 11164 330832 11220
rect 330856 11164 330912 11220
rect 330936 11164 330992 11220
rect 331016 11164 331072 11220
rect 330776 11084 330832 11140
rect 330856 11084 330912 11140
rect 330936 11084 330992 11140
rect 331016 11084 331072 11140
rect 330776 11004 330832 11060
rect 330856 11004 330912 11060
rect 330936 11004 330992 11060
rect 331016 11004 331072 11060
rect 330776 8932 330832 8988
rect 330856 8932 330912 8988
rect 330936 8932 330992 8988
rect 331016 8932 331072 8988
rect 330776 8852 330832 8908
rect 330856 8852 330912 8908
rect 330936 8852 330992 8908
rect 331016 8852 331072 8908
rect 330776 8772 330832 8828
rect 330856 8772 330912 8828
rect 330936 8772 330992 8828
rect 331016 8772 331072 8828
rect 330776 8692 330832 8748
rect 330856 8692 330912 8748
rect 330936 8692 330992 8748
rect 331016 8692 331072 8748
rect 330776 7046 330822 7084
rect 330822 7046 330832 7084
rect 330856 7046 330886 7084
rect 330886 7046 330898 7084
rect 330898 7046 330912 7084
rect 330936 7046 330950 7084
rect 330950 7046 330962 7084
rect 330962 7046 330992 7084
rect 331016 7046 331026 7084
rect 331026 7046 331072 7084
rect 330776 7028 330832 7046
rect 330856 7028 330912 7046
rect 330936 7028 330992 7046
rect 331016 7028 331072 7046
rect 330776 6948 330832 7004
rect 330856 6948 330912 7004
rect 330936 6948 330992 7004
rect 331016 6948 331072 7004
rect 330776 6868 330832 6924
rect 330856 6868 330912 6924
rect 330936 6868 330992 6924
rect 331016 6868 331072 6924
rect 330776 6788 330832 6844
rect 330856 6788 330912 6844
rect 330936 6788 330992 6844
rect 331016 6788 331072 6844
rect 330776 5124 330832 5180
rect 330856 5124 330912 5180
rect 330936 5124 330992 5180
rect 331016 5124 331072 5180
rect 330776 5044 330832 5100
rect 330856 5044 330912 5100
rect 330936 5044 330992 5100
rect 331016 5044 331072 5100
rect 330776 4964 330832 5020
rect 330856 4964 330912 5020
rect 330936 4964 330992 5020
rect 331016 4964 331072 5020
rect 330776 4922 330832 4940
rect 330856 4922 330912 4940
rect 330936 4922 330992 4940
rect 331016 4922 331072 4940
rect 330776 4884 330822 4922
rect 330822 4884 330832 4922
rect 330856 4884 330886 4922
rect 330886 4884 330898 4922
rect 330898 4884 330912 4922
rect 330936 4884 330950 4922
rect 330950 4884 330962 4922
rect 330962 4884 330992 4922
rect 331016 4884 331026 4922
rect 331026 4884 331072 4922
rect 330776 3220 330832 3276
rect 330856 3220 330912 3276
rect 330936 3220 330992 3276
rect 331016 3220 331072 3276
rect 330776 3140 330832 3196
rect 330856 3140 330912 3196
rect 330936 3140 330992 3196
rect 331016 3140 331072 3196
rect 330776 3060 330832 3116
rect 330856 3060 330912 3116
rect 330936 3060 330992 3116
rect 331016 3060 331072 3116
rect 330776 2980 330832 3036
rect 330856 2980 330912 3036
rect 330936 2980 330992 3036
rect 331016 2980 331072 3036
rect 282274 1400 282330 1456
rect 283194 1420 283250 1456
rect 283194 1400 283196 1420
rect 283196 1400 283248 1420
rect 283248 1400 283250 1420
rect 291014 1128 291070 1184
rect 292210 1264 292266 1320
rect 292302 1148 292358 1184
rect 292302 1128 292304 1148
rect 292304 1128 292356 1148
rect 292356 1128 292358 1148
rect 297546 1264 297602 1320
rect 293866 484 293868 504
rect 293868 484 293920 504
rect 293920 484 293922 504
rect 293866 448 293922 484
rect 298558 448 298614 504
rect 300398 448 300454 504
rect 309046 448 309102 504
rect 311898 1264 311954 1320
rect 311070 1128 311126 1184
rect 311990 1148 312046 1184
rect 311990 1128 311992 1148
rect 311992 1128 312044 1148
rect 312044 1128 312046 1148
rect 318062 1264 318118 1320
rect 315302 448 315358 504
rect 318246 448 318302 504
rect 331436 11904 331492 11960
rect 331516 11904 331572 11960
rect 331596 11904 331652 11960
rect 331676 11904 331732 11960
rect 331436 11824 331492 11880
rect 331516 11824 331572 11880
rect 331596 11824 331652 11880
rect 331676 11824 331732 11880
rect 331436 11744 331492 11800
rect 331516 11744 331572 11800
rect 331596 11744 331652 11800
rect 331676 11744 331732 11800
rect 331436 11664 331492 11720
rect 331516 11664 331572 11720
rect 331596 11664 331652 11720
rect 331676 11664 331732 11720
rect 331436 9592 331492 9648
rect 331516 9592 331572 9648
rect 331596 9592 331652 9648
rect 331676 9592 331732 9648
rect 331436 9512 331492 9568
rect 331516 9512 331572 9568
rect 331596 9512 331652 9568
rect 331676 9512 331732 9568
rect 331436 9432 331492 9488
rect 331516 9432 331572 9488
rect 331596 9432 331652 9488
rect 331676 9432 331732 9488
rect 331436 9352 331492 9408
rect 331516 9352 331572 9408
rect 331596 9352 331652 9408
rect 331676 9352 331732 9408
rect 331436 7688 331492 7744
rect 331516 7688 331572 7744
rect 331596 7688 331652 7744
rect 331676 7688 331732 7744
rect 331436 7642 331492 7664
rect 331516 7642 331572 7664
rect 331596 7642 331652 7664
rect 331676 7642 331732 7664
rect 331436 7608 331482 7642
rect 331482 7608 331492 7642
rect 331516 7608 331546 7642
rect 331546 7608 331558 7642
rect 331558 7608 331572 7642
rect 331596 7608 331610 7642
rect 331610 7608 331622 7642
rect 331622 7608 331652 7642
rect 331676 7608 331686 7642
rect 331686 7608 331732 7642
rect 331436 7528 331492 7584
rect 331516 7528 331572 7584
rect 331596 7528 331652 7584
rect 331676 7528 331732 7584
rect 331436 7448 331492 7504
rect 331516 7448 331572 7504
rect 331596 7448 331652 7504
rect 331676 7448 331732 7504
rect 359922 11464 359978 11520
rect 363142 11484 363198 11520
rect 363142 11464 363144 11484
rect 363144 11464 363196 11484
rect 363196 11464 363198 11484
rect 359738 10784 359794 10840
rect 360566 10784 360622 10840
rect 359554 10512 359610 10568
rect 360198 10648 360254 10704
rect 360106 10376 360162 10432
rect 331436 5784 331492 5840
rect 331516 5784 331572 5840
rect 331596 5784 331652 5840
rect 331676 5784 331732 5840
rect 331436 5704 331492 5760
rect 331516 5704 331572 5760
rect 331596 5704 331652 5760
rect 331676 5704 331732 5760
rect 331436 5624 331492 5680
rect 331516 5624 331572 5680
rect 331596 5624 331652 5680
rect 331676 5624 331732 5680
rect 331436 5544 331492 5600
rect 331516 5544 331572 5600
rect 331596 5544 331652 5600
rect 331676 5544 331732 5600
rect 331436 3880 331492 3936
rect 331516 3880 331572 3936
rect 331596 3880 331652 3936
rect 331676 3880 331732 3936
rect 331436 3800 331492 3856
rect 331516 3800 331572 3856
rect 331596 3800 331652 3856
rect 331676 3800 331732 3856
rect 331436 3720 331492 3776
rect 331516 3720 331572 3776
rect 331596 3720 331652 3776
rect 331676 3720 331732 3776
rect 331436 3640 331492 3696
rect 331516 3640 331572 3696
rect 331596 3640 331652 3696
rect 331676 3640 331732 3696
rect 352930 2508 352986 2544
rect 352930 2488 352932 2508
rect 352932 2488 352984 2508
rect 352984 2488 352986 2508
rect 350354 2372 350410 2408
rect 350354 2352 350356 2372
rect 350356 2352 350408 2372
rect 350408 2352 350410 2372
rect 330776 908 330832 964
rect 330856 908 330912 964
rect 330936 908 330992 964
rect 331016 908 331072 964
rect 330776 828 330832 884
rect 330856 828 330912 884
rect 330936 828 330992 884
rect 331016 828 331072 884
rect 330776 748 330832 804
rect 330856 748 330912 804
rect 330936 748 330992 804
rect 331016 748 331072 804
rect 330776 668 330832 724
rect 330856 668 330912 724
rect 330936 668 330992 724
rect 331016 668 331072 724
rect 199508 8 199564 64
rect 199588 8 199644 64
rect 199668 8 199724 64
rect 199748 8 199804 64
rect 331436 248 331492 304
rect 331516 248 331572 304
rect 331596 248 331652 304
rect 331676 248 331732 304
rect 331436 168 331492 224
rect 331516 168 331572 224
rect 331596 168 331652 224
rect 331676 168 331732 224
rect 331436 88 331492 144
rect 331516 88 331572 144
rect 331596 88 331652 144
rect 331676 88 331732 144
rect 361302 10512 361358 10568
rect 363326 10648 363382 10704
rect 366730 10376 366786 10432
rect 390558 2352 390614 2408
rect 393962 2488 394018 2544
rect 462704 11244 462760 11300
rect 462784 11244 462840 11300
rect 462864 11244 462920 11300
rect 462944 11244 463000 11300
rect 462704 11164 462760 11220
rect 462784 11164 462840 11220
rect 462864 11164 462920 11220
rect 462944 11164 463000 11220
rect 462704 11084 462760 11140
rect 462784 11084 462840 11140
rect 462864 11084 462920 11140
rect 462944 11084 463000 11140
rect 462704 11004 462760 11060
rect 462784 11004 462840 11060
rect 462864 11004 462920 11060
rect 462944 11004 463000 11060
rect 462704 8932 462760 8988
rect 462784 8932 462840 8988
rect 462864 8932 462920 8988
rect 462944 8932 463000 8988
rect 462704 8852 462760 8908
rect 462784 8852 462840 8908
rect 462864 8852 462920 8908
rect 462944 8852 463000 8908
rect 462704 8772 462760 8828
rect 462784 8772 462840 8828
rect 462864 8772 462920 8828
rect 462944 8772 463000 8828
rect 462704 8692 462760 8748
rect 462784 8692 462840 8748
rect 462864 8692 462920 8748
rect 462944 8692 463000 8748
rect 462704 7046 462750 7084
rect 462750 7046 462760 7084
rect 462784 7046 462814 7084
rect 462814 7046 462826 7084
rect 462826 7046 462840 7084
rect 462864 7046 462878 7084
rect 462878 7046 462890 7084
rect 462890 7046 462920 7084
rect 462944 7046 462954 7084
rect 462954 7046 463000 7084
rect 462704 7028 462760 7046
rect 462784 7028 462840 7046
rect 462864 7028 462920 7046
rect 462944 7028 463000 7046
rect 462704 6948 462760 7004
rect 462784 6948 462840 7004
rect 462864 6948 462920 7004
rect 462944 6948 463000 7004
rect 462704 6868 462760 6924
rect 462784 6868 462840 6924
rect 462864 6868 462920 6924
rect 462944 6868 463000 6924
rect 462704 6788 462760 6844
rect 462784 6788 462840 6844
rect 462864 6788 462920 6844
rect 462944 6788 463000 6844
rect 462704 5124 462760 5180
rect 462784 5124 462840 5180
rect 462864 5124 462920 5180
rect 462944 5124 463000 5180
rect 462704 5044 462760 5100
rect 462784 5044 462840 5100
rect 462864 5044 462920 5100
rect 462944 5044 463000 5100
rect 462704 4964 462760 5020
rect 462784 4964 462840 5020
rect 462864 4964 462920 5020
rect 462944 4964 463000 5020
rect 462704 4922 462760 4940
rect 462784 4922 462840 4940
rect 462864 4922 462920 4940
rect 462944 4922 463000 4940
rect 462704 4884 462750 4922
rect 462750 4884 462760 4922
rect 462784 4884 462814 4922
rect 462814 4884 462826 4922
rect 462826 4884 462840 4922
rect 462864 4884 462878 4922
rect 462878 4884 462890 4922
rect 462890 4884 462920 4922
rect 462944 4884 462954 4922
rect 462954 4884 463000 4922
rect 462704 3220 462760 3276
rect 462784 3220 462840 3276
rect 462864 3220 462920 3276
rect 462944 3220 463000 3276
rect 462704 3140 462760 3196
rect 462784 3140 462840 3196
rect 462864 3140 462920 3196
rect 462944 3140 463000 3196
rect 462704 3060 462760 3116
rect 462784 3060 462840 3116
rect 462864 3060 462920 3116
rect 462944 3060 463000 3116
rect 462704 2980 462760 3036
rect 462784 2980 462840 3036
rect 462864 2980 462920 3036
rect 462944 2980 463000 3036
rect 462704 908 462760 964
rect 462784 908 462840 964
rect 462864 908 462920 964
rect 462944 908 463000 964
rect 462704 828 462760 884
rect 462784 828 462840 884
rect 462864 828 462920 884
rect 462944 828 463000 884
rect 462704 748 462760 804
rect 462784 748 462840 804
rect 462864 748 462920 804
rect 462944 748 463000 804
rect 462704 668 462760 724
rect 462784 668 462840 724
rect 462864 668 462920 724
rect 462944 668 463000 724
rect 331436 8 331492 64
rect 331516 8 331572 64
rect 331596 8 331652 64
rect 331676 8 331732 64
rect 463364 11904 463420 11960
rect 463444 11904 463500 11960
rect 463524 11904 463580 11960
rect 463604 11904 463660 11960
rect 463364 11824 463420 11880
rect 463444 11824 463500 11880
rect 463524 11824 463580 11880
rect 463604 11824 463660 11880
rect 463364 11744 463420 11800
rect 463444 11744 463500 11800
rect 463524 11744 463580 11800
rect 463604 11744 463660 11800
rect 463364 11664 463420 11720
rect 463444 11664 463500 11720
rect 463524 11664 463580 11720
rect 463604 11664 463660 11720
rect 530688 11904 530744 11960
rect 530768 11904 530824 11960
rect 530848 11904 530904 11960
rect 530928 11904 530984 11960
rect 530688 11824 530744 11880
rect 530768 11824 530824 11880
rect 530848 11824 530904 11880
rect 530928 11824 530984 11880
rect 530688 11744 530744 11800
rect 530768 11744 530824 11800
rect 530848 11744 530904 11800
rect 530928 11744 530984 11800
rect 530688 11664 530744 11720
rect 530768 11664 530824 11720
rect 530848 11664 530904 11720
rect 530928 11664 530984 11720
rect 463364 9592 463420 9648
rect 463444 9592 463500 9648
rect 463524 9592 463580 9648
rect 463604 9592 463660 9648
rect 463364 9512 463420 9568
rect 463444 9512 463500 9568
rect 463524 9512 463580 9568
rect 463604 9512 463660 9568
rect 463364 9432 463420 9488
rect 463444 9432 463500 9488
rect 463524 9432 463580 9488
rect 463604 9432 463660 9488
rect 463364 9352 463420 9408
rect 463444 9352 463500 9408
rect 463524 9352 463580 9408
rect 463604 9352 463660 9408
rect 463364 7688 463420 7744
rect 463444 7688 463500 7744
rect 463524 7688 463580 7744
rect 463604 7688 463660 7744
rect 463364 7642 463420 7664
rect 463444 7642 463500 7664
rect 463524 7642 463580 7664
rect 463604 7642 463660 7664
rect 463364 7608 463410 7642
rect 463410 7608 463420 7642
rect 463444 7608 463474 7642
rect 463474 7608 463486 7642
rect 463486 7608 463500 7642
rect 463524 7608 463538 7642
rect 463538 7608 463550 7642
rect 463550 7608 463580 7642
rect 463604 7608 463614 7642
rect 463614 7608 463660 7642
rect 463364 7528 463420 7584
rect 463444 7528 463500 7584
rect 463524 7528 463580 7584
rect 463604 7528 463660 7584
rect 463364 7448 463420 7504
rect 463444 7448 463500 7504
rect 463524 7448 463580 7504
rect 463604 7448 463660 7504
rect 463364 5784 463420 5840
rect 463444 5784 463500 5840
rect 463524 5784 463580 5840
rect 463604 5784 463660 5840
rect 463364 5704 463420 5760
rect 463444 5704 463500 5760
rect 463524 5704 463580 5760
rect 463604 5704 463660 5760
rect 463364 5624 463420 5680
rect 463444 5624 463500 5680
rect 463524 5624 463580 5680
rect 463604 5624 463660 5680
rect 463364 5544 463420 5600
rect 463444 5544 463500 5600
rect 463524 5544 463580 5600
rect 463604 5544 463660 5600
rect 463364 3880 463420 3936
rect 463444 3880 463500 3936
rect 463524 3880 463580 3936
rect 463604 3880 463660 3936
rect 463364 3800 463420 3856
rect 463444 3800 463500 3856
rect 463524 3800 463580 3856
rect 463604 3800 463660 3856
rect 463364 3720 463420 3776
rect 463444 3720 463500 3776
rect 463524 3720 463580 3776
rect 463604 3720 463660 3776
rect 463364 3640 463420 3696
rect 463444 3640 463500 3696
rect 463524 3640 463580 3696
rect 463604 3640 463660 3696
rect 530028 11244 530084 11300
rect 530108 11244 530164 11300
rect 530188 11244 530244 11300
rect 530268 11244 530324 11300
rect 530028 11164 530084 11220
rect 530108 11164 530164 11220
rect 530188 11164 530244 11220
rect 530268 11164 530324 11220
rect 530028 11084 530084 11140
rect 530108 11084 530164 11140
rect 530188 11084 530244 11140
rect 530268 11084 530324 11140
rect 530028 11004 530084 11060
rect 530108 11004 530164 11060
rect 530188 11004 530244 11060
rect 530268 11004 530324 11060
rect 530028 8932 530084 8988
rect 530108 8932 530164 8988
rect 530188 8932 530244 8988
rect 530268 8932 530324 8988
rect 530028 8852 530084 8908
rect 530108 8852 530164 8908
rect 530188 8852 530244 8908
rect 530268 8852 530324 8908
rect 530028 8772 530084 8828
rect 530108 8772 530164 8828
rect 530188 8772 530244 8828
rect 530268 8772 530324 8828
rect 530028 8692 530084 8748
rect 530108 8692 530164 8748
rect 530188 8692 530244 8748
rect 530268 8692 530324 8748
rect 530028 7028 530084 7084
rect 530108 7028 530164 7084
rect 530188 7028 530244 7084
rect 530268 7028 530324 7084
rect 530028 6948 530084 7004
rect 530108 6948 530164 7004
rect 530188 6948 530244 7004
rect 530268 6948 530324 7004
rect 530028 6868 530084 6924
rect 530108 6868 530164 6924
rect 530188 6868 530244 6924
rect 530268 6868 530324 6924
rect 530028 6788 530084 6844
rect 530108 6788 530164 6844
rect 530188 6788 530244 6844
rect 530268 6788 530324 6844
rect 530028 5124 530084 5180
rect 530108 5124 530164 5180
rect 530188 5124 530244 5180
rect 530268 5124 530324 5180
rect 530028 5044 530084 5100
rect 530108 5044 530164 5100
rect 530188 5044 530244 5100
rect 530268 5044 530324 5100
rect 530028 4964 530084 5020
rect 530108 4964 530164 5020
rect 530188 4964 530244 5020
rect 530268 4964 530324 5020
rect 530028 4884 530084 4940
rect 530108 4884 530164 4940
rect 530188 4884 530244 4940
rect 530268 4884 530324 4940
rect 530028 3220 530084 3276
rect 530108 3220 530164 3276
rect 530188 3220 530244 3276
rect 530268 3220 530324 3276
rect 530028 3140 530084 3196
rect 530108 3140 530164 3196
rect 530188 3140 530244 3196
rect 530268 3140 530324 3196
rect 530028 3060 530084 3116
rect 530108 3060 530164 3116
rect 530188 3060 530244 3116
rect 530268 3060 530324 3116
rect 530028 2980 530084 3036
rect 530108 2980 530164 3036
rect 530188 2980 530244 3036
rect 530268 2980 530324 3036
rect 463364 248 463420 304
rect 463444 248 463500 304
rect 463524 248 463580 304
rect 463604 248 463660 304
rect 463364 168 463420 224
rect 463444 168 463500 224
rect 463524 168 463580 224
rect 463604 168 463660 224
rect 463364 88 463420 144
rect 463444 88 463500 144
rect 463524 88 463580 144
rect 463604 88 463660 144
rect 530028 908 530084 964
rect 530108 908 530164 964
rect 530188 908 530244 964
rect 530268 908 530324 964
rect 530028 828 530084 884
rect 530108 828 530164 884
rect 530188 828 530244 884
rect 530268 828 530324 884
rect 530028 748 530084 804
rect 530108 748 530164 804
rect 530188 748 530244 804
rect 530268 748 530324 804
rect 530028 668 530084 724
rect 530108 668 530164 724
rect 530188 668 530244 724
rect 530268 668 530324 724
rect 530688 9592 530744 9648
rect 530768 9592 530824 9648
rect 530848 9592 530904 9648
rect 530928 9592 530984 9648
rect 530688 9512 530744 9568
rect 530768 9512 530824 9568
rect 530848 9512 530904 9568
rect 530928 9512 530984 9568
rect 530688 9432 530744 9488
rect 530768 9432 530824 9488
rect 530848 9432 530904 9488
rect 530928 9432 530984 9488
rect 530688 9352 530744 9408
rect 530768 9352 530824 9408
rect 530848 9352 530904 9408
rect 530928 9352 530984 9408
rect 530688 7688 530744 7744
rect 530768 7688 530824 7744
rect 530848 7688 530904 7744
rect 530928 7688 530984 7744
rect 530688 7608 530744 7664
rect 530768 7608 530824 7664
rect 530848 7608 530904 7664
rect 530928 7608 530984 7664
rect 530688 7528 530744 7584
rect 530768 7528 530824 7584
rect 530848 7528 530904 7584
rect 530928 7528 530984 7584
rect 530688 7448 530744 7504
rect 530768 7448 530824 7504
rect 530848 7448 530904 7504
rect 530928 7448 530984 7504
rect 530688 5784 530744 5840
rect 530768 5784 530824 5840
rect 530848 5784 530904 5840
rect 530928 5784 530984 5840
rect 530688 5704 530744 5760
rect 530768 5704 530824 5760
rect 530848 5704 530904 5760
rect 530928 5704 530984 5760
rect 530688 5624 530744 5680
rect 530768 5624 530824 5680
rect 530848 5624 530904 5680
rect 530928 5624 530984 5680
rect 530688 5544 530744 5600
rect 530768 5544 530824 5600
rect 530848 5544 530904 5600
rect 530928 5544 530984 5600
rect 530688 3880 530744 3936
rect 530768 3880 530824 3936
rect 530848 3880 530904 3936
rect 530928 3880 530984 3936
rect 530688 3800 530744 3856
rect 530768 3800 530824 3856
rect 530848 3800 530904 3856
rect 530928 3800 530984 3856
rect 530688 3720 530744 3776
rect 530768 3720 530824 3776
rect 530848 3720 530904 3776
rect 530928 3720 530984 3776
rect 530688 3640 530744 3696
rect 530768 3640 530824 3696
rect 530848 3640 530904 3696
rect 530928 3640 530984 3696
rect 530688 248 530744 304
rect 530768 248 530824 304
rect 530848 248 530904 304
rect 530928 248 530984 304
rect 530688 168 530744 224
rect 530768 168 530824 224
rect 530848 168 530904 224
rect 530928 168 530984 224
rect 530688 88 530744 144
rect 530768 88 530824 144
rect 530848 88 530904 144
rect 530928 88 530984 144
rect 463364 8 463420 64
rect 463444 8 463500 64
rect 463524 8 463580 64
rect 463604 8 463660 64
rect 530688 8 530744 64
rect 530768 8 530824 64
rect 530848 8 530904 64
rect 530928 8 530984 64
<< metal3 >>
rect -1076 11960 530996 11972
rect -1076 11904 -1064 11960
rect -1008 11904 -984 11960
rect -928 11904 -904 11960
rect -848 11904 -824 11960
rect -768 11904 67580 11960
rect 67636 11904 67660 11960
rect 67716 11904 67740 11960
rect 67796 11904 67820 11960
rect 67876 11904 199508 11960
rect 199564 11904 199588 11960
rect 199644 11904 199668 11960
rect 199724 11904 199748 11960
rect 199804 11904 331436 11960
rect 331492 11904 331516 11960
rect 331572 11904 331596 11960
rect 331652 11904 331676 11960
rect 331732 11904 463364 11960
rect 463420 11904 463444 11960
rect 463500 11904 463524 11960
rect 463580 11904 463604 11960
rect 463660 11904 530688 11960
rect 530744 11904 530768 11960
rect 530824 11904 530848 11960
rect 530904 11904 530928 11960
rect 530984 11904 530996 11960
rect -1076 11880 530996 11904
rect -1076 11824 -1064 11880
rect -1008 11824 -984 11880
rect -928 11824 -904 11880
rect -848 11824 -824 11880
rect -768 11824 67580 11880
rect 67636 11824 67660 11880
rect 67716 11824 67740 11880
rect 67796 11824 67820 11880
rect 67876 11824 199508 11880
rect 199564 11824 199588 11880
rect 199644 11824 199668 11880
rect 199724 11824 199748 11880
rect 199804 11824 331436 11880
rect 331492 11824 331516 11880
rect 331572 11824 331596 11880
rect 331652 11824 331676 11880
rect 331732 11824 463364 11880
rect 463420 11824 463444 11880
rect 463500 11824 463524 11880
rect 463580 11824 463604 11880
rect 463660 11824 530688 11880
rect 530744 11824 530768 11880
rect 530824 11824 530848 11880
rect 530904 11824 530928 11880
rect 530984 11824 530996 11880
rect -1076 11800 530996 11824
rect -1076 11744 -1064 11800
rect -1008 11744 -984 11800
rect -928 11744 -904 11800
rect -848 11744 -824 11800
rect -768 11744 67580 11800
rect 67636 11744 67660 11800
rect 67716 11744 67740 11800
rect 67796 11744 67820 11800
rect 67876 11744 199508 11800
rect 199564 11744 199588 11800
rect 199644 11744 199668 11800
rect 199724 11744 199748 11800
rect 199804 11744 331436 11800
rect 331492 11744 331516 11800
rect 331572 11744 331596 11800
rect 331652 11744 331676 11800
rect 331732 11744 463364 11800
rect 463420 11744 463444 11800
rect 463500 11744 463524 11800
rect 463580 11744 463604 11800
rect 463660 11744 530688 11800
rect 530744 11744 530768 11800
rect 530824 11744 530848 11800
rect 530904 11744 530928 11800
rect 530984 11744 530996 11800
rect -1076 11720 530996 11744
rect -1076 11664 -1064 11720
rect -1008 11664 -984 11720
rect -928 11664 -904 11720
rect -848 11664 -824 11720
rect -768 11664 67580 11720
rect 67636 11664 67660 11720
rect 67716 11664 67740 11720
rect 67796 11664 67820 11720
rect 67876 11664 199508 11720
rect 199564 11664 199588 11720
rect 199644 11664 199668 11720
rect 199724 11664 199748 11720
rect 199804 11664 331436 11720
rect 331492 11664 331516 11720
rect 331572 11664 331596 11720
rect 331652 11664 331676 11720
rect 331732 11664 463364 11720
rect 463420 11664 463444 11720
rect 463500 11664 463524 11720
rect 463580 11664 463604 11720
rect 463660 11664 530688 11720
rect 530744 11664 530768 11720
rect 530824 11664 530848 11720
rect 530904 11664 530928 11720
rect 530984 11664 530996 11720
rect -1076 11652 530996 11664
rect 199377 11522 199443 11525
rect 202045 11522 202111 11525
rect 199377 11520 202111 11522
rect 199377 11464 199382 11520
rect 199438 11464 202050 11520
rect 202106 11464 202111 11520
rect 199377 11462 202111 11464
rect 199377 11459 199443 11462
rect 202045 11459 202111 11462
rect 205449 11522 205515 11525
rect 207289 11522 207355 11525
rect 205449 11520 207355 11522
rect 205449 11464 205454 11520
rect 205510 11464 207294 11520
rect 207350 11464 207355 11520
rect 205449 11462 207355 11464
rect 205449 11459 205515 11462
rect 207289 11459 207355 11462
rect 213637 11522 213703 11525
rect 214373 11522 214439 11525
rect 213637 11520 214439 11522
rect 213637 11464 213642 11520
rect 213698 11464 214378 11520
rect 214434 11464 214439 11520
rect 213637 11462 214439 11464
rect 213637 11459 213703 11462
rect 214373 11459 214439 11462
rect 359917 11522 359983 11525
rect 363137 11522 363203 11525
rect 359917 11520 363203 11522
rect 359917 11464 359922 11520
rect 359978 11464 363142 11520
rect 363198 11464 363203 11520
rect 359917 11462 363203 11464
rect 359917 11459 359983 11462
rect 363137 11459 363203 11462
rect -416 11300 530336 11312
rect -416 11244 -404 11300
rect -348 11244 -324 11300
rect -268 11244 -244 11300
rect -188 11244 -164 11300
rect -108 11244 66920 11300
rect 66976 11244 67000 11300
rect 67056 11244 67080 11300
rect 67136 11244 67160 11300
rect 67216 11244 198848 11300
rect 198904 11244 198928 11300
rect 198984 11244 199008 11300
rect 199064 11244 199088 11300
rect 199144 11244 330776 11300
rect 330832 11244 330856 11300
rect 330912 11244 330936 11300
rect 330992 11244 331016 11300
rect 331072 11244 462704 11300
rect 462760 11244 462784 11300
rect 462840 11244 462864 11300
rect 462920 11244 462944 11300
rect 463000 11244 530028 11300
rect 530084 11244 530108 11300
rect 530164 11244 530188 11300
rect 530244 11244 530268 11300
rect 530324 11244 530336 11300
rect -416 11220 530336 11244
rect -416 11164 -404 11220
rect -348 11164 -324 11220
rect -268 11164 -244 11220
rect -188 11164 -164 11220
rect -108 11164 66920 11220
rect 66976 11164 67000 11220
rect 67056 11164 67080 11220
rect 67136 11164 67160 11220
rect 67216 11164 198848 11220
rect 198904 11164 198928 11220
rect 198984 11164 199008 11220
rect 199064 11164 199088 11220
rect 199144 11164 330776 11220
rect 330832 11164 330856 11220
rect 330912 11164 330936 11220
rect 330992 11164 331016 11220
rect 331072 11164 462704 11220
rect 462760 11164 462784 11220
rect 462840 11164 462864 11220
rect 462920 11164 462944 11220
rect 463000 11164 530028 11220
rect 530084 11164 530108 11220
rect 530164 11164 530188 11220
rect 530244 11164 530268 11220
rect 530324 11164 530336 11220
rect -416 11140 530336 11164
rect -416 11084 -404 11140
rect -348 11084 -324 11140
rect -268 11084 -244 11140
rect -188 11084 -164 11140
rect -108 11084 66920 11140
rect 66976 11084 67000 11140
rect 67056 11084 67080 11140
rect 67136 11084 67160 11140
rect 67216 11084 198848 11140
rect 198904 11084 198928 11140
rect 198984 11084 199008 11140
rect 199064 11084 199088 11140
rect 199144 11084 330776 11140
rect 330832 11084 330856 11140
rect 330912 11084 330936 11140
rect 330992 11084 331016 11140
rect 331072 11084 462704 11140
rect 462760 11084 462784 11140
rect 462840 11084 462864 11140
rect 462920 11084 462944 11140
rect 463000 11084 530028 11140
rect 530084 11084 530108 11140
rect 530164 11084 530188 11140
rect 530244 11084 530268 11140
rect 530324 11084 530336 11140
rect -416 11060 530336 11084
rect -416 11004 -404 11060
rect -348 11004 -324 11060
rect -268 11004 -244 11060
rect -188 11004 -164 11060
rect -108 11004 66920 11060
rect 66976 11004 67000 11060
rect 67056 11004 67080 11060
rect 67136 11004 67160 11060
rect 67216 11004 198848 11060
rect 198904 11004 198928 11060
rect 198984 11004 199008 11060
rect 199064 11004 199088 11060
rect 199144 11004 330776 11060
rect 330832 11004 330856 11060
rect 330912 11004 330936 11060
rect 330992 11004 331016 11060
rect 331072 11004 462704 11060
rect 462760 11004 462784 11060
rect 462840 11004 462864 11060
rect 462920 11004 462944 11060
rect 463000 11004 530028 11060
rect 530084 11004 530108 11060
rect 530164 11004 530188 11060
rect 530244 11004 530268 11060
rect 530324 11004 530336 11060
rect -416 10992 530336 11004
rect 198641 10842 198707 10845
rect 200941 10842 201007 10845
rect 198641 10840 201007 10842
rect 198641 10784 198646 10840
rect 198702 10784 200946 10840
rect 201002 10784 201007 10840
rect 198641 10782 201007 10784
rect 198641 10779 198707 10782
rect 200941 10779 201007 10782
rect 359733 10842 359799 10845
rect 360561 10842 360627 10845
rect 359733 10840 360627 10842
rect 359733 10784 359738 10840
rect 359794 10784 360566 10840
rect 360622 10784 360627 10840
rect 359733 10782 360627 10784
rect 359733 10779 359799 10782
rect 360561 10779 360627 10782
rect 199285 10706 199351 10709
rect 205725 10706 205791 10709
rect 199285 10704 205791 10706
rect 199285 10648 199290 10704
rect 199346 10648 205730 10704
rect 205786 10648 205791 10704
rect 199285 10646 205791 10648
rect 199285 10643 199351 10646
rect 205725 10643 205791 10646
rect 360193 10706 360259 10709
rect 363321 10706 363387 10709
rect 360193 10704 363387 10706
rect 360193 10648 360198 10704
rect 360254 10648 363326 10704
rect 363382 10648 363387 10704
rect 360193 10646 363387 10648
rect 360193 10643 360259 10646
rect 363321 10643 363387 10646
rect 199285 10570 199351 10573
rect 203977 10570 204043 10573
rect 199285 10568 204043 10570
rect 199285 10512 199290 10568
rect 199346 10512 203982 10568
rect 204038 10512 204043 10568
rect 199285 10510 204043 10512
rect 199285 10507 199351 10510
rect 203977 10507 204043 10510
rect 205817 10570 205883 10573
rect 207381 10570 207447 10573
rect 205817 10568 207447 10570
rect 205817 10512 205822 10568
rect 205878 10512 207386 10568
rect 207442 10512 207447 10568
rect 205817 10510 207447 10512
rect 205817 10507 205883 10510
rect 207381 10507 207447 10510
rect 359549 10570 359615 10573
rect 361297 10570 361363 10573
rect 359549 10568 361363 10570
rect 359549 10512 359554 10568
rect 359610 10512 361302 10568
rect 361358 10512 361363 10568
rect 359549 10510 361363 10512
rect 359549 10507 359615 10510
rect 361297 10507 361363 10510
rect 201493 10434 201559 10437
rect 206185 10434 206251 10437
rect 210325 10434 210391 10437
rect 201493 10432 206251 10434
rect 201493 10376 201498 10432
rect 201554 10376 206190 10432
rect 206246 10376 206251 10432
rect 201493 10374 206251 10376
rect 201493 10371 201559 10374
rect 206185 10371 206251 10374
rect 206326 10432 210391 10434
rect 206326 10376 210330 10432
rect 210386 10376 210391 10432
rect 206326 10374 210391 10376
rect 203701 10298 203767 10301
rect 206326 10298 206386 10374
rect 210325 10371 210391 10374
rect 360101 10434 360167 10437
rect 366725 10434 366791 10437
rect 360101 10432 366791 10434
rect 360101 10376 360106 10432
rect 360162 10376 366730 10432
rect 366786 10376 366791 10432
rect 360101 10374 366791 10376
rect 360101 10371 360167 10374
rect 366725 10371 366791 10374
rect 203701 10296 206386 10298
rect 203701 10240 203706 10296
rect 203762 10240 206386 10296
rect 203701 10238 206386 10240
rect 206737 10298 206803 10301
rect 210141 10298 210207 10301
rect 206737 10296 210207 10298
rect 206737 10240 206742 10296
rect 206798 10240 210146 10296
rect 210202 10240 210207 10296
rect 206737 10238 210207 10240
rect 203701 10235 203767 10238
rect 206737 10235 206803 10238
rect 210141 10235 210207 10238
rect 198641 10162 198707 10165
rect 203517 10162 203583 10165
rect 198641 10160 203583 10162
rect 198641 10104 198646 10160
rect 198702 10104 203522 10160
rect 203578 10104 203583 10160
rect 198641 10102 203583 10104
rect 198641 10099 198707 10102
rect 203517 10099 203583 10102
rect 208669 10162 208735 10165
rect 214097 10162 214163 10165
rect 208669 10160 214163 10162
rect 208669 10104 208674 10160
rect 208730 10104 214102 10160
rect 214158 10104 214163 10160
rect 208669 10102 214163 10104
rect 208669 10099 208735 10102
rect 214097 10099 214163 10102
rect 198365 10026 198431 10029
rect 204529 10026 204595 10029
rect 198365 10024 204595 10026
rect 198365 9968 198370 10024
rect 198426 9968 204534 10024
rect 204590 9968 204595 10024
rect 198365 9966 204595 9968
rect 198365 9963 198431 9966
rect 204529 9963 204595 9966
rect 205633 10026 205699 10029
rect 207289 10026 207355 10029
rect 205633 10024 207355 10026
rect 205633 9968 205638 10024
rect 205694 9968 207294 10024
rect 207350 9968 207355 10024
rect 205633 9966 207355 9968
rect 205633 9963 205699 9966
rect 207289 9963 207355 9966
rect 197813 9890 197879 9893
rect 205541 9890 205607 9893
rect 197813 9888 205607 9890
rect 197813 9832 197818 9888
rect 197874 9832 205546 9888
rect 205602 9832 205607 9888
rect 197813 9830 205607 9832
rect 197813 9827 197879 9830
rect 205541 9827 205607 9830
rect 206277 9890 206343 9893
rect 210233 9890 210299 9893
rect 206277 9888 210299 9890
rect 206277 9832 206282 9888
rect 206338 9832 210238 9888
rect 210294 9832 210299 9888
rect 206277 9830 210299 9832
rect 206277 9827 206343 9830
rect 210233 9827 210299 9830
rect -1076 9648 530996 9660
rect -1076 9592 -1064 9648
rect -1008 9592 -984 9648
rect -928 9592 -904 9648
rect -848 9592 -824 9648
rect -768 9592 67580 9648
rect 67636 9592 67660 9648
rect 67716 9592 67740 9648
rect 67796 9592 67820 9648
rect 67876 9592 199508 9648
rect 199564 9592 199588 9648
rect 199644 9592 199668 9648
rect 199724 9592 199748 9648
rect 199804 9592 331436 9648
rect 331492 9592 331516 9648
rect 331572 9592 331596 9648
rect 331652 9592 331676 9648
rect 331732 9592 463364 9648
rect 463420 9592 463444 9648
rect 463500 9592 463524 9648
rect 463580 9592 463604 9648
rect 463660 9592 530688 9648
rect 530744 9592 530768 9648
rect 530824 9592 530848 9648
rect 530904 9592 530928 9648
rect 530984 9592 530996 9648
rect -1076 9568 530996 9592
rect -1076 9512 -1064 9568
rect -1008 9512 -984 9568
rect -928 9512 -904 9568
rect -848 9512 -824 9568
rect -768 9512 67580 9568
rect 67636 9512 67660 9568
rect 67716 9512 67740 9568
rect 67796 9512 67820 9568
rect 67876 9512 199508 9568
rect 199564 9512 199588 9568
rect 199644 9512 199668 9568
rect 199724 9512 199748 9568
rect 199804 9512 331436 9568
rect 331492 9512 331516 9568
rect 331572 9512 331596 9568
rect 331652 9512 331676 9568
rect 331732 9512 463364 9568
rect 463420 9512 463444 9568
rect 463500 9512 463524 9568
rect 463580 9512 463604 9568
rect 463660 9512 530688 9568
rect 530744 9512 530768 9568
rect 530824 9512 530848 9568
rect 530904 9512 530928 9568
rect 530984 9512 530996 9568
rect -1076 9488 530996 9512
rect -1076 9432 -1064 9488
rect -1008 9432 -984 9488
rect -928 9432 -904 9488
rect -848 9432 -824 9488
rect -768 9432 67580 9488
rect 67636 9432 67660 9488
rect 67716 9432 67740 9488
rect 67796 9432 67820 9488
rect 67876 9432 199508 9488
rect 199564 9432 199588 9488
rect 199644 9432 199668 9488
rect 199724 9432 199748 9488
rect 199804 9432 331436 9488
rect 331492 9432 331516 9488
rect 331572 9432 331596 9488
rect 331652 9432 331676 9488
rect 331732 9432 463364 9488
rect 463420 9432 463444 9488
rect 463500 9432 463524 9488
rect 463580 9432 463604 9488
rect 463660 9432 530688 9488
rect 530744 9432 530768 9488
rect 530824 9432 530848 9488
rect 530904 9432 530928 9488
rect 530984 9432 530996 9488
rect -1076 9408 530996 9432
rect -1076 9352 -1064 9408
rect -1008 9352 -984 9408
rect -928 9352 -904 9408
rect -848 9352 -824 9408
rect -768 9352 67580 9408
rect 67636 9352 67660 9408
rect 67716 9352 67740 9408
rect 67796 9352 67820 9408
rect 67876 9352 199508 9408
rect 199564 9352 199588 9408
rect 199644 9352 199668 9408
rect 199724 9352 199748 9408
rect 199804 9352 331436 9408
rect 331492 9352 331516 9408
rect 331572 9352 331596 9408
rect 331652 9352 331676 9408
rect 331732 9352 463364 9408
rect 463420 9352 463444 9408
rect 463500 9352 463524 9408
rect 463580 9352 463604 9408
rect 463660 9352 530688 9408
rect 530744 9352 530768 9408
rect 530824 9352 530848 9408
rect 530904 9352 530928 9408
rect 530984 9352 530996 9408
rect -1076 9340 530996 9352
rect 103053 9210 103119 9213
rect 210233 9210 210299 9213
rect 103053 9208 210299 9210
rect 103053 9152 103058 9208
rect 103114 9152 210238 9208
rect 210294 9152 210299 9208
rect 103053 9150 210299 9152
rect 103053 9147 103119 9150
rect 210233 9147 210299 9150
rect -1076 8988 530996 9000
rect -1076 8932 -404 8988
rect -348 8932 -324 8988
rect -268 8932 -244 8988
rect -188 8932 -164 8988
rect -108 8932 66920 8988
rect 66976 8932 67000 8988
rect 67056 8932 67080 8988
rect 67136 8932 67160 8988
rect 67216 8932 198848 8988
rect 198904 8932 198928 8988
rect 198984 8932 199008 8988
rect 199064 8932 199088 8988
rect 199144 8932 330776 8988
rect 330832 8932 330856 8988
rect 330912 8932 330936 8988
rect 330992 8932 331016 8988
rect 331072 8932 462704 8988
rect 462760 8932 462784 8988
rect 462840 8932 462864 8988
rect 462920 8932 462944 8988
rect 463000 8932 530028 8988
rect 530084 8932 530108 8988
rect 530164 8932 530188 8988
rect 530244 8932 530268 8988
rect 530324 8932 530996 8988
rect -1076 8908 530996 8932
rect -1076 8852 -404 8908
rect -348 8852 -324 8908
rect -268 8852 -244 8908
rect -188 8852 -164 8908
rect -108 8852 66920 8908
rect 66976 8852 67000 8908
rect 67056 8852 67080 8908
rect 67136 8852 67160 8908
rect 67216 8852 198848 8908
rect 198904 8852 198928 8908
rect 198984 8852 199008 8908
rect 199064 8852 199088 8908
rect 199144 8852 330776 8908
rect 330832 8852 330856 8908
rect 330912 8852 330936 8908
rect 330992 8852 331016 8908
rect 331072 8852 462704 8908
rect 462760 8852 462784 8908
rect 462840 8852 462864 8908
rect 462920 8852 462944 8908
rect 463000 8852 530028 8908
rect 530084 8852 530108 8908
rect 530164 8852 530188 8908
rect 530244 8852 530268 8908
rect 530324 8852 530996 8908
rect -1076 8828 530996 8852
rect -1076 8772 -404 8828
rect -348 8772 -324 8828
rect -268 8772 -244 8828
rect -188 8772 -164 8828
rect -108 8772 66920 8828
rect 66976 8772 67000 8828
rect 67056 8772 67080 8828
rect 67136 8772 67160 8828
rect 67216 8772 198848 8828
rect 198904 8772 198928 8828
rect 198984 8772 199008 8828
rect 199064 8772 199088 8828
rect 199144 8772 330776 8828
rect 330832 8772 330856 8828
rect 330912 8772 330936 8828
rect 330992 8772 331016 8828
rect 331072 8772 462704 8828
rect 462760 8772 462784 8828
rect 462840 8772 462864 8828
rect 462920 8772 462944 8828
rect 463000 8772 530028 8828
rect 530084 8772 530108 8828
rect 530164 8772 530188 8828
rect 530244 8772 530268 8828
rect 530324 8772 530996 8828
rect -1076 8748 530996 8772
rect -1076 8692 -404 8748
rect -348 8692 -324 8748
rect -268 8692 -244 8748
rect -188 8692 -164 8748
rect -108 8692 66920 8748
rect 66976 8692 67000 8748
rect 67056 8692 67080 8748
rect 67136 8692 67160 8748
rect 67216 8692 198848 8748
rect 198904 8692 198928 8748
rect 198984 8692 199008 8748
rect 199064 8692 199088 8748
rect 199144 8692 330776 8748
rect 330832 8692 330856 8748
rect 330912 8692 330936 8748
rect 330992 8692 331016 8748
rect 331072 8692 462704 8748
rect 462760 8692 462784 8748
rect 462840 8692 462864 8748
rect 462920 8692 462944 8748
rect 463000 8692 530028 8748
rect 530084 8692 530108 8748
rect 530164 8692 530188 8748
rect 530244 8692 530268 8748
rect 530324 8692 530996 8748
rect -1076 8680 530996 8692
rect 67265 8530 67331 8533
rect 175273 8530 175339 8533
rect 67265 8528 175339 8530
rect 67265 8472 67270 8528
rect 67326 8472 175278 8528
rect 175334 8472 175339 8528
rect 67265 8470 175339 8472
rect 67265 8467 67331 8470
rect 175273 8467 175339 8470
rect 184197 8530 184263 8533
rect 215569 8530 215635 8533
rect 184197 8528 215635 8530
rect 184197 8472 184202 8528
rect 184258 8472 215574 8528
rect 215630 8472 215635 8528
rect 184197 8470 215635 8472
rect 184197 8467 184263 8470
rect 215569 8467 215635 8470
rect 172513 8394 172579 8397
rect 224677 8394 224743 8397
rect 172513 8392 224743 8394
rect 172513 8336 172518 8392
rect 172574 8336 224682 8392
rect 224738 8336 224743 8392
rect 172513 8334 224743 8336
rect 172513 8331 172579 8334
rect 224677 8331 224743 8334
rect 176653 8258 176719 8261
rect 202965 8258 203031 8261
rect 176653 8256 203031 8258
rect 176653 8200 176658 8256
rect 176714 8200 202970 8256
rect 203026 8200 203031 8256
rect 176653 8198 203031 8200
rect 176653 8195 176719 8198
rect 202965 8195 203031 8198
rect 101857 8122 101923 8125
rect 210049 8122 210115 8125
rect 101857 8120 210115 8122
rect 101857 8064 101862 8120
rect 101918 8064 210054 8120
rect 210110 8064 210115 8120
rect 101857 8062 210115 8064
rect 101857 8059 101923 8062
rect 210049 8059 210115 8062
rect 93485 7986 93551 7989
rect 202505 7986 202571 7989
rect 93485 7984 202571 7986
rect 93485 7928 93490 7984
rect 93546 7928 202510 7984
rect 202566 7928 202571 7984
rect 93485 7926 202571 7928
rect 93485 7923 93551 7926
rect 202505 7923 202571 7926
rect 202689 7986 202755 7989
rect 270953 7986 271019 7989
rect 202689 7984 271019 7986
rect 202689 7928 202694 7984
rect 202750 7928 270958 7984
rect 271014 7928 271019 7984
rect 202689 7926 271019 7928
rect 202689 7923 202755 7926
rect 270953 7923 271019 7926
rect -1076 7744 530996 7756
rect -1076 7688 -1064 7744
rect -1008 7688 -984 7744
rect -928 7688 -904 7744
rect -848 7688 -824 7744
rect -768 7688 67580 7744
rect 67636 7688 67660 7744
rect 67716 7688 67740 7744
rect 67796 7688 67820 7744
rect 67876 7688 199508 7744
rect 199564 7688 199588 7744
rect 199644 7688 199668 7744
rect 199724 7688 199748 7744
rect 199804 7688 331436 7744
rect 331492 7688 331516 7744
rect 331572 7688 331596 7744
rect 331652 7688 331676 7744
rect 331732 7688 463364 7744
rect 463420 7688 463444 7744
rect 463500 7688 463524 7744
rect 463580 7688 463604 7744
rect 463660 7688 530688 7744
rect 530744 7688 530768 7744
rect 530824 7688 530848 7744
rect 530904 7688 530928 7744
rect 530984 7688 530996 7744
rect -1076 7664 530996 7688
rect -1076 7608 -1064 7664
rect -1008 7608 -984 7664
rect -928 7608 -904 7664
rect -848 7608 -824 7664
rect -768 7608 67580 7664
rect 67636 7608 67660 7664
rect 67716 7608 67740 7664
rect 67796 7608 67820 7664
rect 67876 7608 199508 7664
rect 199564 7608 199588 7664
rect 199644 7608 199668 7664
rect 199724 7608 199748 7664
rect 199804 7608 331436 7664
rect 331492 7608 331516 7664
rect 331572 7608 331596 7664
rect 331652 7608 331676 7664
rect 331732 7608 463364 7664
rect 463420 7608 463444 7664
rect 463500 7608 463524 7664
rect 463580 7608 463604 7664
rect 463660 7608 530688 7664
rect 530744 7608 530768 7664
rect 530824 7608 530848 7664
rect 530904 7608 530928 7664
rect 530984 7608 530996 7664
rect -1076 7584 530996 7608
rect -1076 7528 -1064 7584
rect -1008 7528 -984 7584
rect -928 7528 -904 7584
rect -848 7528 -824 7584
rect -768 7528 67580 7584
rect 67636 7528 67660 7584
rect 67716 7528 67740 7584
rect 67796 7528 67820 7584
rect 67876 7528 199508 7584
rect 199564 7528 199588 7584
rect 199644 7528 199668 7584
rect 199724 7528 199748 7584
rect 199804 7528 331436 7584
rect 331492 7528 331516 7584
rect 331572 7528 331596 7584
rect 331652 7528 331676 7584
rect 331732 7528 463364 7584
rect 463420 7528 463444 7584
rect 463500 7528 463524 7584
rect 463580 7528 463604 7584
rect 463660 7528 530688 7584
rect 530744 7528 530768 7584
rect 530824 7528 530848 7584
rect 530904 7528 530928 7584
rect 530984 7528 530996 7584
rect -1076 7504 530996 7528
rect -1076 7448 -1064 7504
rect -1008 7448 -984 7504
rect -928 7448 -904 7504
rect -848 7448 -824 7504
rect -768 7448 67580 7504
rect 67636 7448 67660 7504
rect 67716 7448 67740 7504
rect 67796 7448 67820 7504
rect 67876 7448 199508 7504
rect 199564 7448 199588 7504
rect 199644 7448 199668 7504
rect 199724 7448 199748 7504
rect 199804 7448 331436 7504
rect 331492 7448 331516 7504
rect 331572 7448 331596 7504
rect 331652 7448 331676 7504
rect 331732 7448 463364 7504
rect 463420 7448 463444 7504
rect 463500 7448 463524 7504
rect 463580 7448 463604 7504
rect 463660 7448 530688 7504
rect 530744 7448 530768 7504
rect 530824 7448 530848 7504
rect 530904 7448 530928 7504
rect 530984 7448 530996 7504
rect -1076 7436 530996 7448
rect 182909 7306 182975 7309
rect 291193 7306 291259 7309
rect 182909 7304 291259 7306
rect 182909 7248 182914 7304
rect 182970 7248 291198 7304
rect 291254 7248 291259 7304
rect 182909 7246 291259 7248
rect 182909 7243 182975 7246
rect 291193 7243 291259 7246
rect -1076 7084 530996 7096
rect -1076 7028 -404 7084
rect -348 7028 -324 7084
rect -268 7028 -244 7084
rect -188 7028 -164 7084
rect -108 7028 66920 7084
rect 66976 7028 67000 7084
rect 67056 7028 67080 7084
rect 67136 7028 67160 7084
rect 67216 7028 198848 7084
rect 198904 7028 198928 7084
rect 198984 7028 199008 7084
rect 199064 7028 199088 7084
rect 199144 7028 330776 7084
rect 330832 7028 330856 7084
rect 330912 7028 330936 7084
rect 330992 7028 331016 7084
rect 331072 7028 462704 7084
rect 462760 7028 462784 7084
rect 462840 7028 462864 7084
rect 462920 7028 462944 7084
rect 463000 7028 530028 7084
rect 530084 7028 530108 7084
rect 530164 7028 530188 7084
rect 530244 7028 530268 7084
rect 530324 7028 530996 7084
rect -1076 7004 530996 7028
rect -1076 6948 -404 7004
rect -348 6948 -324 7004
rect -268 6948 -244 7004
rect -188 6948 -164 7004
rect -108 6948 66920 7004
rect 66976 6948 67000 7004
rect 67056 6948 67080 7004
rect 67136 6948 67160 7004
rect 67216 6948 198848 7004
rect 198904 6948 198928 7004
rect 198984 6948 199008 7004
rect 199064 6948 199088 7004
rect 199144 6948 330776 7004
rect 330832 6948 330856 7004
rect 330912 6948 330936 7004
rect 330992 6948 331016 7004
rect 331072 6948 462704 7004
rect 462760 6948 462784 7004
rect 462840 6948 462864 7004
rect 462920 6948 462944 7004
rect 463000 6948 530028 7004
rect 530084 6948 530108 7004
rect 530164 6948 530188 7004
rect 530244 6948 530268 7004
rect 530324 6948 530996 7004
rect -1076 6924 530996 6948
rect -1076 6868 -404 6924
rect -348 6868 -324 6924
rect -268 6868 -244 6924
rect -188 6868 -164 6924
rect -108 6868 66920 6924
rect 66976 6868 67000 6924
rect 67056 6868 67080 6924
rect 67136 6868 67160 6924
rect 67216 6868 198848 6924
rect 198904 6868 198928 6924
rect 198984 6868 199008 6924
rect 199064 6868 199088 6924
rect 199144 6868 330776 6924
rect 330832 6868 330856 6924
rect 330912 6868 330936 6924
rect 330992 6868 331016 6924
rect 331072 6868 462704 6924
rect 462760 6868 462784 6924
rect 462840 6868 462864 6924
rect 462920 6868 462944 6924
rect 463000 6868 530028 6924
rect 530084 6868 530108 6924
rect 530164 6868 530188 6924
rect 530244 6868 530268 6924
rect 530324 6868 530996 6924
rect -1076 6844 530996 6868
rect -1076 6788 -404 6844
rect -348 6788 -324 6844
rect -268 6788 -244 6844
rect -188 6788 -164 6844
rect -108 6788 66920 6844
rect 66976 6788 67000 6844
rect 67056 6788 67080 6844
rect 67136 6788 67160 6844
rect 67216 6788 198848 6844
rect 198904 6788 198928 6844
rect 198984 6788 199008 6844
rect 199064 6788 199088 6844
rect 199144 6788 330776 6844
rect 330832 6788 330856 6844
rect 330912 6788 330936 6844
rect 330992 6788 331016 6844
rect 331072 6788 462704 6844
rect 462760 6788 462784 6844
rect 462840 6788 462864 6844
rect 462920 6788 462944 6844
rect 463000 6788 530028 6844
rect 530084 6788 530108 6844
rect 530164 6788 530188 6844
rect 530244 6788 530268 6844
rect 530324 6788 530996 6844
rect -1076 6776 530996 6788
rect 114185 6626 114251 6629
rect 222193 6626 222259 6629
rect 114185 6624 222259 6626
rect 114185 6568 114190 6624
rect 114246 6568 222198 6624
rect 222254 6568 222259 6624
rect 114185 6566 222259 6568
rect 114185 6563 114251 6566
rect 222193 6563 222259 6566
rect 125501 6354 125567 6357
rect 233417 6354 233483 6357
rect 125501 6352 233483 6354
rect 125501 6296 125506 6352
rect 125562 6296 233422 6352
rect 233478 6296 233483 6352
rect 125501 6294 233483 6296
rect 125501 6291 125567 6294
rect 233417 6291 233483 6294
rect 130929 6218 130995 6221
rect 238293 6218 238359 6221
rect 130929 6216 238359 6218
rect 130929 6160 130934 6216
rect 130990 6160 238298 6216
rect 238354 6160 238359 6216
rect 130929 6158 238359 6160
rect 130929 6155 130995 6158
rect 238293 6155 238359 6158
rect 135529 6082 135595 6085
rect 242893 6082 242959 6085
rect 135529 6080 242959 6082
rect 135529 6024 135534 6080
rect 135590 6024 242898 6080
rect 242954 6024 242959 6080
rect 135529 6022 242959 6024
rect 135529 6019 135595 6022
rect 242893 6019 242959 6022
rect -1076 5840 530996 5852
rect -1076 5784 -1064 5840
rect -1008 5784 -984 5840
rect -928 5784 -904 5840
rect -848 5784 -824 5840
rect -768 5784 67580 5840
rect 67636 5784 67660 5840
rect 67716 5784 67740 5840
rect 67796 5784 67820 5840
rect 67876 5784 199508 5840
rect 199564 5784 199588 5840
rect 199644 5784 199668 5840
rect 199724 5784 199748 5840
rect 199804 5784 331436 5840
rect 331492 5784 331516 5840
rect 331572 5784 331596 5840
rect 331652 5784 331676 5840
rect 331732 5784 463364 5840
rect 463420 5784 463444 5840
rect 463500 5784 463524 5840
rect 463580 5784 463604 5840
rect 463660 5784 530688 5840
rect 530744 5784 530768 5840
rect 530824 5784 530848 5840
rect 530904 5784 530928 5840
rect 530984 5784 530996 5840
rect -1076 5760 530996 5784
rect -1076 5704 -1064 5760
rect -1008 5704 -984 5760
rect -928 5704 -904 5760
rect -848 5704 -824 5760
rect -768 5704 67580 5760
rect 67636 5704 67660 5760
rect 67716 5704 67740 5760
rect 67796 5704 67820 5760
rect 67876 5704 199508 5760
rect 199564 5704 199588 5760
rect 199644 5704 199668 5760
rect 199724 5704 199748 5760
rect 199804 5704 331436 5760
rect 331492 5704 331516 5760
rect 331572 5704 331596 5760
rect 331652 5704 331676 5760
rect 331732 5704 463364 5760
rect 463420 5704 463444 5760
rect 463500 5704 463524 5760
rect 463580 5704 463604 5760
rect 463660 5704 530688 5760
rect 530744 5704 530768 5760
rect 530824 5704 530848 5760
rect 530904 5704 530928 5760
rect 530984 5704 530996 5760
rect -1076 5680 530996 5704
rect -1076 5624 -1064 5680
rect -1008 5624 -984 5680
rect -928 5624 -904 5680
rect -848 5624 -824 5680
rect -768 5624 67580 5680
rect 67636 5624 67660 5680
rect 67716 5624 67740 5680
rect 67796 5624 67820 5680
rect 67876 5624 199508 5680
rect 199564 5624 199588 5680
rect 199644 5624 199668 5680
rect 199724 5624 199748 5680
rect 199804 5624 331436 5680
rect 331492 5624 331516 5680
rect 331572 5624 331596 5680
rect 331652 5624 331676 5680
rect 331732 5624 463364 5680
rect 463420 5624 463444 5680
rect 463500 5624 463524 5680
rect 463580 5624 463604 5680
rect 463660 5624 530688 5680
rect 530744 5624 530768 5680
rect 530824 5624 530848 5680
rect 530904 5624 530928 5680
rect 530984 5624 530996 5680
rect -1076 5600 530996 5624
rect -1076 5544 -1064 5600
rect -1008 5544 -984 5600
rect -928 5544 -904 5600
rect -848 5544 -824 5600
rect -768 5544 67580 5600
rect 67636 5544 67660 5600
rect 67716 5544 67740 5600
rect 67796 5544 67820 5600
rect 67876 5544 199508 5600
rect 199564 5544 199588 5600
rect 199644 5544 199668 5600
rect 199724 5544 199748 5600
rect 199804 5544 331436 5600
rect 331492 5544 331516 5600
rect 331572 5544 331596 5600
rect 331652 5544 331676 5600
rect 331732 5544 463364 5600
rect 463420 5544 463444 5600
rect 463500 5544 463524 5600
rect 463580 5544 463604 5600
rect 463660 5544 530688 5600
rect 530744 5544 530768 5600
rect 530824 5544 530848 5600
rect 530904 5544 530928 5600
rect 530984 5544 530996 5600
rect -1076 5532 530996 5544
rect 141325 5402 141391 5405
rect 248505 5402 248571 5405
rect 141325 5400 248571 5402
rect 141325 5344 141330 5400
rect 141386 5344 248510 5400
rect 248566 5344 248571 5400
rect 141325 5342 248571 5344
rect 141325 5339 141391 5342
rect 248505 5339 248571 5342
rect -1076 5180 530996 5192
rect -1076 5124 -404 5180
rect -348 5124 -324 5180
rect -268 5124 -244 5180
rect -188 5124 -164 5180
rect -108 5124 66920 5180
rect 66976 5124 67000 5180
rect 67056 5124 67080 5180
rect 67136 5124 67160 5180
rect 67216 5124 198848 5180
rect 198904 5124 198928 5180
rect 198984 5124 199008 5180
rect 199064 5124 199088 5180
rect 199144 5124 330776 5180
rect 330832 5124 330856 5180
rect 330912 5124 330936 5180
rect 330992 5124 331016 5180
rect 331072 5124 462704 5180
rect 462760 5124 462784 5180
rect 462840 5124 462864 5180
rect 462920 5124 462944 5180
rect 463000 5124 530028 5180
rect 530084 5124 530108 5180
rect 530164 5124 530188 5180
rect 530244 5124 530268 5180
rect 530324 5124 530996 5180
rect -1076 5100 530996 5124
rect -1076 5044 -404 5100
rect -348 5044 -324 5100
rect -268 5044 -244 5100
rect -188 5044 -164 5100
rect -108 5044 66920 5100
rect 66976 5044 67000 5100
rect 67056 5044 67080 5100
rect 67136 5044 67160 5100
rect 67216 5044 198848 5100
rect 198904 5044 198928 5100
rect 198984 5044 199008 5100
rect 199064 5044 199088 5100
rect 199144 5044 330776 5100
rect 330832 5044 330856 5100
rect 330912 5044 330936 5100
rect 330992 5044 331016 5100
rect 331072 5044 462704 5100
rect 462760 5044 462784 5100
rect 462840 5044 462864 5100
rect 462920 5044 462944 5100
rect 463000 5044 530028 5100
rect 530084 5044 530108 5100
rect 530164 5044 530188 5100
rect 530244 5044 530268 5100
rect 530324 5044 530996 5100
rect -1076 5020 530996 5044
rect -1076 4964 -404 5020
rect -348 4964 -324 5020
rect -268 4964 -244 5020
rect -188 4964 -164 5020
rect -108 4964 66920 5020
rect 66976 4964 67000 5020
rect 67056 4964 67080 5020
rect 67136 4964 67160 5020
rect 67216 4964 198848 5020
rect 198904 4964 198928 5020
rect 198984 4964 199008 5020
rect 199064 4964 199088 5020
rect 199144 4964 330776 5020
rect 330832 4964 330856 5020
rect 330912 4964 330936 5020
rect 330992 4964 331016 5020
rect 331072 4964 462704 5020
rect 462760 4964 462784 5020
rect 462840 4964 462864 5020
rect 462920 4964 462944 5020
rect 463000 4964 530028 5020
rect 530084 4964 530108 5020
rect 530164 4964 530188 5020
rect 530244 4964 530268 5020
rect 530324 4964 530996 5020
rect -1076 4940 530996 4964
rect -1076 4884 -404 4940
rect -348 4884 -324 4940
rect -268 4884 -244 4940
rect -188 4884 -164 4940
rect -108 4884 66920 4940
rect 66976 4884 67000 4940
rect 67056 4884 67080 4940
rect 67136 4884 67160 4940
rect 67216 4884 198848 4940
rect 198904 4884 198928 4940
rect 198984 4884 199008 4940
rect 199064 4884 199088 4940
rect 199144 4884 330776 4940
rect 330832 4884 330856 4940
rect 330912 4884 330936 4940
rect 330992 4884 331016 4940
rect 331072 4884 462704 4940
rect 462760 4884 462784 4940
rect 462840 4884 462864 4940
rect 462920 4884 462944 4940
rect 463000 4884 530028 4940
rect 530084 4884 530108 4940
rect 530164 4884 530188 4940
rect 530244 4884 530268 4940
rect 530324 4884 530996 4940
rect -1076 4872 530996 4884
rect 81709 4722 81775 4725
rect 125685 4722 125751 4725
rect 81709 4720 125751 4722
rect 81709 4664 81714 4720
rect 81770 4664 125690 4720
rect 125746 4664 125751 4720
rect 81709 4662 125751 4664
rect 81709 4659 81775 4662
rect 125685 4659 125751 4662
rect 133505 4722 133571 4725
rect 240133 4722 240199 4725
rect 133505 4720 240199 4722
rect 133505 4664 133510 4720
rect 133566 4664 240138 4720
rect 240194 4664 240199 4720
rect 133505 4662 240199 4664
rect 133505 4659 133571 4662
rect 240133 4659 240199 4662
rect 92381 4586 92447 4589
rect 131205 4586 131271 4589
rect 92381 4584 131271 4586
rect 92381 4528 92386 4584
rect 92442 4528 131210 4584
rect 131266 4528 131271 4584
rect 92381 4526 131271 4528
rect 92381 4523 92447 4526
rect 131205 4523 131271 4526
rect 145925 4586 145991 4589
rect 252737 4586 252803 4589
rect 145925 4584 252803 4586
rect 145925 4528 145930 4584
rect 145986 4528 252742 4584
rect 252798 4528 252803 4584
rect 145925 4526 252803 4528
rect 145925 4523 145991 4526
rect 252737 4523 252803 4526
rect 137829 4450 137895 4453
rect 245009 4450 245075 4453
rect 137829 4448 245075 4450
rect 137829 4392 137834 4448
rect 137890 4392 245014 4448
rect 245070 4392 245075 4448
rect 137829 4390 245075 4392
rect 137829 4387 137895 4390
rect 245009 4387 245075 4390
rect 144821 4314 144887 4317
rect 251541 4314 251607 4317
rect 144821 4312 251607 4314
rect 144821 4256 144826 4312
rect 144882 4256 251546 4312
rect 251602 4256 251607 4312
rect 144821 4254 251607 4256
rect 144821 4251 144887 4254
rect 251541 4251 251607 4254
rect -1076 3936 530996 3948
rect -1076 3880 -1064 3936
rect -1008 3880 -984 3936
rect -928 3880 -904 3936
rect -848 3880 -824 3936
rect -768 3880 67580 3936
rect 67636 3880 67660 3936
rect 67716 3880 67740 3936
rect 67796 3880 67820 3936
rect 67876 3880 199508 3936
rect 199564 3880 199588 3936
rect 199644 3880 199668 3936
rect 199724 3880 199748 3936
rect 199804 3880 331436 3936
rect 331492 3880 331516 3936
rect 331572 3880 331596 3936
rect 331652 3880 331676 3936
rect 331732 3880 463364 3936
rect 463420 3880 463444 3936
rect 463500 3880 463524 3936
rect 463580 3880 463604 3936
rect 463660 3880 530688 3936
rect 530744 3880 530768 3936
rect 530824 3880 530848 3936
rect 530904 3880 530928 3936
rect 530984 3880 530996 3936
rect -1076 3856 530996 3880
rect -1076 3800 -1064 3856
rect -1008 3800 -984 3856
rect -928 3800 -904 3856
rect -848 3800 -824 3856
rect -768 3800 67580 3856
rect 67636 3800 67660 3856
rect 67716 3800 67740 3856
rect 67796 3800 67820 3856
rect 67876 3800 199508 3856
rect 199564 3800 199588 3856
rect 199644 3800 199668 3856
rect 199724 3800 199748 3856
rect 199804 3800 331436 3856
rect 331492 3800 331516 3856
rect 331572 3800 331596 3856
rect 331652 3800 331676 3856
rect 331732 3800 463364 3856
rect 463420 3800 463444 3856
rect 463500 3800 463524 3856
rect 463580 3800 463604 3856
rect 463660 3800 530688 3856
rect 530744 3800 530768 3856
rect 530824 3800 530848 3856
rect 530904 3800 530928 3856
rect 530984 3800 530996 3856
rect -1076 3776 530996 3800
rect -1076 3720 -1064 3776
rect -1008 3720 -984 3776
rect -928 3720 -904 3776
rect -848 3720 -824 3776
rect -768 3720 67580 3776
rect 67636 3720 67660 3776
rect 67716 3720 67740 3776
rect 67796 3720 67820 3776
rect 67876 3720 199508 3776
rect 199564 3720 199588 3776
rect 199644 3720 199668 3776
rect 199724 3720 199748 3776
rect 199804 3720 331436 3776
rect 331492 3720 331516 3776
rect 331572 3720 331596 3776
rect 331652 3720 331676 3776
rect 331732 3720 463364 3776
rect 463420 3720 463444 3776
rect 463500 3720 463524 3776
rect 463580 3720 463604 3776
rect 463660 3720 530688 3776
rect 530744 3720 530768 3776
rect 530824 3720 530848 3776
rect 530904 3720 530928 3776
rect 530984 3720 530996 3776
rect -1076 3696 530996 3720
rect -1076 3640 -1064 3696
rect -1008 3640 -984 3696
rect -928 3640 -904 3696
rect -848 3640 -824 3696
rect -768 3640 67580 3696
rect 67636 3640 67660 3696
rect 67716 3640 67740 3696
rect 67796 3640 67820 3696
rect 67876 3640 199508 3696
rect 199564 3640 199588 3696
rect 199644 3640 199668 3696
rect 199724 3640 199748 3696
rect 199804 3640 331436 3696
rect 331492 3640 331516 3696
rect 331572 3640 331596 3696
rect 331652 3640 331676 3696
rect 331732 3640 463364 3696
rect 463420 3640 463444 3696
rect 463500 3640 463524 3696
rect 463580 3640 463604 3696
rect 463660 3640 530688 3696
rect 530744 3640 530768 3696
rect 530824 3640 530848 3696
rect 530904 3640 530928 3696
rect 530984 3640 530996 3696
rect -1076 3628 530996 3640
rect 32765 3498 32831 3501
rect 104433 3498 104499 3501
rect 32765 3496 104499 3498
rect 32765 3440 32770 3496
rect 32826 3440 104438 3496
rect 104494 3440 104499 3496
rect 32765 3438 104499 3440
rect 32765 3435 32831 3438
rect 104433 3435 104499 3438
rect 105077 3498 105143 3501
rect 105629 3498 105695 3501
rect 195973 3498 196039 3501
rect 105077 3496 196039 3498
rect 105077 3440 105082 3496
rect 105138 3440 105634 3496
rect 105690 3440 195978 3496
rect 196034 3440 196039 3496
rect 105077 3438 196039 3440
rect 105077 3435 105143 3438
rect 105629 3435 105695 3438
rect 195973 3435 196039 3438
rect 196157 3498 196223 3501
rect 286133 3498 286199 3501
rect 196157 3496 286199 3498
rect 196157 3440 196162 3496
rect 196218 3440 286138 3496
rect 286194 3440 286199 3496
rect 196157 3438 286199 3440
rect 196157 3435 196223 3438
rect 286133 3435 286199 3438
rect -1076 3276 530996 3288
rect -1076 3220 -404 3276
rect -348 3220 -324 3276
rect -268 3220 -244 3276
rect -188 3220 -164 3276
rect -108 3220 66920 3276
rect 66976 3220 67000 3276
rect 67056 3220 67080 3276
rect 67136 3220 67160 3276
rect 67216 3220 198848 3276
rect 198904 3220 198928 3276
rect 198984 3220 199008 3276
rect 199064 3220 199088 3276
rect 199144 3220 330776 3276
rect 330832 3220 330856 3276
rect 330912 3220 330936 3276
rect 330992 3220 331016 3276
rect 331072 3220 462704 3276
rect 462760 3220 462784 3276
rect 462840 3220 462864 3276
rect 462920 3220 462944 3276
rect 463000 3220 530028 3276
rect 530084 3220 530108 3276
rect 530164 3220 530188 3276
rect 530244 3220 530268 3276
rect 530324 3220 530996 3276
rect -1076 3196 530996 3220
rect -1076 3140 -404 3196
rect -348 3140 -324 3196
rect -268 3140 -244 3196
rect -188 3140 -164 3196
rect -108 3140 66920 3196
rect 66976 3140 67000 3196
rect 67056 3140 67080 3196
rect 67136 3140 67160 3196
rect 67216 3140 198848 3196
rect 198904 3140 198928 3196
rect 198984 3140 199008 3196
rect 199064 3140 199088 3196
rect 199144 3140 330776 3196
rect 330832 3140 330856 3196
rect 330912 3140 330936 3196
rect 330992 3140 331016 3196
rect 331072 3140 462704 3196
rect 462760 3140 462784 3196
rect 462840 3140 462864 3196
rect 462920 3140 462944 3196
rect 463000 3140 530028 3196
rect 530084 3140 530108 3196
rect 530164 3140 530188 3196
rect 530244 3140 530268 3196
rect 530324 3140 530996 3196
rect -1076 3116 530996 3140
rect -1076 3060 -404 3116
rect -348 3060 -324 3116
rect -268 3060 -244 3116
rect -188 3060 -164 3116
rect -108 3060 66920 3116
rect 66976 3060 67000 3116
rect 67056 3060 67080 3116
rect 67136 3060 67160 3116
rect 67216 3060 198848 3116
rect 198904 3060 198928 3116
rect 198984 3060 199008 3116
rect 199064 3060 199088 3116
rect 199144 3060 330776 3116
rect 330832 3060 330856 3116
rect 330912 3060 330936 3116
rect 330992 3060 331016 3116
rect 331072 3060 462704 3116
rect 462760 3060 462784 3116
rect 462840 3060 462864 3116
rect 462920 3060 462944 3116
rect 463000 3060 530028 3116
rect 530084 3060 530108 3116
rect 530164 3060 530188 3116
rect 530244 3060 530268 3116
rect 530324 3060 530996 3116
rect -1076 3036 530996 3060
rect -1076 2980 -404 3036
rect -348 2980 -324 3036
rect -268 2980 -244 3036
rect -188 2980 -164 3036
rect -108 2980 66920 3036
rect 66976 2980 67000 3036
rect 67056 2980 67080 3036
rect 67136 2980 67160 3036
rect 67216 2980 198848 3036
rect 198904 2980 198928 3036
rect 198984 2980 199008 3036
rect 199064 2980 199088 3036
rect 199144 2980 330776 3036
rect 330832 2980 330856 3036
rect 330912 2980 330936 3036
rect 330992 2980 331016 3036
rect 331072 2980 462704 3036
rect 462760 2980 462784 3036
rect 462840 2980 462864 3036
rect 462920 2980 462944 3036
rect 463000 2980 530028 3036
rect 530084 2980 530108 3036
rect 530164 2980 530188 3036
rect 530244 2980 530268 3036
rect 530324 2980 530996 3036
rect -1076 2968 530996 2980
rect 55949 2818 56015 2821
rect 112989 2818 113055 2821
rect 55949 2816 113055 2818
rect 55949 2760 55954 2816
rect 56010 2760 112994 2816
rect 113050 2760 113055 2816
rect 55949 2758 113055 2760
rect 55949 2755 56015 2758
rect 112989 2755 113055 2758
rect 113173 2818 113239 2821
rect 119337 2818 119403 2821
rect 113173 2816 119403 2818
rect 113173 2760 113178 2816
rect 113234 2760 119342 2816
rect 119398 2760 119403 2816
rect 113173 2758 119403 2760
rect 113173 2755 113239 2758
rect 119337 2755 119403 2758
rect 121085 2818 121151 2821
rect 228265 2818 228331 2821
rect 121085 2816 228331 2818
rect 121085 2760 121090 2816
rect 121146 2760 228270 2816
rect 228326 2760 228331 2816
rect 121085 2758 228331 2760
rect 121085 2755 121151 2758
rect 228265 2755 228331 2758
rect 48957 2682 49023 2685
rect 156689 2682 156755 2685
rect 48957 2680 156755 2682
rect 48957 2624 48962 2680
rect 49018 2624 156694 2680
rect 156750 2624 156755 2680
rect 48957 2622 156755 2624
rect 48957 2619 49023 2622
rect 156689 2619 156755 2622
rect 164141 2682 164207 2685
rect 256325 2682 256391 2685
rect 164141 2680 256391 2682
rect 164141 2624 164146 2680
rect 164202 2624 256330 2680
rect 256386 2624 256391 2680
rect 164141 2622 256391 2624
rect 164141 2619 164207 2622
rect 256325 2619 256391 2622
rect 41229 2546 41295 2549
rect 149053 2546 149119 2549
rect 41229 2544 149119 2546
rect 41229 2488 41234 2544
rect 41290 2488 149058 2544
rect 149114 2488 149119 2544
rect 41229 2486 149119 2488
rect 41229 2483 41295 2486
rect 149053 2483 149119 2486
rect 158897 2546 158963 2549
rect 254577 2546 254643 2549
rect 158897 2544 254643 2546
rect 158897 2488 158902 2544
rect 158958 2488 254582 2544
rect 254638 2488 254643 2544
rect 158897 2486 254643 2488
rect 158897 2483 158963 2486
rect 254577 2483 254643 2486
rect 352925 2546 352991 2549
rect 393957 2546 394023 2549
rect 352925 2544 394023 2546
rect 352925 2488 352930 2544
rect 352986 2488 393962 2544
rect 394018 2488 394023 2544
rect 352925 2486 394023 2488
rect 352925 2483 352991 2486
rect 393957 2483 394023 2486
rect 28349 2410 28415 2413
rect 136633 2410 136699 2413
rect 28349 2408 136699 2410
rect 28349 2352 28354 2408
rect 28410 2352 136638 2408
rect 136694 2352 136699 2408
rect 28349 2350 136699 2352
rect 28349 2347 28415 2350
rect 136633 2347 136699 2350
rect 146845 2410 146911 2413
rect 255773 2410 255839 2413
rect 146845 2408 255839 2410
rect 146845 2352 146850 2408
rect 146906 2352 255778 2408
rect 255834 2352 255839 2408
rect 146845 2350 255839 2352
rect 146845 2347 146911 2350
rect 255773 2347 255839 2350
rect 350349 2410 350415 2413
rect 390553 2410 390619 2413
rect 350349 2408 390619 2410
rect 350349 2352 350354 2408
rect 350410 2352 390558 2408
rect 390614 2352 390619 2408
rect 350349 2350 390619 2352
rect 350349 2347 350415 2350
rect 390553 2347 390619 2350
rect 99005 2274 99071 2277
rect 111885 2274 111951 2277
rect 99005 2272 111951 2274
rect 99005 2216 99010 2272
rect 99066 2216 111890 2272
rect 111946 2216 111951 2272
rect 99005 2214 111951 2216
rect 99005 2211 99071 2214
rect 111885 2211 111951 2214
rect 169293 2274 169359 2277
rect 257521 2274 257587 2277
rect 169293 2272 257587 2274
rect 169293 2216 169298 2272
rect 169354 2216 257526 2272
rect 257582 2216 257587 2272
rect 169293 2214 257587 2216
rect 169293 2211 169359 2214
rect 257521 2211 257587 2214
rect 64413 2138 64479 2141
rect 171225 2138 171291 2141
rect 64413 2136 171291 2138
rect 64413 2080 64418 2136
rect 64474 2080 171230 2136
rect 171286 2080 171291 2136
rect 64413 2078 171291 2080
rect 64413 2075 64479 2078
rect 171225 2075 171291 2078
rect 174445 2138 174511 2141
rect 258993 2138 259059 2141
rect 174445 2136 259059 2138
rect 174445 2080 174450 2136
rect 174506 2080 258998 2136
rect 259054 2080 259059 2136
rect 174445 2078 259059 2080
rect 174445 2075 174511 2078
rect 258993 2075 259059 2078
rect 99373 2002 99439 2005
rect 112345 2002 112411 2005
rect 99373 2000 112411 2002
rect 99373 1944 99378 2000
rect 99434 1944 112350 2000
rect 112406 1944 112411 2000
rect 99373 1942 112411 1944
rect 99373 1939 99439 1942
rect 112345 1939 112411 1942
rect 118601 2002 118667 2005
rect 124489 2002 124555 2005
rect 118601 2000 124555 2002
rect 118601 1944 118606 2000
rect 118662 1944 124494 2000
rect 124550 1944 124555 2000
rect 118601 1942 124555 1944
rect 118601 1939 118667 1942
rect 124489 1939 124555 1942
rect 126237 2002 126303 2005
rect 232037 2002 232103 2005
rect 126237 2000 232103 2002
rect 126237 1944 126242 2000
rect 126298 1944 232042 2000
rect 232098 1944 232103 2000
rect 126237 1942 232103 1944
rect 126237 1939 126303 1942
rect 232037 1939 232103 1942
rect 95325 1866 95391 1869
rect 190453 1866 190519 1869
rect 95325 1864 190519 1866
rect 95325 1808 95330 1864
rect 95386 1808 190458 1864
rect 190514 1808 190519 1864
rect 95325 1806 190519 1808
rect 95325 1803 95391 1806
rect 190453 1803 190519 1806
rect 191097 1866 191163 1869
rect 251449 1866 251515 1869
rect 191097 1864 251515 1866
rect 191097 1808 191102 1864
rect 191158 1808 251454 1864
rect 251510 1808 251515 1864
rect 191097 1806 251515 1808
rect 191097 1803 191163 1806
rect 251449 1803 251515 1806
rect 72141 1730 72207 1733
rect 158713 1730 158779 1733
rect 72141 1728 158779 1730
rect 72141 1672 72146 1728
rect 72202 1672 158718 1728
rect 158774 1672 158779 1728
rect 72141 1670 158779 1672
rect 72141 1667 72207 1670
rect 158713 1667 158779 1670
rect 168189 1730 168255 1733
rect 178033 1730 178099 1733
rect 168189 1728 178099 1730
rect 168189 1672 168194 1728
rect 168250 1672 178038 1728
rect 178094 1672 178099 1728
rect 168189 1670 178099 1672
rect 168189 1667 168255 1670
rect 178033 1667 178099 1670
rect 178677 1730 178743 1733
rect 187325 1730 187391 1733
rect 251357 1730 251423 1733
rect 178677 1728 186330 1730
rect 178677 1672 178682 1728
rect 178738 1672 186330 1728
rect 178677 1670 186330 1672
rect 178677 1667 178743 1670
rect 79869 1594 79935 1597
rect 186129 1594 186195 1597
rect 79869 1592 186195 1594
rect 79869 1536 79874 1592
rect 79930 1536 186134 1592
rect 186190 1536 186195 1592
rect 79869 1534 186195 1536
rect 186270 1594 186330 1670
rect 187325 1728 251423 1730
rect 187325 1672 187330 1728
rect 187386 1672 251362 1728
rect 251418 1672 251423 1728
rect 187325 1670 251423 1672
rect 187325 1667 187391 1670
rect 251357 1667 251423 1670
rect 189073 1594 189139 1597
rect 195145 1594 195211 1597
rect 186270 1592 189139 1594
rect 186270 1536 189078 1592
rect 189134 1536 189139 1592
rect 186270 1534 189139 1536
rect 79869 1531 79935 1534
rect 186129 1531 186195 1534
rect 189073 1531 189139 1534
rect 189214 1592 195211 1594
rect 189214 1536 195150 1592
rect 195206 1536 195211 1592
rect 189214 1534 195211 1536
rect 87321 1458 87387 1461
rect 96613 1458 96679 1461
rect 87321 1456 96679 1458
rect 87321 1400 87326 1456
rect 87382 1400 96618 1456
rect 96674 1400 96679 1456
rect 87321 1398 96679 1400
rect 87321 1395 87387 1398
rect 96613 1395 96679 1398
rect 98821 1458 98887 1461
rect 101121 1458 101187 1461
rect 98821 1456 101187 1458
rect 98821 1400 98826 1456
rect 98882 1400 101126 1456
rect 101182 1400 101187 1456
rect 98821 1398 101187 1400
rect 98821 1395 98887 1398
rect 101121 1395 101187 1398
rect 108297 1458 108363 1461
rect 114553 1458 114619 1461
rect 108297 1456 114619 1458
rect 108297 1400 108302 1456
rect 108358 1400 114558 1456
rect 114614 1400 114619 1456
rect 108297 1398 114619 1400
rect 108297 1395 108363 1398
rect 114553 1395 114619 1398
rect 119521 1458 119587 1461
rect 127065 1458 127131 1461
rect 119521 1456 127131 1458
rect 119521 1400 119526 1456
rect 119582 1400 127070 1456
rect 127126 1400 127131 1456
rect 119521 1398 127131 1400
rect 119521 1395 119587 1398
rect 127065 1395 127131 1398
rect 130469 1458 130535 1461
rect 135253 1458 135319 1461
rect 130469 1456 135319 1458
rect 130469 1400 130474 1456
rect 130530 1400 135258 1456
rect 135314 1400 135319 1456
rect 130469 1398 135319 1400
rect 130469 1395 130535 1398
rect 135253 1395 135319 1398
rect 146385 1458 146451 1461
rect 150525 1458 150591 1461
rect 146385 1456 150591 1458
rect 146385 1400 146390 1456
rect 146446 1400 150530 1456
rect 150586 1400 150591 1456
rect 146385 1398 150591 1400
rect 146385 1395 146451 1398
rect 150525 1395 150591 1398
rect 154665 1458 154731 1461
rect 156965 1458 157031 1461
rect 154665 1456 157031 1458
rect 154665 1400 154670 1456
rect 154726 1400 156970 1456
rect 157026 1400 157031 1456
rect 154665 1398 157031 1400
rect 154665 1395 154731 1398
rect 156965 1395 157031 1398
rect 157149 1458 157215 1461
rect 168373 1458 168439 1461
rect 157149 1456 168439 1458
rect 157149 1400 157154 1456
rect 157210 1400 168378 1456
rect 168434 1400 168439 1456
rect 157149 1398 168439 1400
rect 157149 1395 157215 1398
rect 168373 1395 168439 1398
rect 168557 1458 168623 1461
rect 173065 1458 173131 1461
rect 168557 1456 173131 1458
rect 168557 1400 168562 1456
rect 168618 1400 173070 1456
rect 173126 1400 173131 1456
rect 168557 1398 173131 1400
rect 168557 1395 168623 1398
rect 173065 1395 173131 1398
rect 176377 1458 176443 1461
rect 183553 1458 183619 1461
rect 176377 1456 183619 1458
rect 176377 1400 176382 1456
rect 176438 1400 183558 1456
rect 183614 1400 183619 1456
rect 176377 1398 183619 1400
rect 176377 1395 176443 1398
rect 183553 1395 183619 1398
rect 183921 1458 183987 1461
rect 189214 1458 189274 1534
rect 195145 1531 195211 1534
rect 183921 1456 189274 1458
rect 183921 1400 183926 1456
rect 183982 1400 189274 1456
rect 183921 1398 189274 1400
rect 191741 1458 191807 1461
rect 195145 1458 195211 1461
rect 191741 1456 195211 1458
rect 191741 1400 191746 1456
rect 191802 1400 195150 1456
rect 195206 1400 195211 1456
rect 191741 1398 195211 1400
rect 183921 1395 183987 1398
rect 191741 1395 191807 1398
rect 195145 1395 195211 1398
rect 282269 1458 282335 1461
rect 283189 1458 283255 1461
rect 282269 1456 283255 1458
rect 282269 1400 282274 1456
rect 282330 1400 283194 1456
rect 283250 1400 283255 1456
rect 282269 1398 283255 1400
rect 282269 1395 282335 1398
rect 283189 1395 283255 1398
rect 86861 1322 86927 1325
rect 94773 1322 94839 1325
rect 86861 1320 94839 1322
rect 86861 1264 86866 1320
rect 86922 1264 94778 1320
rect 94834 1264 94839 1320
rect 86861 1262 94839 1264
rect 86861 1259 86927 1262
rect 94773 1259 94839 1262
rect 97533 1322 97599 1325
rect 100753 1322 100819 1325
rect 97533 1320 100819 1322
rect 97533 1264 97538 1320
rect 97594 1264 100758 1320
rect 100814 1264 100819 1320
rect 97533 1262 100819 1264
rect 97533 1259 97599 1262
rect 100753 1259 100819 1262
rect 100937 1322 101003 1325
rect 108849 1322 108915 1325
rect 114737 1322 114803 1325
rect 100937 1320 108915 1322
rect 100937 1264 100942 1320
rect 100998 1264 108854 1320
rect 108910 1264 108915 1320
rect 100937 1262 108915 1264
rect 100937 1259 101003 1262
rect 108849 1259 108915 1262
rect 108990 1320 114803 1322
rect 108990 1264 114742 1320
rect 114798 1264 114803 1320
rect 108990 1262 114803 1264
rect 68093 1186 68159 1189
rect 69841 1186 69907 1189
rect 68093 1184 69907 1186
rect 68093 1128 68098 1184
rect 68154 1128 69846 1184
rect 69902 1128 69907 1184
rect 68093 1126 69907 1128
rect 68093 1123 68159 1126
rect 69841 1123 69907 1126
rect 81341 1186 81407 1189
rect 84009 1186 84075 1189
rect 81341 1184 84075 1186
rect 81341 1128 81346 1184
rect 81402 1128 84014 1184
rect 84070 1128 84075 1184
rect 81341 1126 84075 1128
rect 81341 1123 81407 1126
rect 84009 1123 84075 1126
rect 90173 1186 90239 1189
rect 96705 1186 96771 1189
rect 90173 1184 96771 1186
rect 90173 1128 90178 1184
rect 90234 1128 96710 1184
rect 96766 1128 96771 1184
rect 90173 1126 96771 1128
rect 90173 1123 90239 1126
rect 96705 1123 96771 1126
rect 97901 1186 97967 1189
rect 108990 1186 109050 1262
rect 114737 1259 114803 1262
rect 117957 1322 118023 1325
rect 216949 1322 217015 1325
rect 117957 1320 217015 1322
rect 117957 1264 117962 1320
rect 118018 1264 216954 1320
rect 217010 1264 217015 1320
rect 117957 1262 217015 1264
rect 117957 1259 118023 1262
rect 216949 1259 217015 1262
rect 292205 1322 292271 1325
rect 297541 1322 297607 1325
rect 292205 1320 297607 1322
rect 292205 1264 292210 1320
rect 292266 1264 297546 1320
rect 297602 1264 297607 1320
rect 292205 1262 297607 1264
rect 292205 1259 292271 1262
rect 297541 1259 297607 1262
rect 311893 1322 311959 1325
rect 318057 1322 318123 1325
rect 311893 1320 318123 1322
rect 311893 1264 311898 1320
rect 311954 1264 318062 1320
rect 318118 1264 318123 1320
rect 311893 1262 318123 1264
rect 311893 1259 311959 1262
rect 318057 1259 318123 1262
rect 97901 1184 109050 1186
rect 97901 1128 97906 1184
rect 97962 1128 109050 1184
rect 97901 1126 109050 1128
rect 111885 1186 111951 1189
rect 115105 1186 115171 1189
rect 111885 1184 115171 1186
rect 111885 1128 111890 1184
rect 111946 1128 115110 1184
rect 115166 1128 115171 1184
rect 111885 1126 115171 1128
rect 97901 1123 97967 1126
rect 111885 1123 111951 1126
rect 115105 1123 115171 1126
rect 118509 1186 118575 1189
rect 118785 1186 118851 1189
rect 118509 1184 118851 1186
rect 118509 1128 118514 1184
rect 118570 1128 118790 1184
rect 118846 1128 118851 1184
rect 118509 1126 118851 1128
rect 118509 1123 118575 1126
rect 118785 1123 118851 1126
rect 120165 1186 120231 1189
rect 219157 1186 219223 1189
rect 120165 1184 219223 1186
rect 120165 1128 120170 1184
rect 120226 1128 219162 1184
rect 219218 1128 219223 1184
rect 120165 1126 219223 1128
rect 120165 1123 120231 1126
rect 219157 1123 219223 1126
rect 273161 1186 273227 1189
rect 278957 1186 279023 1189
rect 273161 1184 279023 1186
rect 273161 1128 273166 1184
rect 273222 1128 278962 1184
rect 279018 1128 279023 1184
rect 273161 1126 279023 1128
rect 273161 1123 273227 1126
rect 278957 1123 279023 1126
rect 291009 1186 291075 1189
rect 292297 1186 292363 1189
rect 291009 1184 292363 1186
rect 291009 1128 291014 1184
rect 291070 1128 292302 1184
rect 292358 1128 292363 1184
rect 291009 1126 292363 1128
rect 291009 1123 291075 1126
rect 292297 1123 292363 1126
rect 311065 1186 311131 1189
rect 311985 1186 312051 1189
rect 311065 1184 312051 1186
rect 311065 1128 311070 1184
rect 311126 1128 311990 1184
rect 312046 1128 312051 1184
rect 311065 1126 312051 1128
rect 311065 1123 311131 1126
rect 311985 1123 312051 1126
rect -416 964 530336 976
rect -416 908 -404 964
rect -348 908 -324 964
rect -268 908 -244 964
rect -188 908 -164 964
rect -108 908 66920 964
rect 66976 908 67000 964
rect 67056 908 67080 964
rect 67136 908 67160 964
rect 67216 908 198848 964
rect 198904 908 198928 964
rect 198984 908 199008 964
rect 199064 908 199088 964
rect 199144 908 330776 964
rect 330832 908 330856 964
rect 330912 908 330936 964
rect 330992 908 331016 964
rect 331072 908 462704 964
rect 462760 908 462784 964
rect 462840 908 462864 964
rect 462920 908 462944 964
rect 463000 908 530028 964
rect 530084 908 530108 964
rect 530164 908 530188 964
rect 530244 908 530268 964
rect 530324 908 530336 964
rect -416 884 530336 908
rect -416 828 -404 884
rect -348 828 -324 884
rect -268 828 -244 884
rect -188 828 -164 884
rect -108 828 66920 884
rect 66976 828 67000 884
rect 67056 828 67080 884
rect 67136 828 67160 884
rect 67216 828 198848 884
rect 198904 828 198928 884
rect 198984 828 199008 884
rect 199064 828 199088 884
rect 199144 828 330776 884
rect 330832 828 330856 884
rect 330912 828 330936 884
rect 330992 828 331016 884
rect 331072 828 462704 884
rect 462760 828 462784 884
rect 462840 828 462864 884
rect 462920 828 462944 884
rect 463000 828 530028 884
rect 530084 828 530108 884
rect 530164 828 530188 884
rect 530244 828 530268 884
rect 530324 828 530336 884
rect -416 804 530336 828
rect -416 748 -404 804
rect -348 748 -324 804
rect -268 748 -244 804
rect -188 748 -164 804
rect -108 748 66920 804
rect 66976 748 67000 804
rect 67056 748 67080 804
rect 67136 748 67160 804
rect 67216 748 198848 804
rect 198904 748 198928 804
rect 198984 748 199008 804
rect 199064 748 199088 804
rect 199144 748 330776 804
rect 330832 748 330856 804
rect 330912 748 330936 804
rect 330992 748 331016 804
rect 331072 748 462704 804
rect 462760 748 462784 804
rect 462840 748 462864 804
rect 462920 748 462944 804
rect 463000 748 530028 804
rect 530084 748 530108 804
rect 530164 748 530188 804
rect 530244 748 530268 804
rect 530324 748 530336 804
rect -416 724 530336 748
rect -416 668 -404 724
rect -348 668 -324 724
rect -268 668 -244 724
rect -188 668 -164 724
rect -108 668 66920 724
rect 66976 668 67000 724
rect 67056 668 67080 724
rect 67136 668 67160 724
rect 67216 668 198848 724
rect 198904 668 198928 724
rect 198984 668 199008 724
rect 199064 668 199088 724
rect 199144 668 330776 724
rect 330832 668 330856 724
rect 330912 668 330936 724
rect 330992 668 331016 724
rect 331072 668 462704 724
rect 462760 668 462784 724
rect 462840 668 462864 724
rect 462920 668 462944 724
rect 463000 668 530028 724
rect 530084 668 530108 724
rect 530164 668 530188 724
rect 530244 668 530268 724
rect 530324 668 530336 724
rect -416 656 530336 668
rect 89161 506 89227 509
rect 94681 506 94747 509
rect 89161 504 94747 506
rect 89161 448 89166 504
rect 89222 448 94686 504
rect 94742 448 94747 504
rect 89161 446 94747 448
rect 89161 443 89227 446
rect 94681 443 94747 446
rect 97901 506 97967 509
rect 103605 506 103671 509
rect 97901 504 103671 506
rect 97901 448 97906 504
rect 97962 448 103610 504
rect 103666 448 103671 504
rect 97901 446 103671 448
rect 97901 443 97967 446
rect 103605 443 103671 446
rect 108849 506 108915 509
rect 109125 506 109191 509
rect 108849 504 109191 506
rect 108849 448 108854 504
rect 108910 448 109130 504
rect 109186 448 109191 504
rect 108849 446 109191 448
rect 108849 443 108915 446
rect 109125 443 109191 446
rect 110689 506 110755 509
rect 114737 506 114803 509
rect 110689 504 114803 506
rect 110689 448 110694 504
rect 110750 448 114742 504
rect 114798 448 114803 504
rect 110689 446 114803 448
rect 110689 443 110755 446
rect 114737 443 114803 446
rect 116025 506 116091 509
rect 213729 506 213795 509
rect 116025 504 213795 506
rect 116025 448 116030 504
rect 116086 448 213734 504
rect 213790 448 213795 504
rect 116025 446 213795 448
rect 116025 443 116091 446
rect 213729 443 213795 446
rect 252553 506 252619 509
rect 254117 506 254183 509
rect 252553 504 254183 506
rect 252553 448 252558 504
rect 252614 448 254122 504
rect 254178 448 254183 504
rect 252553 446 254183 448
rect 252553 443 252619 446
rect 254117 443 254183 446
rect 254945 506 255011 509
rect 259361 506 259427 509
rect 254945 504 259427 506
rect 254945 448 254950 504
rect 255006 448 259366 504
rect 259422 448 259427 504
rect 254945 446 259427 448
rect 254945 443 255011 446
rect 259361 443 259427 446
rect 293861 506 293927 509
rect 298553 506 298619 509
rect 293861 504 298619 506
rect 293861 448 293866 504
rect 293922 448 298558 504
rect 298614 448 298619 504
rect 293861 446 298619 448
rect 293861 443 293927 446
rect 298553 443 298619 446
rect 300393 506 300459 509
rect 309041 506 309107 509
rect 300393 504 309107 506
rect 300393 448 300398 504
rect 300454 448 309046 504
rect 309102 448 309107 504
rect 300393 446 309107 448
rect 300393 443 300459 446
rect 309041 443 309107 446
rect 315297 506 315363 509
rect 318241 506 318307 509
rect 315297 504 318307 506
rect 315297 448 315302 504
rect 315358 448 318246 504
rect 318302 448 318307 504
rect 315297 446 318307 448
rect 315297 443 315363 446
rect 318241 443 318307 446
rect -1076 304 530996 316
rect -1076 248 -1064 304
rect -1008 248 -984 304
rect -928 248 -904 304
rect -848 248 -824 304
rect -768 248 67580 304
rect 67636 248 67660 304
rect 67716 248 67740 304
rect 67796 248 67820 304
rect 67876 248 199508 304
rect 199564 248 199588 304
rect 199644 248 199668 304
rect 199724 248 199748 304
rect 199804 248 331436 304
rect 331492 248 331516 304
rect 331572 248 331596 304
rect 331652 248 331676 304
rect 331732 248 463364 304
rect 463420 248 463444 304
rect 463500 248 463524 304
rect 463580 248 463604 304
rect 463660 248 530688 304
rect 530744 248 530768 304
rect 530824 248 530848 304
rect 530904 248 530928 304
rect 530984 248 530996 304
rect -1076 224 530996 248
rect -1076 168 -1064 224
rect -1008 168 -984 224
rect -928 168 -904 224
rect -848 168 -824 224
rect -768 168 67580 224
rect 67636 168 67660 224
rect 67716 168 67740 224
rect 67796 168 67820 224
rect 67876 168 199508 224
rect 199564 168 199588 224
rect 199644 168 199668 224
rect 199724 168 199748 224
rect 199804 168 331436 224
rect 331492 168 331516 224
rect 331572 168 331596 224
rect 331652 168 331676 224
rect 331732 168 463364 224
rect 463420 168 463444 224
rect 463500 168 463524 224
rect 463580 168 463604 224
rect 463660 168 530688 224
rect 530744 168 530768 224
rect 530824 168 530848 224
rect 530904 168 530928 224
rect 530984 168 530996 224
rect -1076 144 530996 168
rect -1076 88 -1064 144
rect -1008 88 -984 144
rect -928 88 -904 144
rect -848 88 -824 144
rect -768 88 67580 144
rect 67636 88 67660 144
rect 67716 88 67740 144
rect 67796 88 67820 144
rect 67876 88 199508 144
rect 199564 88 199588 144
rect 199644 88 199668 144
rect 199724 88 199748 144
rect 199804 88 331436 144
rect 331492 88 331516 144
rect 331572 88 331596 144
rect 331652 88 331676 144
rect 331732 88 463364 144
rect 463420 88 463444 144
rect 463500 88 463524 144
rect 463580 88 463604 144
rect 463660 88 530688 144
rect 530744 88 530768 144
rect 530824 88 530848 144
rect 530904 88 530928 144
rect 530984 88 530996 144
rect -1076 64 530996 88
rect -1076 8 -1064 64
rect -1008 8 -984 64
rect -928 8 -904 64
rect -848 8 -824 64
rect -768 8 67580 64
rect 67636 8 67660 64
rect 67716 8 67740 64
rect 67796 8 67820 64
rect 67876 8 199508 64
rect 199564 8 199588 64
rect 199644 8 199668 64
rect 199724 8 199748 64
rect 199804 8 331436 64
rect 331492 8 331516 64
rect 331572 8 331596 64
rect 331652 8 331676 64
rect 331732 8 463364 64
rect 463420 8 463444 64
rect 463500 8 463524 64
rect 463580 8 463604 64
rect 463660 8 530688 64
rect 530744 8 530768 64
rect 530824 8 530848 64
rect 530904 8 530928 64
rect 530984 8 530996 64
rect -1076 -4 530996 8
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[0\].u_buf_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[1\].u_buf_A
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[2\].u_buf_A
timestamp 1676037725
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[3\].u_buf_A
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[4\].u_buf_A
timestamp 1676037725
transform -1 0 6716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[5\].u_buf_A
timestamp 1676037725
transform -1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[6\].u_buf_A
timestamp 1676037725
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[7\].u_buf_A
timestamp 1676037725
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[8\].u_buf_A
timestamp 1676037725
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[9\].u_buf_A
timestamp 1676037725
transform -1 0 11500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[10\].u_buf_A
timestamp 1676037725
transform -1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[11\].u_buf_A
timestamp 1676037725
transform 1 0 14260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[12\].u_buf_A
timestamp 1676037725
transform 1 0 17940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[13\].u_buf_A
timestamp 1676037725
transform -1 0 16652 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[14\].u_buf_A
timestamp 1676037725
transform -1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[15\].u_buf_A
timestamp 1676037725
transform 1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[16\].u_buf_A
timestamp 1676037725
transform 1 0 23092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[17\].u_buf_A
timestamp 1676037725
transform -1 0 21804 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[18\].u_buf_A
timestamp 1676037725
transform -1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[19\].u_buf_A
timestamp 1676037725
transform 1 0 24564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[20\].u_buf_A
timestamp 1676037725
transform 1 0 28244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[21\].u_buf_A
timestamp 1676037725
transform -1 0 26956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[22\].u_buf_A
timestamp 1676037725
transform -1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[23\].u_buf_A
timestamp 1676037725
transform 1 0 29716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[24\].u_buf_A
timestamp 1676037725
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[25\].u_buf_A
timestamp 1676037725
transform -1 0 32108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[26\].u_buf_A
timestamp 1676037725
transform -1 0 35052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[27\].u_buf_A
timestamp 1676037725
transform 1 0 35972 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[28\].u_buf_A
timestamp 1676037725
transform -1 0 37628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[29\].u_buf_A
timestamp 1676037725
transform -1 0 37260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[30\].u_buf_A
timestamp 1676037725
transform 1 0 41124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[31\].u_buf_A
timestamp 1676037725
transform 1 0 40204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[32\].u_buf_A
timestamp 1676037725
transform -1 0 42964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[33\].u_buf_A
timestamp 1676037725
transform 1 0 43700 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[34\].u_buf_A
timestamp 1676037725
transform -1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[35\].u_buf_A
timestamp 1676037725
transform 1 0 45356 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[36\].u_buf_A
timestamp 1676037725
transform 1 0 48852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[37\].u_buf_A
timestamp 1676037725
transform -1 0 47748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[38\].u_buf_A
timestamp 1676037725
transform -1 0 50692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[39\].u_buf_A
timestamp 1676037725
transform 1 0 51428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[40\].u_buf_A
timestamp 1676037725
transform -1 0 53268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[41\].u_buf_A
timestamp 1676037725
transform -1 0 52900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[42\].u_buf_A
timestamp 1676037725
transform 1 0 56580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[43\].u_buf_A
timestamp 1676037725
transform 1 0 55660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[44\].u_buf_A
timestamp 1676037725
transform -1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[45\].u_buf_A
timestamp 1676037725
transform 1 0 59156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[46\].u_buf_A
timestamp 1676037725
transform -1 0 60168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[47\].u_buf_A
timestamp 1676037725
transform 1 0 60812 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[48\].u_buf_A
timestamp 1676037725
transform 1 0 64308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[49\].u_buf_A
timestamp 1676037725
transform -1 0 63204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[50\].u_buf_A
timestamp 1676037725
transform -1 0 66148 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[51\].u_buf_A
timestamp 1676037725
transform 1 0 66884 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[52\].u_buf_A
timestamp 1676037725
transform -1 0 68724 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[53\].u_buf_A
timestamp 1676037725
transform -1 0 68356 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[54\].u_buf_A
timestamp 1676037725
transform 1 0 72036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[55\].u_buf_A
timestamp 1676037725
transform 1 0 71116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[56\].u_buf_A
timestamp 1676037725
transform -1 0 73876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[57\].u_buf_A
timestamp 1676037725
transform 1 0 74612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[58\].u_buf_A
timestamp 1676037725
transform -1 0 75624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[59\].u_buf_A
timestamp 1676037725
transform 1 0 76268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[60\].u_buf_A
timestamp 1676037725
transform 1 0 79764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[61\].u_buf_A
timestamp 1676037725
transform -1 0 78660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[62\].u_buf_A
timestamp 1676037725
transform -1 0 81604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[63\].u_buf_A
timestamp 1676037725
transform 1 0 82340 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[64\].u_buf_A
timestamp 1676037725
transform -1 0 84180 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[65\].u_buf_A
timestamp 1676037725
transform -1 0 83812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[66\].u_buf_A
timestamp 1676037725
transform 1 0 87492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[67\].u_buf_A
timestamp 1676037725
transform 1 0 86572 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[68\].u_buf_A
timestamp 1676037725
transform -1 0 89332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[69\].u_buf_A
timestamp 1676037725
transform 1 0 90068 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[70\].u_buf_A
timestamp 1676037725
transform -1 0 91080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[71\].u_buf_A
timestamp 1676037725
transform 1 0 91724 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[72\].u_buf_A
timestamp 1676037725
transform 1 0 95220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[73\].u_buf_A
timestamp 1676037725
transform -1 0 94116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[74\].u_buf_A
timestamp 1676037725
transform -1 0 97060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[75\].u_buf_A
timestamp 1676037725
transform 1 0 97796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[76\].u_buf_A
timestamp 1676037725
transform -1 0 99636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[77\].u_buf_A
timestamp 1676037725
transform -1 0 99268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[78\].u_buf_A
timestamp 1676037725
transform 1 0 102948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[79\].u_buf_A
timestamp 1676037725
transform 1 0 102028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[80\].u_buf_A
timestamp 1676037725
transform -1 0 104788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[81\].u_buf_A
timestamp 1676037725
transform 1 0 105524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[82\].u_buf_A
timestamp 1676037725
transform -1 0 106536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[83\].u_buf_A
timestamp 1676037725
transform 1 0 107180 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[84\].u_buf_A
timestamp 1676037725
transform 1 0 110676 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[85\].u_buf_A
timestamp 1676037725
transform -1 0 109572 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[86\].u_buf_A
timestamp 1676037725
transform -1 0 112516 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[87\].u_buf_A
timestamp 1676037725
transform 1 0 113252 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[88\].u_buf_A
timestamp 1676037725
transform -1 0 115092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[89\].u_buf_A
timestamp 1676037725
transform -1 0 114724 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[90\].u_buf_A
timestamp 1676037725
transform 1 0 118404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[91\].u_buf_A
timestamp 1676037725
transform 1 0 117484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[92\].u_buf_A
timestamp 1676037725
transform -1 0 120244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[93\].u_buf_A
timestamp 1676037725
transform 1 0 120980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[94\].u_buf_A
timestamp 1676037725
transform -1 0 121992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[95\].u_buf_A
timestamp 1676037725
transform 1 0 122636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[96\].u_buf_A
timestamp 1676037725
transform 1 0 126132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[97\].u_buf_A
timestamp 1676037725
transform -1 0 125028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[98\].u_buf_A
timestamp 1676037725
transform -1 0 127972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[99\].u_buf_A
timestamp 1676037725
transform 1 0 128708 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[100\].u_buf_A
timestamp 1676037725
transform -1 0 131468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[101\].u_buf_A
timestamp 1676037725
transform -1 0 131468 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[102\].u_buf_A
timestamp 1676037725
transform 1 0 133860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[103\].u_buf_A
timestamp 1676037725
transform -1 0 134044 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[104\].u_buf_A
timestamp 1676037725
transform -1 0 136620 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[105\].u_buf_A
timestamp 1676037725
transform 1 0 136436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[106\].u_buf_A
timestamp 1676037725
transform -1 0 138092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[107\].u_buf_A
timestamp 1676037725
transform 1 0 141588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[108\].u_buf_A
timestamp 1676037725
transform -1 0 143244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[109\].u_buf_A
timestamp 1676037725
transform 1 0 146740 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[110\].u_buf_A
timestamp 1676037725
transform -1 0 148396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[111\].u_buf_A
timestamp 1676037725
transform 1 0 151892 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[112\].u_buf_A
timestamp 1676037725
transform -1 0 153548 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[113\].u_buf_A
timestamp 1676037725
transform 1 0 157044 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[114\].u_buf_A
timestamp 1676037725
transform -1 0 158700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[115\].u_buf_A
timestamp 1676037725
transform 1 0 162196 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[116\].u_buf_A
timestamp 1676037725
transform -1 0 163852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[117\].u_buf_A
timestamp 1676037725
transform 1 0 167348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[118\].u_buf_A
timestamp 1676037725
transform -1 0 169004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[119\].u_buf_A
timestamp 1676037725
transform 1 0 172500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[120\].u_buf_A
timestamp 1676037725
transform -1 0 174156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[121\].u_buf_A
timestamp 1676037725
transform 1 0 177652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[122\].u_buf_A
timestamp 1676037725
transform -1 0 179308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[123\].u_buf_A
timestamp 1676037725
transform 1 0 182804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[124\].u_buf_A
timestamp 1676037725
transform -1 0 184460 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[125\].u_buf_A
timestamp 1676037725
transform 1 0 187956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[126\].u_buf_A
timestamp 1676037725
transform -1 0 189612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[127\].u_buf_A
timestamp 1676037725
transform 1 0 193108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[128\].u_buf_A
timestamp 1676037725
transform -1 0 194764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[129\].u_buf_A
timestamp 1676037725
transform 1 0 198260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[130\].u_buf_A
timestamp 1676037725
transform -1 0 200100 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[131\].u_buf_A
timestamp 1676037725
transform 1 0 203412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[132\].u_buf_A
timestamp 1676037725
transform -1 0 205252 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[133\].u_buf_A
timestamp 1676037725
transform 1 0 208564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[134\].u_buf_A
timestamp 1676037725
transform -1 0 210404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[135\].u_buf_A
timestamp 1676037725
transform 1 0 213716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[136\].u_buf_A
timestamp 1676037725
transform -1 0 215556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[137\].u_buf_A
timestamp 1676037725
transform 1 0 218868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[138\].u_buf_A
timestamp 1676037725
transform -1 0 220708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[139\].u_buf_A
timestamp 1676037725
transform 1 0 224020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[140\].u_buf_A
timestamp 1676037725
transform -1 0 225860 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[141\].u_buf_A
timestamp 1676037725
transform 1 0 229172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[142\].u_buf_A
timestamp 1676037725
transform 1 0 231748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[143\].u_buf_A
timestamp 1676037725
transform 1 0 234324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[144\].u_buf_A
timestamp 1676037725
transform 1 0 236900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[145\].u_buf_A
timestamp 1676037725
transform 1 0 239476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[146\].u_buf_A
timestamp 1676037725
transform 1 0 242052 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[147\].u_buf_A
timestamp 1676037725
transform 1 0 244628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[148\].u_buf_A
timestamp 1676037725
transform 1 0 247204 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[149\].u_buf_A
timestamp 1676037725
transform 1 0 249780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[150\].u_buf_A
timestamp 1676037725
transform 1 0 252356 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[151\].u_buf_A
timestamp 1676037725
transform 1 0 254932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[152\].u_buf_A
timestamp 1676037725
transform 1 0 257508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[153\].u_buf_A
timestamp 1676037725
transform 1 0 260084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[154\].u_buf_A
timestamp 1676037725
transform 1 0 262660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[155\].u_buf_A
timestamp 1676037725
transform 1 0 265236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[156\].u_buf_A
timestamp 1676037725
transform 1 0 267812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[157\].u_buf_A
timestamp 1676037725
transform 1 0 270388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[158\].u_buf_A
timestamp 1676037725
transform 1 0 272964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[159\].u_buf_A
timestamp 1676037725
transform 1 0 275540 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[160\].u_buf_A
timestamp 1676037725
transform 1 0 278116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[161\].u_buf_A
timestamp 1676037725
transform 1 0 280692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[162\].u_buf_A
timestamp 1676037725
transform 1 0 283268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[163\].u_buf_A
timestamp 1676037725
transform 1 0 285844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[164\].u_buf_A
timestamp 1676037725
transform 1 0 288420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[165\].u_buf_A
timestamp 1676037725
transform 1 0 290996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[166\].u_buf_A
timestamp 1676037725
transform 1 0 293572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[167\].u_buf_A
timestamp 1676037725
transform 1 0 296148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[168\].u_buf_A
timestamp 1676037725
transform 1 0 298724 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[169\].u_buf_A
timestamp 1676037725
transform 1 0 301300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[170\].u_buf_A
timestamp 1676037725
transform 1 0 303876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[171\].u_buf_A
timestamp 1676037725
transform 1 0 306452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[172\].u_buf_A
timestamp 1676037725
transform 1 0 309028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[173\].u_buf_A
timestamp 1676037725
transform 1 0 311604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[174\].u_buf_A
timestamp 1676037725
transform 1 0 314180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[175\].u_buf_A
timestamp 1676037725
transform 1 0 316756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[176\].u_buf_A
timestamp 1676037725
transform 1 0 319332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[177\].u_buf_A
timestamp 1676037725
transform 1 0 321908 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[178\].u_buf_A
timestamp 1676037725
transform 1 0 324484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[179\].u_buf_A
timestamp 1676037725
transform 1 0 327060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[180\].u_buf_A
timestamp 1676037725
transform 1 0 329636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[181\].u_buf_A
timestamp 1676037725
transform 1 0 332212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[182\].u_buf_A
timestamp 1676037725
transform 1 0 334788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[183\].u_buf_A
timestamp 1676037725
transform 1 0 337364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[184\].u_buf_A
timestamp 1676037725
transform 1 0 339940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[185\].u_buf_A
timestamp 1676037725
transform 1 0 342516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[186\].u_buf_A
timestamp 1676037725
transform 1 0 345092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[187\].u_buf_A
timestamp 1676037725
transform 1 0 347668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[188\].u_buf_A
timestamp 1676037725
transform 1 0 350244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[189\].u_buf_A
timestamp 1676037725
transform 1 0 352820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[190\].u_buf_A
timestamp 1676037725
transform 1 0 355396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[191\].u_buf_A
timestamp 1676037725
transform 1 0 357972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[192\].u_buf_A
timestamp 1676037725
transform 1 0 360548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[193\].u_buf_A
timestamp 1676037725
transform 1 0 363124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[194\].u_buf_A
timestamp 1676037725
transform 1 0 365700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[195\].u_buf_A
timestamp 1676037725
transform 1 0 368276 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[196\].u_buf_A
timestamp 1676037725
transform 1 0 370852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[197\].u_buf_A
timestamp 1676037725
transform 1 0 373428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[198\].u_buf_A
timestamp 1676037725
transform 1 0 376004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[199\].u_buf_A
timestamp 1676037725
transform 1 0 378580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[200\].u_buf_A
timestamp 1676037725
transform 1 0 381156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[201\].u_buf_A
timestamp 1676037725
transform 1 0 383732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[202\].u_buf_A
timestamp 1676037725
transform 1 0 386308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[203\].u_buf_A
timestamp 1676037725
transform 1 0 388884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[204\].u_buf_A
timestamp 1676037725
transform 1 0 391460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[205\].u_buf_A
timestamp 1676037725
transform 1 0 394036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[206\].u_buf_A
timestamp 1676037725
transform 1 0 396612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[207\].u_buf_A
timestamp 1676037725
transform 1 0 399188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[208\].u_buf_A
timestamp 1676037725
transform 1 0 401764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[209\].u_buf_A
timestamp 1676037725
transform 1 0 404340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[210\].u_buf_A
timestamp 1676037725
transform 1 0 406916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[211\].u_buf_A
timestamp 1676037725
transform 1 0 409492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[212\].u_buf_A
timestamp 1676037725
transform 1 0 412068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[213\].u_buf_A
timestamp 1676037725
transform 1 0 414644 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[214\].u_buf_A
timestamp 1676037725
transform 1 0 417220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[215\].u_buf_A
timestamp 1676037725
transform 1 0 419796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[216\].u_buf_A
timestamp 1676037725
transform 1 0 422372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[217\].u_buf_A
timestamp 1676037725
transform 1 0 424948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[218\].u_buf_A
timestamp 1676037725
transform 1 0 427524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[219\].u_buf_A
timestamp 1676037725
transform 1 0 430100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[220\].u_buf_A
timestamp 1676037725
transform 1 0 432676 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[221\].u_buf_A
timestamp 1676037725
transform 1 0 435252 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[222\].u_buf_A
timestamp 1676037725
transform 1 0 437828 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[223\].u_buf_A
timestamp 1676037725
transform 1 0 440404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[224\].u_buf_A
timestamp 1676037725
transform 1 0 442980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[225\].u_buf_A
timestamp 1676037725
transform 1 0 445556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[226\].u_buf_A
timestamp 1676037725
transform 1 0 448132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[227\].u_buf_A
timestamp 1676037725
transform 1 0 450708 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[228\].u_buf_A
timestamp 1676037725
transform 1 0 453284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[229\].u_buf_A
timestamp 1676037725
transform 1 0 455860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[230\].u_buf_A
timestamp 1676037725
transform 1 0 458436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[231\].u_buf_A
timestamp 1676037725
transform 1 0 461012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[232\].u_buf_A
timestamp 1676037725
transform 1 0 463588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[233\].u_buf_A
timestamp 1676037725
transform 1 0 466164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[234\].u_buf_A
timestamp 1676037725
transform 1 0 468740 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[235\].u_buf_A
timestamp 1676037725
transform 1 0 471316 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[236\].u_buf_A
timestamp 1676037725
transform 1 0 473892 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[237\].u_buf_A
timestamp 1676037725
transform 1 0 476468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[238\].u_buf_A
timestamp 1676037725
transform 1 0 479044 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[239\].u_buf_A
timestamp 1676037725
transform 1 0 481620 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[240\].u_buf_A
timestamp 1676037725
transform 1 0 484196 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[241\].u_buf_A
timestamp 1676037725
transform 1 0 485852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[242\].u_buf_A
timestamp 1676037725
transform 1 0 488428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[243\].u_buf_A
timestamp 1676037725
transform 1 0 491004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[244\].u_buf_A
timestamp 1676037725
transform 1 0 493580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[245\].u_buf_A
timestamp 1676037725
transform 1 0 496156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[246\].u_buf_A
timestamp 1676037725
transform 1 0 498732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[247\].u_buf_A
timestamp 1676037725
transform 1 0 501308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[248\].u_buf_A
timestamp 1676037725
transform 1 0 503884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[249\].u_buf_A
timestamp 1676037725
transform 1 0 506460 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[250\].u_buf_A
timestamp 1676037725
transform 1 0 509036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[251\].u_buf_A
timestamp 1676037725
transform 1 0 511612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_u_rp\[252\].u_buf_A
timestamp 1676037725
transform -1 0 514372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire1_A
timestamp 1676037725
transform -1 0 95404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire2_A
timestamp 1676037725
transform 1 0 146648 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire3_A
timestamp 1676037725
transform 1 0 145452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire4_A
timestamp 1676037725
transform 1 0 143980 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire5_A
timestamp 1676037725
transform 1 0 144992 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire6_A
timestamp 1676037725
transform 1 0 143152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire7_A
timestamp 1676037725
transform -1 0 142140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire8_A
timestamp 1676037725
transform 1 0 140484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire9_A
timestamp 1676037725
transform 1 0 141128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire10_A
timestamp 1676037725
transform -1 0 139840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire11_A
timestamp 1676037725
transform -1 0 138368 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire12_A
timestamp 1676037725
transform 1 0 136988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire13_A
timestamp 1676037725
transform 1 0 137724 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire14_A
timestamp 1676037725
transform -1 0 136344 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire15_A
timestamp 1676037725
transform -1 0 94208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire16_A
timestamp 1676037725
transform -1 0 135516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire17_A
timestamp 1676037725
transform -1 0 133768 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire18_A
timestamp 1676037725
transform 1 0 134136 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire19_A
timestamp 1676037725
transform 1 0 132664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire20_A
timestamp 1676037725
transform -1 0 131744 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire21_A
timestamp 1676037725
transform -1 0 130272 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire22_A
timestamp 1676037725
transform 1 0 131192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire23_A
timestamp 1676037725
transform 1 0 94300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire24_A
timestamp 1676037725
transform 1 0 129536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire25_A
timestamp 1676037725
transform 1 0 128156 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire26_A
timestamp 1676037725
transform 1 0 126592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire27_A
timestamp 1676037725
transform -1 0 127788 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire28_A
timestamp 1676037725
transform 1 0 125672 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire29_A
timestamp 1676037725
transform -1 0 125028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire30_A
timestamp 1676037725
transform 1 0 92276 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire31_A
timestamp 1676037725
transform 1 0 123188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire32_A
timestamp 1676037725
transform 1 0 123832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire33_A
timestamp 1676037725
transform 1 0 122636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire34_A
timestamp 1676037725
transform -1 0 121532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire35_A
timestamp 1676037725
transform -1 0 120336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire36_A
timestamp 1676037725
transform 1 0 120428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire37_A
timestamp 1676037725
transform -1 0 119048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire38_A
timestamp 1676037725
transform -1 0 92920 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire39_A
timestamp 1676037725
transform 1 0 117576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire40_A
timestamp 1676037725
transform -1 0 116840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire41_A
timestamp 1676037725
transform 1 0 117116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire42_A
timestamp 1676037725
transform -1 0 115644 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire43_A
timestamp 1676037725
transform 1 0 114724 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire44_A
timestamp 1676037725
transform -1 0 113528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire45_A
timestamp 1676037725
transform 1 0 113252 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire46_A
timestamp 1676037725
transform -1 0 91816 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire47_A
timestamp 1676037725
transform 1 0 111688 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire48_A
timestamp 1676037725
transform -1 0 111688 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire49_A
timestamp 1676037725
transform -1 0 109848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire50_A
timestamp 1676037725
transform 1 0 109756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire51_A
timestamp 1676037725
transform -1 0 108836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire52_A
timestamp 1676037725
transform -1 0 107548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire53_A
timestamp 1676037725
transform -1 0 108192 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire54_A
timestamp 1676037725
transform -1 0 106536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire55_A
timestamp 1676037725
transform 1 0 105064 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire56_A
timestamp 1676037725
transform 1 0 104420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire57_A
timestamp 1676037725
transform -1 0 103408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire58_A
timestamp 1676037725
transform 1 0 102580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire59_A
timestamp 1676037725
transform -1 0 101384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire60_A
timestamp 1676037725
transform 1 0 90528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire61_A
timestamp 1676037725
transform -1 0 101200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire62_A
timestamp 1676037725
transform 1 0 100740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire63_A
timestamp 1676037725
transform 1 0 99452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire64_A
timestamp 1676037725
transform -1 0 98532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire65_A
timestamp 1676037725
transform 1 0 98624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire66_A
timestamp 1676037725
transform 1 0 270480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire67_A
timestamp 1676037725
transform -1 0 97796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire68_A
timestamp 1676037725
transform 1 0 269652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire69_A
timestamp 1676037725
transform 1 0 268364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire70_A
timestamp 1676037725
transform -1 0 266984 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire71_A
timestamp 1676037725
transform 1 0 265972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire72_A
timestamp 1676037725
transform 1 0 264316 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire73_A
timestamp 1676037725
transform -1 0 263304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire74_A
timestamp 1676037725
transform 1 0 262292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire75_A
timestamp 1676037725
transform 1 0 260728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire76_A
timestamp 1676037725
transform 1 0 259900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire77_A
timestamp 1676037725
transform -1 0 259164 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire78_A
timestamp 1676037725
transform -1 0 96876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire79_A
timestamp 1676037725
transform 1 0 257508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire80_A
timestamp 1676037725
transform 1 0 256312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire81_A
timestamp 1676037725
transform -1 0 254748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire82_A
timestamp 1676037725
transform 1 0 253920 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire83_A
timestamp 1676037725
transform -1 0 252540 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire84_A
timestamp 1676037725
transform 1 0 96600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire85_A
timestamp 1676037725
transform -1 0 251436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire86_A
timestamp 1676037725
transform 1 0 249596 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire89_A
timestamp 1676037725
transform 1 0 147476 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire90_A
timestamp 1676037725
transform 1 0 148212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire91_A
timestamp 1676037725
transform -1 0 91080 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire92_A
timestamp 1676037725
transform -1 0 236900 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire93_A
timestamp 1676037725
transform -1 0 233404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire94_A
timestamp 1676037725
transform -1 0 229172 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire95_A
timestamp 1676037725
transform -1 0 225676 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire96_A
timestamp 1676037725
transform 1 0 122452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire97_A
timestamp 1676037725
transform -1 0 221444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire98_A
timestamp 1676037725
transform -1 0 218868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire99_A
timestamp 1676037725
transform -1 0 213900 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire100_A
timestamp 1676037725
transform -1 0 211140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire101_A
timestamp 1676037725
transform -1 0 206356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire102_A
timestamp 1676037725
transform -1 0 203688 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire103_A
timestamp 1676037725
transform -1 0 199088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire104_A
timestamp 1676037725
transform -1 0 195960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire105_A
timestamp 1676037725
transform -1 0 191544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire106_A
timestamp 1676037725
transform 1 0 188140 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire107_A
timestamp 1676037725
transform -1 0 184460 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire108_A
timestamp 1676037725
transform 1 0 180504 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire109_A
timestamp 1676037725
transform 1 0 176180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire110_A
timestamp 1676037725
transform 1 0 172960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire111_A
timestamp 1676037725
transform 1 0 168820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire112_A
timestamp 1676037725
transform -1 0 165600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire113_A
timestamp 1676037725
transform 1 0 161000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire114_A
timestamp 1676037725
transform -1 0 157964 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire115_A
timestamp 1676037725
transform 1 0 153364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire116_A
timestamp 1676037725
transform -1 0 150052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire117_A
timestamp 1676037725
transform 1 0 114724 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire118_A
timestamp 1676037725
transform -1 0 145820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire119_A
timestamp 1676037725
transform -1 0 142784 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire120_A
timestamp 1676037725
transform 1 0 137908 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire121_A
timestamp 1676037725
transform 1 0 132756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire122_A
timestamp 1676037725
transform -1 0 384100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire123_A
timestamp 1676037725
transform -1 0 381708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire124_A
timestamp 1676037725
transform -1 0 379224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire125_A
timestamp 1676037725
transform -1 0 376832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire126_A
timestamp 1676037725
transform -1 0 374348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire127_A
timestamp 1676037725
transform -1 0 371588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire128_A
timestamp 1676037725
transform -1 0 369932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire129_A
timestamp 1676037725
transform -1 0 367356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire130_A
timestamp 1676037725
transform -1 0 364780 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire131_A
timestamp 1676037725
transform -1 0 362204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire132_A
timestamp 1676037725
transform -1 0 359628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire133_A
timestamp 1676037725
transform -1 0 357972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire134_A
timestamp 1676037725
transform -1 0 355396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire135_A
timestamp 1676037725
transform -1 0 352820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire136_A
timestamp 1676037725
transform -1 0 350244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire137_A
timestamp 1676037725
transform -1 0 347668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire138_A
timestamp 1676037725
transform -1 0 345368 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire139_A
timestamp 1676037725
transform -1 0 342792 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire140_A
timestamp 1676037725
transform -1 0 340216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire141_A
timestamp 1676037725
transform 1 0 337364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire142_A
timestamp 1676037725
transform 1 0 332396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire143_A
timestamp 1676037725
transform 1 0 327428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire144_A
timestamp 1676037725
transform 1 0 322368 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire145_A
timestamp 1676037725
transform -1 0 317584 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire146_A
timestamp 1676037725
transform -1 0 312524 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire147_A
timestamp 1676037725
transform 1 0 127604 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire148_A
timestamp 1676037725
transform -1 0 307556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire149_A
timestamp 1676037725
transform -1 0 302496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire150_A
timestamp 1676037725
transform 1 0 297620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire151_A
timestamp 1676037725
transform 1 0 292468 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire152_A
timestamp 1676037725
transform 1 0 287316 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire153_A
timestamp 1676037725
transform 1 0 282164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire154_A
timestamp 1676037725
transform 1 0 277012 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire155_A
timestamp 1676037725
transform -1 0 272228 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire156_A
timestamp 1676037725
transform -1 0 267168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire157_A
timestamp 1676037725
transform -1 0 262108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire158_A
timestamp 1676037725
transform -1 0 257048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire159_A
timestamp 1676037725
transform 1 0 252448 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire160_A
timestamp 1676037725
transform -1 0 244628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire161_A
timestamp 1676037725
transform -1 0 240212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1676037725
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45
timestamp 1676037725
transform 1 0 5244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95
timestamp 1676037725
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1676037725
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123
timestamp 1676037725
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_129
timestamp 1676037725
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135
timestamp 1676037725
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151
timestamp 1676037725
transform 1 0 14996 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1676037725
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1676037725
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_185
timestamp 1676037725
transform 1 0 18124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_191
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_207
timestamp 1676037725
transform 1 0 20148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1676037725
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1676037725
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_235
timestamp 1676037725
transform 1 0 22724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_241
timestamp 1676037725
transform 1 0 23276 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_263
timestamp 1676037725
transform 1 0 25300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1676037725
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1676037725
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1676037725
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_297
timestamp 1676037725
transform 1 0 28428 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_303
timestamp 1676037725
transform 1 0 28980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1676037725
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_319
timestamp 1676037725
transform 1 0 30452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1676037725
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1676037725
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1676037725
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 1676037725
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_375
timestamp 1676037725
transform 1 0 35604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_387
timestamp 1676037725
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_403
timestamp 1676037725
transform 1 0 38180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1676037725
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1676037725
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_437
timestamp 1676037725
transform 1 0 41308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_459
timestamp 1676037725
transform 1 0 43332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_471
timestamp 1676037725
transform 1 0 44436 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1676037725
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_487
timestamp 1676037725
transform 1 0 45908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_499
timestamp 1676037725
transform 1 0 47012 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1676037725
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1676037725
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_521
timestamp 1676037725
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1676037725
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_543
timestamp 1676037725
transform 1 0 51060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_555
timestamp 1676037725
transform 1 0 52164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1676037725
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_561
timestamp 1676037725
transform 1 0 52716 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_571
timestamp 1676037725
transform 1 0 53636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_583
timestamp 1676037725
transform 1 0 54740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1676037725
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1676037725
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_605
timestamp 1676037725
transform 1 0 56764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1676037725
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_617
timestamp 1676037725
transform 1 0 57868 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_627
timestamp 1676037725
transform 1 0 58788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_639
timestamp 1676037725
transform 1 0 59892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_642
timestamp 1676037725
transform 1 0 60168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_645
timestamp 1676037725
transform 1 0 60444 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_655
timestamp 1676037725
transform 1 0 61364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_667
timestamp 1676037725
transform 1 0 62468 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_671
timestamp 1676037725
transform 1 0 62836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_673
timestamp 1676037725
transform 1 0 63020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_683
timestamp 1676037725
transform 1 0 63940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_689
timestamp 1676037725
transform 1 0 64492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1676037725
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_701
timestamp 1676037725
transform 1 0 65596 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_711
timestamp 1676037725
transform 1 0 66516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_723
timestamp 1676037725
transform 1 0 67620 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_727
timestamp 1676037725
transform 1 0 67988 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_729
timestamp 1676037725
transform 1 0 68172 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_739
timestamp 1676037725
transform 1 0 69092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_751
timestamp 1676037725
transform 1 0 70196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_755
timestamp 1676037725
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_757
timestamp 1676037725
transform 1 0 70748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_767
timestamp 1676037725
transform 1 0 71668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_773
timestamp 1676037725
transform 1 0 72220 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1676037725
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_785
timestamp 1676037725
transform 1 0 73324 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_795
timestamp 1676037725
transform 1 0 74244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_807
timestamp 1676037725
transform 1 0 75348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_810
timestamp 1676037725
transform 1 0 75624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_813
timestamp 1676037725
transform 1 0 75900 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_823
timestamp 1676037725
transform 1 0 76820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_835
timestamp 1676037725
transform 1 0 77924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_839
timestamp 1676037725
transform 1 0 78292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_841
timestamp 1676037725
transform 1 0 78476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_851
timestamp 1676037725
transform 1 0 79396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_857
timestamp 1676037725
transform 1 0 79948 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1676037725
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_869
timestamp 1676037725
transform 1 0 81052 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_879
timestamp 1676037725
transform 1 0 81972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_891
timestamp 1676037725
transform 1 0 83076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_895
timestamp 1676037725
transform 1 0 83444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_897
timestamp 1676037725
transform 1 0 83628 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_907
timestamp 1676037725
transform 1 0 84548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_919
timestamp 1676037725
transform 1 0 85652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_923
timestamp 1676037725
transform 1 0 86020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_925
timestamp 1676037725
transform 1 0 86204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_935
timestamp 1676037725
transform 1 0 87124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_941
timestamp 1676037725
transform 1 0 87676 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1676037725
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_953
timestamp 1676037725
transform 1 0 88780 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_963
timestamp 1676037725
transform 1 0 89700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_975
timestamp 1676037725
transform 1 0 90804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_978
timestamp 1676037725
transform 1 0 91080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_981
timestamp 1676037725
transform 1 0 91356 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_991
timestamp 1676037725
transform 1 0 92276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1003
timestamp 1676037725
transform 1 0 93380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1007
timestamp 1676037725
transform 1 0 93748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1009
timestamp 1676037725
transform 1 0 93932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1019
timestamp 1676037725
transform 1 0 94852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1025
timestamp 1676037725
transform 1 0 95404 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1676037725
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1037
timestamp 1676037725
transform 1 0 96508 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1047
timestamp 1676037725
transform 1 0 97428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1059
timestamp 1676037725
transform 1 0 98532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1063
timestamp 1676037725
transform 1 0 98900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1065
timestamp 1676037725
transform 1 0 99084 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1075
timestamp 1676037725
transform 1 0 100004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1087
timestamp 1676037725
transform 1 0 101108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1091
timestamp 1676037725
transform 1 0 101476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1093
timestamp 1676037725
transform 1 0 101660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1103
timestamp 1676037725
transform 1 0 102580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1109
timestamp 1676037725
transform 1 0 103132 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1676037725
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1121
timestamp 1676037725
transform 1 0 104236 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1131
timestamp 1676037725
transform 1 0 105156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1143
timestamp 1676037725
transform 1 0 106260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1146
timestamp 1676037725
transform 1 0 106536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1149
timestamp 1676037725
transform 1 0 106812 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1159
timestamp 1676037725
transform 1 0 107732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1171
timestamp 1676037725
transform 1 0 108836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1175
timestamp 1676037725
transform 1 0 109204 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1177
timestamp 1676037725
transform 1 0 109388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1187
timestamp 1676037725
transform 1 0 110308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1193
timestamp 1676037725
transform 1 0 110860 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1201
timestamp 1676037725
transform 1 0 111596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1205
timestamp 1676037725
transform 1 0 111964 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1215
timestamp 1676037725
transform 1 0 112884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1227
timestamp 1676037725
transform 1 0 113988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1231
timestamp 1676037725
transform 1 0 114356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1233
timestamp 1676037725
transform 1 0 114540 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1243
timestamp 1676037725
transform 1 0 115460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1255
timestamp 1676037725
transform 1 0 116564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1259
timestamp 1676037725
transform 1 0 116932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1261
timestamp 1676037725
transform 1 0 117116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1271
timestamp 1676037725
transform 1 0 118036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1277
timestamp 1676037725
transform 1 0 118588 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1285
timestamp 1676037725
transform 1 0 119324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1289
timestamp 1676037725
transform 1 0 119692 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1299
timestamp 1676037725
transform 1 0 120612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1311
timestamp 1676037725
transform 1 0 121716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1314
timestamp 1676037725
transform 1 0 121992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1317
timestamp 1676037725
transform 1 0 122268 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1327
timestamp 1676037725
transform 1 0 123188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1339
timestamp 1676037725
transform 1 0 124292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1343
timestamp 1676037725
transform 1 0 124660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1345
timestamp 1676037725
transform 1 0 124844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1355
timestamp 1676037725
transform 1 0 125764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1361
timestamp 1676037725
transform 1 0 126316 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1369
timestamp 1676037725
transform 1 0 127052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1373
timestamp 1676037725
transform 1 0 127420 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1383
timestamp 1676037725
transform 1 0 128340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1395
timestamp 1676037725
transform 1 0 129444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1399
timestamp 1676037725
transform 1 0 129812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1401
timestamp 1676037725
transform 1 0 129996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1407
timestamp 1676037725
transform 1 0 130548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1411
timestamp 1676037725
transform 1 0 130916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1417
timestamp 1676037725
transform 1 0 131468 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1425
timestamp 1676037725
transform 1 0 132204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1429
timestamp 1676037725
transform 1 0 132572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1439
timestamp 1676037725
transform 1 0 133492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1445
timestamp 1676037725
transform 1 0 134044 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1453
timestamp 1676037725
transform 1 0 134780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1457
timestamp 1676037725
transform 1 0 135148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1463
timestamp 1676037725
transform 1 0 135700 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1467
timestamp 1676037725
transform 1 0 136068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1473
timestamp 1676037725
transform 1 0 136620 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1481
timestamp 1676037725
transform 1 0 137356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1485
timestamp 1676037725
transform 1 0 137724 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1495
timestamp 1676037725
transform 1 0 138644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1507
timestamp 1676037725
transform 1 0 139748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1511
timestamp 1676037725
transform 1 0 140116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1513
timestamp 1676037725
transform 1 0 140300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1523
timestamp 1676037725
transform 1 0 141220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1529
timestamp 1676037725
transform 1 0 141772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1537
timestamp 1676037725
transform 1 0 142508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1541
timestamp 1676037725
transform 1 0 142876 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1551
timestamp 1676037725
transform 1 0 143796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1563
timestamp 1676037725
transform 1 0 144900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1567
timestamp 1676037725
transform 1 0 145268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1569
timestamp 1676037725
transform 1 0 145452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1579
timestamp 1676037725
transform 1 0 146372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1585
timestamp 1676037725
transform 1 0 146924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1593
timestamp 1676037725
transform 1 0 147660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1597
timestamp 1676037725
transform 1 0 148028 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1607
timestamp 1676037725
transform 1 0 148948 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1619
timestamp 1676037725
transform 1 0 150052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1623
timestamp 1676037725
transform 1 0 150420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1625
timestamp 1676037725
transform 1 0 150604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1635
timestamp 1676037725
transform 1 0 151524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1641
timestamp 1676037725
transform 1 0 152076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1649
timestamp 1676037725
transform 1 0 152812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1653
timestamp 1676037725
transform 1 0 153180 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1663
timestamp 1676037725
transform 1 0 154100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1675
timestamp 1676037725
transform 1 0 155204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1679
timestamp 1676037725
transform 1 0 155572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1681
timestamp 1676037725
transform 1 0 155756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1691
timestamp 1676037725
transform 1 0 156676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1697
timestamp 1676037725
transform 1 0 157228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1705
timestamp 1676037725
transform 1 0 157964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1709
timestamp 1676037725
transform 1 0 158332 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1719
timestamp 1676037725
transform 1 0 159252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1731
timestamp 1676037725
transform 1 0 160356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1735
timestamp 1676037725
transform 1 0 160724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1737
timestamp 1676037725
transform 1 0 160908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1747
timestamp 1676037725
transform 1 0 161828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1753
timestamp 1676037725
transform 1 0 162380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1761
timestamp 1676037725
transform 1 0 163116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1765
timestamp 1676037725
transform 1 0 163484 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1775
timestamp 1676037725
transform 1 0 164404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1787
timestamp 1676037725
transform 1 0 165508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1791
timestamp 1676037725
transform 1 0 165876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1793
timestamp 1676037725
transform 1 0 166060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1803
timestamp 1676037725
transform 1 0 166980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1809
timestamp 1676037725
transform 1 0 167532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1817
timestamp 1676037725
transform 1 0 168268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1821
timestamp 1676037725
transform 1 0 168636 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1831
timestamp 1676037725
transform 1 0 169556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1843
timestamp 1676037725
transform 1 0 170660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1847
timestamp 1676037725
transform 1 0 171028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1849
timestamp 1676037725
transform 1 0 171212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1859
timestamp 1676037725
transform 1 0 172132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1865
timestamp 1676037725
transform 1 0 172684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1873
timestamp 1676037725
transform 1 0 173420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1877
timestamp 1676037725
transform 1 0 173788 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1887
timestamp 1676037725
transform 1 0 174708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1899
timestamp 1676037725
transform 1 0 175812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1903
timestamp 1676037725
transform 1 0 176180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1905
timestamp 1676037725
transform 1 0 176364 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1915
timestamp 1676037725
transform 1 0 177284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1921
timestamp 1676037725
transform 1 0 177836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1929
timestamp 1676037725
transform 1 0 178572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1933
timestamp 1676037725
transform 1 0 178940 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1943
timestamp 1676037725
transform 1 0 179860 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1955
timestamp 1676037725
transform 1 0 180964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1959
timestamp 1676037725
transform 1 0 181332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1961
timestamp 1676037725
transform 1 0 181516 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1971
timestamp 1676037725
transform 1 0 182436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1977
timestamp 1676037725
transform 1 0 182988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1985
timestamp 1676037725
transform 1 0 183724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1989
timestamp 1676037725
transform 1 0 184092 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1999
timestamp 1676037725
transform 1 0 185012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2011
timestamp 1676037725
transform 1 0 186116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2015
timestamp 1676037725
transform 1 0 186484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2017
timestamp 1676037725
transform 1 0 186668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2027
timestamp 1676037725
transform 1 0 187588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2033
timestamp 1676037725
transform 1 0 188140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2041
timestamp 1676037725
transform 1 0 188876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2045
timestamp 1676037725
transform 1 0 189244 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2055
timestamp 1676037725
transform 1 0 190164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2067
timestamp 1676037725
transform 1 0 191268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2071
timestamp 1676037725
transform 1 0 191636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2073
timestamp 1676037725
transform 1 0 191820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2083
timestamp 1676037725
transform 1 0 192740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2089
timestamp 1676037725
transform 1 0 193292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2097
timestamp 1676037725
transform 1 0 194028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2101
timestamp 1676037725
transform 1 0 194396 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2111
timestamp 1676037725
transform 1 0 195316 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2123
timestamp 1676037725
transform 1 0 196420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2127
timestamp 1676037725
transform 1 0 196788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2129
timestamp 1676037725
transform 1 0 196972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2139
timestamp 1676037725
transform 1 0 197892 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2145
timestamp 1676037725
transform 1 0 198444 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2153
timestamp 1676037725
transform 1 0 199180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2157
timestamp 1676037725
transform 1 0 199548 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2167
timestamp 1676037725
transform 1 0 200468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2179
timestamp 1676037725
transform 1 0 201572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2183
timestamp 1676037725
transform 1 0 201940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2185
timestamp 1676037725
transform 1 0 202124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2195
timestamp 1676037725
transform 1 0 203044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2201
timestamp 1676037725
transform 1 0 203596 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2209
timestamp 1676037725
transform 1 0 204332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2213
timestamp 1676037725
transform 1 0 204700 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2223
timestamp 1676037725
transform 1 0 205620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2235
timestamp 1676037725
transform 1 0 206724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2239
timestamp 1676037725
transform 1 0 207092 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2241
timestamp 1676037725
transform 1 0 207276 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2251
timestamp 1676037725
transform 1 0 208196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2257
timestamp 1676037725
transform 1 0 208748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2265
timestamp 1676037725
transform 1 0 209484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2269
timestamp 1676037725
transform 1 0 209852 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2279
timestamp 1676037725
transform 1 0 210772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2291
timestamp 1676037725
transform 1 0 211876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2295
timestamp 1676037725
transform 1 0 212244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2297
timestamp 1676037725
transform 1 0 212428 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2307
timestamp 1676037725
transform 1 0 213348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2313
timestamp 1676037725
transform 1 0 213900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2321
timestamp 1676037725
transform 1 0 214636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2325
timestamp 1676037725
transform 1 0 215004 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2335
timestamp 1676037725
transform 1 0 215924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2347
timestamp 1676037725
transform 1 0 217028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2351
timestamp 1676037725
transform 1 0 217396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2353
timestamp 1676037725
transform 1 0 217580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2363
timestamp 1676037725
transform 1 0 218500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2369
timestamp 1676037725
transform 1 0 219052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2377
timestamp 1676037725
transform 1 0 219788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2381
timestamp 1676037725
transform 1 0 220156 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2391
timestamp 1676037725
transform 1 0 221076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2403
timestamp 1676037725
transform 1 0 222180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2407
timestamp 1676037725
transform 1 0 222548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2409
timestamp 1676037725
transform 1 0 222732 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2419
timestamp 1676037725
transform 1 0 223652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2425
timestamp 1676037725
transform 1 0 224204 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2433
timestamp 1676037725
transform 1 0 224940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2437
timestamp 1676037725
transform 1 0 225308 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2447
timestamp 1676037725
transform 1 0 226228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2459
timestamp 1676037725
transform 1 0 227332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2463
timestamp 1676037725
transform 1 0 227700 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2465
timestamp 1676037725
transform 1 0 227884 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2475
timestamp 1676037725
transform 1 0 228804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2481
timestamp 1676037725
transform 1 0 229356 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2489
timestamp 1676037725
transform 1 0 230092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2493
timestamp 1676037725
transform 1 0 230460 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2503
timestamp 1676037725
transform 1 0 231380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2509
timestamp 1676037725
transform 1 0 231932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2517
timestamp 1676037725
transform 1 0 232668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2521
timestamp 1676037725
transform 1 0 233036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2531
timestamp 1676037725
transform 1 0 233956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2537
timestamp 1676037725
transform 1 0 234508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2545
timestamp 1676037725
transform 1 0 235244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2549
timestamp 1676037725
transform 1 0 235612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2559
timestamp 1676037725
transform 1 0 236532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2565
timestamp 1676037725
transform 1 0 237084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2573
timestamp 1676037725
transform 1 0 237820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2577
timestamp 1676037725
transform 1 0 238188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2587
timestamp 1676037725
transform 1 0 239108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2593
timestamp 1676037725
transform 1 0 239660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2601
timestamp 1676037725
transform 1 0 240396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2605
timestamp 1676037725
transform 1 0 240764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2615
timestamp 1676037725
transform 1 0 241684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2621
timestamp 1676037725
transform 1 0 242236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2629
timestamp 1676037725
transform 1 0 242972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2633
timestamp 1676037725
transform 1 0 243340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2643
timestamp 1676037725
transform 1 0 244260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2649
timestamp 1676037725
transform 1 0 244812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2657
timestamp 1676037725
transform 1 0 245548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2661
timestamp 1676037725
transform 1 0 245916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2671
timestamp 1676037725
transform 1 0 246836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2677
timestamp 1676037725
transform 1 0 247388 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2685
timestamp 1676037725
transform 1 0 248124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2689
timestamp 1676037725
transform 1 0 248492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2699
timestamp 1676037725
transform 1 0 249412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2705
timestamp 1676037725
transform 1 0 249964 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2713
timestamp 1676037725
transform 1 0 250700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2717
timestamp 1676037725
transform 1 0 251068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2727
timestamp 1676037725
transform 1 0 251988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2733
timestamp 1676037725
transform 1 0 252540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2741
timestamp 1676037725
transform 1 0 253276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2745
timestamp 1676037725
transform 1 0 253644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2755
timestamp 1676037725
transform 1 0 254564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2761
timestamp 1676037725
transform 1 0 255116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2769
timestamp 1676037725
transform 1 0 255852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2773
timestamp 1676037725
transform 1 0 256220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2783
timestamp 1676037725
transform 1 0 257140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2789
timestamp 1676037725
transform 1 0 257692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2797
timestamp 1676037725
transform 1 0 258428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2801
timestamp 1676037725
transform 1 0 258796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2811
timestamp 1676037725
transform 1 0 259716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2817
timestamp 1676037725
transform 1 0 260268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2825
timestamp 1676037725
transform 1 0 261004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2829
timestamp 1676037725
transform 1 0 261372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2839
timestamp 1676037725
transform 1 0 262292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2845
timestamp 1676037725
transform 1 0 262844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2853
timestamp 1676037725
transform 1 0 263580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2857
timestamp 1676037725
transform 1 0 263948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2867
timestamp 1676037725
transform 1 0 264868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2873
timestamp 1676037725
transform 1 0 265420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2881
timestamp 1676037725
transform 1 0 266156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2885
timestamp 1676037725
transform 1 0 266524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2895
timestamp 1676037725
transform 1 0 267444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2901
timestamp 1676037725
transform 1 0 267996 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2909
timestamp 1676037725
transform 1 0 268732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2913
timestamp 1676037725
transform 1 0 269100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2923
timestamp 1676037725
transform 1 0 270020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2929
timestamp 1676037725
transform 1 0 270572 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2937
timestamp 1676037725
transform 1 0 271308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2941
timestamp 1676037725
transform 1 0 271676 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2951
timestamp 1676037725
transform 1 0 272596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2957
timestamp 1676037725
transform 1 0 273148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2965
timestamp 1676037725
transform 1 0 273884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2969
timestamp 1676037725
transform 1 0 274252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2979
timestamp 1676037725
transform 1 0 275172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2985
timestamp 1676037725
transform 1 0 275724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2993
timestamp 1676037725
transform 1 0 276460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2997
timestamp 1676037725
transform 1 0 276828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3007
timestamp 1676037725
transform 1 0 277748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3013
timestamp 1676037725
transform 1 0 278300 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3021
timestamp 1676037725
transform 1 0 279036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3025
timestamp 1676037725
transform 1 0 279404 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3035
timestamp 1676037725
transform 1 0 280324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3041
timestamp 1676037725
transform 1 0 280876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3049
timestamp 1676037725
transform 1 0 281612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3053
timestamp 1676037725
transform 1 0 281980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3063
timestamp 1676037725
transform 1 0 282900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3069
timestamp 1676037725
transform 1 0 283452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3077
timestamp 1676037725
transform 1 0 284188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3081
timestamp 1676037725
transform 1 0 284556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3091
timestamp 1676037725
transform 1 0 285476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3097
timestamp 1676037725
transform 1 0 286028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3105
timestamp 1676037725
transform 1 0 286764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3109
timestamp 1676037725
transform 1 0 287132 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3119
timestamp 1676037725
transform 1 0 288052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3125
timestamp 1676037725
transform 1 0 288604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3133
timestamp 1676037725
transform 1 0 289340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3137
timestamp 1676037725
transform 1 0 289708 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3147
timestamp 1676037725
transform 1 0 290628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3153
timestamp 1676037725
transform 1 0 291180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3161
timestamp 1676037725
transform 1 0 291916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3165
timestamp 1676037725
transform 1 0 292284 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3175
timestamp 1676037725
transform 1 0 293204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3181
timestamp 1676037725
transform 1 0 293756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3189
timestamp 1676037725
transform 1 0 294492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3193
timestamp 1676037725
transform 1 0 294860 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3203
timestamp 1676037725
transform 1 0 295780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3209
timestamp 1676037725
transform 1 0 296332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3217
timestamp 1676037725
transform 1 0 297068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3221
timestamp 1676037725
transform 1 0 297436 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3231
timestamp 1676037725
transform 1 0 298356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3237
timestamp 1676037725
transform 1 0 298908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3245
timestamp 1676037725
transform 1 0 299644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3249
timestamp 1676037725
transform 1 0 300012 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3259
timestamp 1676037725
transform 1 0 300932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3265
timestamp 1676037725
transform 1 0 301484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3273
timestamp 1676037725
transform 1 0 302220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3277
timestamp 1676037725
transform 1 0 302588 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3287
timestamp 1676037725
transform 1 0 303508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3293
timestamp 1676037725
transform 1 0 304060 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3301
timestamp 1676037725
transform 1 0 304796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3305
timestamp 1676037725
transform 1 0 305164 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3315
timestamp 1676037725
transform 1 0 306084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3321
timestamp 1676037725
transform 1 0 306636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3329
timestamp 1676037725
transform 1 0 307372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3333
timestamp 1676037725
transform 1 0 307740 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3343
timestamp 1676037725
transform 1 0 308660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3349
timestamp 1676037725
transform 1 0 309212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3357
timestamp 1676037725
transform 1 0 309948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3361
timestamp 1676037725
transform 1 0 310316 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3371
timestamp 1676037725
transform 1 0 311236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3377
timestamp 1676037725
transform 1 0 311788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3385
timestamp 1676037725
transform 1 0 312524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3389
timestamp 1676037725
transform 1 0 312892 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3399
timestamp 1676037725
transform 1 0 313812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3405
timestamp 1676037725
transform 1 0 314364 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3413
timestamp 1676037725
transform 1 0 315100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3417
timestamp 1676037725
transform 1 0 315468 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3427
timestamp 1676037725
transform 1 0 316388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3433
timestamp 1676037725
transform 1 0 316940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3441
timestamp 1676037725
transform 1 0 317676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3445
timestamp 1676037725
transform 1 0 318044 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3455
timestamp 1676037725
transform 1 0 318964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3461
timestamp 1676037725
transform 1 0 319516 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3469
timestamp 1676037725
transform 1 0 320252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3473
timestamp 1676037725
transform 1 0 320620 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3483
timestamp 1676037725
transform 1 0 321540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3489
timestamp 1676037725
transform 1 0 322092 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3497
timestamp 1676037725
transform 1 0 322828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3501
timestamp 1676037725
transform 1 0 323196 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3511
timestamp 1676037725
transform 1 0 324116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3517
timestamp 1676037725
transform 1 0 324668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3525
timestamp 1676037725
transform 1 0 325404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3529
timestamp 1676037725
transform 1 0 325772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3539
timestamp 1676037725
transform 1 0 326692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3545
timestamp 1676037725
transform 1 0 327244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3553
timestamp 1676037725
transform 1 0 327980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3557
timestamp 1676037725
transform 1 0 328348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3567
timestamp 1676037725
transform 1 0 329268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3573
timestamp 1676037725
transform 1 0 329820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3581
timestamp 1676037725
transform 1 0 330556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3585
timestamp 1676037725
transform 1 0 330924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3595
timestamp 1676037725
transform 1 0 331844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3601
timestamp 1676037725
transform 1 0 332396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3609
timestamp 1676037725
transform 1 0 333132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3613
timestamp 1676037725
transform 1 0 333500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3623
timestamp 1676037725
transform 1 0 334420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3629
timestamp 1676037725
transform 1 0 334972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3637
timestamp 1676037725
transform 1 0 335708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3641
timestamp 1676037725
transform 1 0 336076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3651
timestamp 1676037725
transform 1 0 336996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3657
timestamp 1676037725
transform 1 0 337548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3665
timestamp 1676037725
transform 1 0 338284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3669
timestamp 1676037725
transform 1 0 338652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3679
timestamp 1676037725
transform 1 0 339572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3685
timestamp 1676037725
transform 1 0 340124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3693
timestamp 1676037725
transform 1 0 340860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3697
timestamp 1676037725
transform 1 0 341228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3707
timestamp 1676037725
transform 1 0 342148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3713
timestamp 1676037725
transform 1 0 342700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3721
timestamp 1676037725
transform 1 0 343436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3725
timestamp 1676037725
transform 1 0 343804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3735
timestamp 1676037725
transform 1 0 344724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3741
timestamp 1676037725
transform 1 0 345276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3749
timestamp 1676037725
transform 1 0 346012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3753
timestamp 1676037725
transform 1 0 346380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3763
timestamp 1676037725
transform 1 0 347300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3769
timestamp 1676037725
transform 1 0 347852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3777
timestamp 1676037725
transform 1 0 348588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3781
timestamp 1676037725
transform 1 0 348956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3791
timestamp 1676037725
transform 1 0 349876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3797
timestamp 1676037725
transform 1 0 350428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3805
timestamp 1676037725
transform 1 0 351164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3809
timestamp 1676037725
transform 1 0 351532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3819
timestamp 1676037725
transform 1 0 352452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3825
timestamp 1676037725
transform 1 0 353004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3833
timestamp 1676037725
transform 1 0 353740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3837
timestamp 1676037725
transform 1 0 354108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3847
timestamp 1676037725
transform 1 0 355028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3853
timestamp 1676037725
transform 1 0 355580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3861
timestamp 1676037725
transform 1 0 356316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3865
timestamp 1676037725
transform 1 0 356684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3875
timestamp 1676037725
transform 1 0 357604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3881
timestamp 1676037725
transform 1 0 358156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3889
timestamp 1676037725
transform 1 0 358892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3893
timestamp 1676037725
transform 1 0 359260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3903
timestamp 1676037725
transform 1 0 360180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3909
timestamp 1676037725
transform 1 0 360732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3917
timestamp 1676037725
transform 1 0 361468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3921
timestamp 1676037725
transform 1 0 361836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3931
timestamp 1676037725
transform 1 0 362756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3937
timestamp 1676037725
transform 1 0 363308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3945
timestamp 1676037725
transform 1 0 364044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3949
timestamp 1676037725
transform 1 0 364412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3959
timestamp 1676037725
transform 1 0 365332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3965
timestamp 1676037725
transform 1 0 365884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3973
timestamp 1676037725
transform 1 0 366620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3977
timestamp 1676037725
transform 1 0 366988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3987
timestamp 1676037725
transform 1 0 367908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3993
timestamp 1676037725
transform 1 0 368460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4001
timestamp 1676037725
transform 1 0 369196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4005
timestamp 1676037725
transform 1 0 369564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4015
timestamp 1676037725
transform 1 0 370484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4021
timestamp 1676037725
transform 1 0 371036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4029
timestamp 1676037725
transform 1 0 371772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4033
timestamp 1676037725
transform 1 0 372140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4043
timestamp 1676037725
transform 1 0 373060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4049
timestamp 1676037725
transform 1 0 373612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4057
timestamp 1676037725
transform 1 0 374348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4061
timestamp 1676037725
transform 1 0 374716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4071
timestamp 1676037725
transform 1 0 375636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4077
timestamp 1676037725
transform 1 0 376188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4085
timestamp 1676037725
transform 1 0 376924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4089
timestamp 1676037725
transform 1 0 377292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4099
timestamp 1676037725
transform 1 0 378212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4105
timestamp 1676037725
transform 1 0 378764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4113
timestamp 1676037725
transform 1 0 379500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4117
timestamp 1676037725
transform 1 0 379868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4127
timestamp 1676037725
transform 1 0 380788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4133
timestamp 1676037725
transform 1 0 381340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4141
timestamp 1676037725
transform 1 0 382076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4145
timestamp 1676037725
transform 1 0 382444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4155
timestamp 1676037725
transform 1 0 383364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4161
timestamp 1676037725
transform 1 0 383916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4169
timestamp 1676037725
transform 1 0 384652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4173
timestamp 1676037725
transform 1 0 385020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4183
timestamp 1676037725
transform 1 0 385940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4189
timestamp 1676037725
transform 1 0 386492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4197
timestamp 1676037725
transform 1 0 387228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4201
timestamp 1676037725
transform 1 0 387596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4211
timestamp 1676037725
transform 1 0 388516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4217
timestamp 1676037725
transform 1 0 389068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4225
timestamp 1676037725
transform 1 0 389804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4229
timestamp 1676037725
transform 1 0 390172 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4239
timestamp 1676037725
transform 1 0 391092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4245
timestamp 1676037725
transform 1 0 391644 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4253
timestamp 1676037725
transform 1 0 392380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4257
timestamp 1676037725
transform 1 0 392748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4267
timestamp 1676037725
transform 1 0 393668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4273
timestamp 1676037725
transform 1 0 394220 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4281
timestamp 1676037725
transform 1 0 394956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4285
timestamp 1676037725
transform 1 0 395324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4295
timestamp 1676037725
transform 1 0 396244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4301
timestamp 1676037725
transform 1 0 396796 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4309
timestamp 1676037725
transform 1 0 397532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4313
timestamp 1676037725
transform 1 0 397900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4323
timestamp 1676037725
transform 1 0 398820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4329
timestamp 1676037725
transform 1 0 399372 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4337
timestamp 1676037725
transform 1 0 400108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4341
timestamp 1676037725
transform 1 0 400476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4351
timestamp 1676037725
transform 1 0 401396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4357
timestamp 1676037725
transform 1 0 401948 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4365
timestamp 1676037725
transform 1 0 402684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4369
timestamp 1676037725
transform 1 0 403052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4379
timestamp 1676037725
transform 1 0 403972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4385
timestamp 1676037725
transform 1 0 404524 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4393
timestamp 1676037725
transform 1 0 405260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4397
timestamp 1676037725
transform 1 0 405628 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4407
timestamp 1676037725
transform 1 0 406548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4413
timestamp 1676037725
transform 1 0 407100 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4421
timestamp 1676037725
transform 1 0 407836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4425
timestamp 1676037725
transform 1 0 408204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4435
timestamp 1676037725
transform 1 0 409124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4441
timestamp 1676037725
transform 1 0 409676 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4449
timestamp 1676037725
transform 1 0 410412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4453
timestamp 1676037725
transform 1 0 410780 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4463
timestamp 1676037725
transform 1 0 411700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4469
timestamp 1676037725
transform 1 0 412252 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4477
timestamp 1676037725
transform 1 0 412988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4481
timestamp 1676037725
transform 1 0 413356 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4491
timestamp 1676037725
transform 1 0 414276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4497
timestamp 1676037725
transform 1 0 414828 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4505
timestamp 1676037725
transform 1 0 415564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4509
timestamp 1676037725
transform 1 0 415932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4519
timestamp 1676037725
transform 1 0 416852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4525
timestamp 1676037725
transform 1 0 417404 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4533
timestamp 1676037725
transform 1 0 418140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4537
timestamp 1676037725
transform 1 0 418508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4547
timestamp 1676037725
transform 1 0 419428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4553
timestamp 1676037725
transform 1 0 419980 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4561
timestamp 1676037725
transform 1 0 420716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4565
timestamp 1676037725
transform 1 0 421084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4575
timestamp 1676037725
transform 1 0 422004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4581
timestamp 1676037725
transform 1 0 422556 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4589
timestamp 1676037725
transform 1 0 423292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4593
timestamp 1676037725
transform 1 0 423660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4603
timestamp 1676037725
transform 1 0 424580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4609
timestamp 1676037725
transform 1 0 425132 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4617
timestamp 1676037725
transform 1 0 425868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4621
timestamp 1676037725
transform 1 0 426236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4631
timestamp 1676037725
transform 1 0 427156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4637
timestamp 1676037725
transform 1 0 427708 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4645
timestamp 1676037725
transform 1 0 428444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4649
timestamp 1676037725
transform 1 0 428812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4659
timestamp 1676037725
transform 1 0 429732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4665
timestamp 1676037725
transform 1 0 430284 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4673
timestamp 1676037725
transform 1 0 431020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4677
timestamp 1676037725
transform 1 0 431388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4687
timestamp 1676037725
transform 1 0 432308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4693
timestamp 1676037725
transform 1 0 432860 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4701
timestamp 1676037725
transform 1 0 433596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4705
timestamp 1676037725
transform 1 0 433964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4715
timestamp 1676037725
transform 1 0 434884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4721
timestamp 1676037725
transform 1 0 435436 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4729
timestamp 1676037725
transform 1 0 436172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4733
timestamp 1676037725
transform 1 0 436540 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4743
timestamp 1676037725
transform 1 0 437460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4749
timestamp 1676037725
transform 1 0 438012 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4757
timestamp 1676037725
transform 1 0 438748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4761
timestamp 1676037725
transform 1 0 439116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4771
timestamp 1676037725
transform 1 0 440036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4777
timestamp 1676037725
transform 1 0 440588 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4785
timestamp 1676037725
transform 1 0 441324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4789
timestamp 1676037725
transform 1 0 441692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4799
timestamp 1676037725
transform 1 0 442612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4805
timestamp 1676037725
transform 1 0 443164 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4813
timestamp 1676037725
transform 1 0 443900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4817
timestamp 1676037725
transform 1 0 444268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4827
timestamp 1676037725
transform 1 0 445188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4833
timestamp 1676037725
transform 1 0 445740 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4841
timestamp 1676037725
transform 1 0 446476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4845
timestamp 1676037725
transform 1 0 446844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4855
timestamp 1676037725
transform 1 0 447764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4861
timestamp 1676037725
transform 1 0 448316 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4869
timestamp 1676037725
transform 1 0 449052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4873
timestamp 1676037725
transform 1 0 449420 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4883
timestamp 1676037725
transform 1 0 450340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4889
timestamp 1676037725
transform 1 0 450892 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4897
timestamp 1676037725
transform 1 0 451628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4901
timestamp 1676037725
transform 1 0 451996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4911
timestamp 1676037725
transform 1 0 452916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4917
timestamp 1676037725
transform 1 0 453468 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4925
timestamp 1676037725
transform 1 0 454204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4929
timestamp 1676037725
transform 1 0 454572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4939
timestamp 1676037725
transform 1 0 455492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4945
timestamp 1676037725
transform 1 0 456044 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4953
timestamp 1676037725
transform 1 0 456780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4957
timestamp 1676037725
transform 1 0 457148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4967
timestamp 1676037725
transform 1 0 458068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4973
timestamp 1676037725
transform 1 0 458620 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4981
timestamp 1676037725
transform 1 0 459356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4985
timestamp 1676037725
transform 1 0 459724 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4995
timestamp 1676037725
transform 1 0 460644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5001
timestamp 1676037725
transform 1 0 461196 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5009
timestamp 1676037725
transform 1 0 461932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5013
timestamp 1676037725
transform 1 0 462300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5023
timestamp 1676037725
transform 1 0 463220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5029
timestamp 1676037725
transform 1 0 463772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5037
timestamp 1676037725
transform 1 0 464508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5041
timestamp 1676037725
transform 1 0 464876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5051
timestamp 1676037725
transform 1 0 465796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5057
timestamp 1676037725
transform 1 0 466348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5065
timestamp 1676037725
transform 1 0 467084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5069
timestamp 1676037725
transform 1 0 467452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5079
timestamp 1676037725
transform 1 0 468372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5085
timestamp 1676037725
transform 1 0 468924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5093
timestamp 1676037725
transform 1 0 469660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5097
timestamp 1676037725
transform 1 0 470028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5107
timestamp 1676037725
transform 1 0 470948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5113
timestamp 1676037725
transform 1 0 471500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5121
timestamp 1676037725
transform 1 0 472236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5125
timestamp 1676037725
transform 1 0 472604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5135
timestamp 1676037725
transform 1 0 473524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5141
timestamp 1676037725
transform 1 0 474076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5149
timestamp 1676037725
transform 1 0 474812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5153
timestamp 1676037725
transform 1 0 475180 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5163
timestamp 1676037725
transform 1 0 476100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5169
timestamp 1676037725
transform 1 0 476652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5177
timestamp 1676037725
transform 1 0 477388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5181
timestamp 1676037725
transform 1 0 477756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5191
timestamp 1676037725
transform 1 0 478676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5197
timestamp 1676037725
transform 1 0 479228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5205
timestamp 1676037725
transform 1 0 479964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5209
timestamp 1676037725
transform 1 0 480332 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5219
timestamp 1676037725
transform 1 0 481252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5225
timestamp 1676037725
transform 1 0 481804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5233
timestamp 1676037725
transform 1 0 482540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5237
timestamp 1676037725
transform 1 0 482908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5247
timestamp 1676037725
transform 1 0 483828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5253
timestamp 1676037725
transform 1 0 484380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5261
timestamp 1676037725
transform 1 0 485116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5265
timestamp 1676037725
transform 1 0 485484 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5275
timestamp 1676037725
transform 1 0 486404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5287
timestamp 1676037725
transform 1 0 487508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5291
timestamp 1676037725
transform 1 0 487876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5293
timestamp 1676037725
transform 1 0 488060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5303
timestamp 1676037725
transform 1 0 488980 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5315
timestamp 1676037725
transform 1 0 490084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5319
timestamp 1676037725
transform 1 0 490452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5321
timestamp 1676037725
transform 1 0 490636 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5331
timestamp 1676037725
transform 1 0 491556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5343
timestamp 1676037725
transform 1 0 492660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5347
timestamp 1676037725
transform 1 0 493028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5349
timestamp 1676037725
transform 1 0 493212 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5359
timestamp 1676037725
transform 1 0 494132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5371
timestamp 1676037725
transform 1 0 495236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5375
timestamp 1676037725
transform 1 0 495604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5377
timestamp 1676037725
transform 1 0 495788 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5387
timestamp 1676037725
transform 1 0 496708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5399
timestamp 1676037725
transform 1 0 497812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5403
timestamp 1676037725
transform 1 0 498180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5405
timestamp 1676037725
transform 1 0 498364 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5415
timestamp 1676037725
transform 1 0 499284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5427
timestamp 1676037725
transform 1 0 500388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5431
timestamp 1676037725
transform 1 0 500756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5433
timestamp 1676037725
transform 1 0 500940 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5443
timestamp 1676037725
transform 1 0 501860 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5455
timestamp 1676037725
transform 1 0 502964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5459
timestamp 1676037725
transform 1 0 503332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5461
timestamp 1676037725
transform 1 0 503516 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5471
timestamp 1676037725
transform 1 0 504436 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5483
timestamp 1676037725
transform 1 0 505540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5487
timestamp 1676037725
transform 1 0 505908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5489
timestamp 1676037725
transform 1 0 506092 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5499
timestamp 1676037725
transform 1 0 507012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5511
timestamp 1676037725
transform 1 0 508116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5515
timestamp 1676037725
transform 1 0 508484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5517
timestamp 1676037725
transform 1 0 508668 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5527
timestamp 1676037725
transform 1 0 509588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5539
timestamp 1676037725
transform 1 0 510692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5543
timestamp 1676037725
transform 1 0 511060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5545
timestamp 1676037725
transform 1 0 511244 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5555
timestamp 1676037725
transform 1 0 512164 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5567
timestamp 1676037725
transform 1 0 513268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5571
timestamp 1676037725
transform 1 0 513636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5573
timestamp 1676037725
transform 1 0 513820 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5583
timestamp 1676037725
transform 1 0 514740 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5595
timestamp 1676037725
transform 1 0 515844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5599
timestamp 1676037725
transform 1 0 516212 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5601
timestamp 1676037725
transform 1 0 516396 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5613
timestamp 1676037725
transform 1 0 517500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5625
timestamp 1676037725
transform 1 0 518604 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5629
timestamp 1676037725
transform 1 0 518972 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5641
timestamp 1676037725
transform 1 0 520076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5653
timestamp 1676037725
transform 1 0 521180 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5657
timestamp 1676037725
transform 1 0 521548 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5669
timestamp 1676037725
transform 1 0 522652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5681
timestamp 1676037725
transform 1 0 523756 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5685
timestamp 1676037725
transform 1 0 524124 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5697
timestamp 1676037725
transform 1 0 525228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5709
timestamp 1676037725
transform 1 0 526332 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5713
timestamp 1676037725
transform 1 0 526700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5725
timestamp 1676037725
transform 1 0 527804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7
timestamp 1676037725
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1676037725
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_45
timestamp 1676037725
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1676037725
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_61
timestamp 1676037725
transform 1 0 6716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_73
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1676037725
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_89
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1676037725
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 1676037725
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_201
timestamp 1676037725
transform 1 0 19596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_213
timestamp 1676037725
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1676037725
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_257
timestamp 1676037725
transform 1 0 24748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1676037725
transform 1 0 25852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1676037725
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_313
timestamp 1676037725
transform 1 0 29900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_325
timestamp 1676037725
transform 1 0 31004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1676037725
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_369
timestamp 1676037725
transform 1 0 35052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_381
timestamp 1676037725
transform 1 0 36156 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_389
timestamp 1676037725
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_397
timestamp 1676037725
transform 1 0 37628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_409
timestamp 1676037725
transform 1 0 38732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_421
timestamp 1676037725
transform 1 0 39836 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_427
timestamp 1676037725
transform 1 0 40388 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_439
timestamp 1676037725
transform 1 0 41492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_455
timestamp 1676037725
transform 1 0 42964 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_467
timestamp 1676037725
transform 1 0 44068 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_479
timestamp 1676037725
transform 1 0 45172 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_483
timestamp 1676037725
transform 1 0 45540 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_495
timestamp 1676037725
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_529
timestamp 1676037725
transform 1 0 49772 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_539
timestamp 1676037725
transform 1 0 50692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_551
timestamp 1676037725
transform 1 0 51796 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1676037725
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_567
timestamp 1676037725
transform 1 0 53268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_579
timestamp 1676037725
transform 1 0 54372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_591
timestamp 1676037725
transform 1 0 55476 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_595
timestamp 1676037725
transform 1 0 55844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_607
timestamp 1676037725
transform 1 0 56948 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1676037725
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_623
timestamp 1676037725
transform 1 0 58420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_635
timestamp 1676037725
transform 1 0 59524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_647
timestamp 1676037725
transform 1 0 60628 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_651
timestamp 1676037725
transform 1 0 60996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_663
timestamp 1676037725
transform 1 0 62100 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1676037725
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1676037725
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1676037725
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_697
timestamp 1676037725
transform 1 0 65228 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_707
timestamp 1676037725
transform 1 0 66148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_719
timestamp 1676037725
transform 1 0 67252 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1676037725
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1676037725
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_735
timestamp 1676037725
transform 1 0 68724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_747
timestamp 1676037725
transform 1 0 69828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_759
timestamp 1676037725
transform 1 0 70932 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_763
timestamp 1676037725
transform 1 0 71300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_775
timestamp 1676037725
transform 1 0 72404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1676037725
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_785
timestamp 1676037725
transform 1 0 73324 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_791
timestamp 1676037725
transform 1 0 73876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_803
timestamp 1676037725
transform 1 0 74980 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_815
timestamp 1676037725
transform 1 0 76084 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_819
timestamp 1676037725
transform 1 0 76452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_831
timestamp 1676037725
transform 1 0 77556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1676037725
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1676037725
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1676037725
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_865
timestamp 1676037725
transform 1 0 80684 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_875
timestamp 1676037725
transform 1 0 81604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_887
timestamp 1676037725
transform 1 0 82708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1676037725
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_897
timestamp 1676037725
transform 1 0 83628 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_903
timestamp 1676037725
transform 1 0 84180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_915
timestamp 1676037725
transform 1 0 85284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_927
timestamp 1676037725
transform 1 0 86388 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_931
timestamp 1676037725
transform 1 0 86756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_943
timestamp 1676037725
transform 1 0 87860 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1676037725
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_953
timestamp 1676037725
transform 1 0 88780 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_959
timestamp 1676037725
transform 1 0 89332 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_971
timestamp 1676037725
transform 1 0 90436 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_983
timestamp 1676037725
transform 1 0 91540 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_987
timestamp 1676037725
transform 1 0 91908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_999
timestamp 1676037725
transform 1 0 93012 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1676037725
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1676037725
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1676037725
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1033
timestamp 1676037725
transform 1 0 96140 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1043
timestamp 1676037725
transform 1 0 97060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1055
timestamp 1676037725
transform 1 0 98164 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1676037725
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1065
timestamp 1676037725
transform 1 0 99084 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1071
timestamp 1676037725
transform 1 0 99636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1083
timestamp 1676037725
transform 1 0 100740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1095
timestamp 1676037725
transform 1 0 101844 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1099
timestamp 1676037725
transform 1 0 102212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1111
timestamp 1676037725
transform 1 0 103316 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1676037725
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1121
timestamp 1676037725
transform 1 0 104236 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1127
timestamp 1676037725
transform 1 0 104788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1139
timestamp 1676037725
transform 1 0 105892 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1151
timestamp 1676037725
transform 1 0 106996 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1155
timestamp 1676037725
transform 1 0 107364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1167
timestamp 1676037725
transform 1 0 108468 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1676037725
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1177
timestamp 1676037725
transform 1 0 109388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1189
timestamp 1676037725
transform 1 0 110492 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1201
timestamp 1676037725
transform 1 0 111596 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1211
timestamp 1676037725
transform 1 0 112516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1223
timestamp 1676037725
transform 1 0 113620 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1676037725
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1233
timestamp 1676037725
transform 1 0 114540 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1239
timestamp 1676037725
transform 1 0 115092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1251
timestamp 1676037725
transform 1 0 116196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1263
timestamp 1676037725
transform 1 0 117300 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1267
timestamp 1676037725
transform 1 0 117668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1279
timestamp 1676037725
transform 1 0 118772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1287
timestamp 1676037725
transform 1 0 119508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1289
timestamp 1676037725
transform 1 0 119692 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1295
timestamp 1676037725
transform 1 0 120244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1307
timestamp 1676037725
transform 1 0 121348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1319
timestamp 1676037725
transform 1 0 122452 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1323
timestamp 1676037725
transform 1 0 122820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1335
timestamp 1676037725
transform 1 0 123924 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1343
timestamp 1676037725
transform 1 0 124660 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1345
timestamp 1676037725
transform 1 0 124844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1357
timestamp 1676037725
transform 1 0 125948 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1369
timestamp 1676037725
transform 1 0 127052 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1379
timestamp 1676037725
transform 1 0 127972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1391
timestamp 1676037725
transform 1 0 129076 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1399
timestamp 1676037725
transform 1 0 129812 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1401
timestamp 1676037725
transform 1 0 129996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1413
timestamp 1676037725
transform 1 0 131100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1425
timestamp 1676037725
transform 1 0 132204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1437
timestamp 1676037725
transform 1 0 133308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1449
timestamp 1676037725
transform 1 0 134412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1455
timestamp 1676037725
transform 1 0 134964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1457
timestamp 1676037725
transform 1 0 135148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1469
timestamp 1676037725
transform 1 0 136252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1481
timestamp 1676037725
transform 1 0 137356 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1489
timestamp 1676037725
transform 1 0 138092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1501
timestamp 1676037725
transform 1 0 139196 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1509
timestamp 1676037725
transform 1 0 139932 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1513
timestamp 1676037725
transform 1 0 140300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1525
timestamp 1676037725
transform 1 0 141404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1537
timestamp 1676037725
transform 1 0 142508 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1545
timestamp 1676037725
transform 1 0 143244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1557
timestamp 1676037725
transform 1 0 144348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1565
timestamp 1676037725
transform 1 0 145084 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1569
timestamp 1676037725
transform 1 0 145452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1581
timestamp 1676037725
transform 1 0 146556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1593
timestamp 1676037725
transform 1 0 147660 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1601
timestamp 1676037725
transform 1 0 148396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1613
timestamp 1676037725
transform 1 0 149500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1621
timestamp 1676037725
transform 1 0 150236 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1625
timestamp 1676037725
transform 1 0 150604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1637
timestamp 1676037725
transform 1 0 151708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1649
timestamp 1676037725
transform 1 0 152812 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1657
timestamp 1676037725
transform 1 0 153548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1669
timestamp 1676037725
transform 1 0 154652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1677
timestamp 1676037725
transform 1 0 155388 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1681
timestamp 1676037725
transform 1 0 155756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1693
timestamp 1676037725
transform 1 0 156860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1705
timestamp 1676037725
transform 1 0 157964 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1713
timestamp 1676037725
transform 1 0 158700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1725
timestamp 1676037725
transform 1 0 159804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1733
timestamp 1676037725
transform 1 0 160540 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1737
timestamp 1676037725
transform 1 0 160908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1749
timestamp 1676037725
transform 1 0 162012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1761
timestamp 1676037725
transform 1 0 163116 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1769
timestamp 1676037725
transform 1 0 163852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1781
timestamp 1676037725
transform 1 0 164956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1789
timestamp 1676037725
transform 1 0 165692 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1793
timestamp 1676037725
transform 1 0 166060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1805
timestamp 1676037725
transform 1 0 167164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1817
timestamp 1676037725
transform 1 0 168268 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1825
timestamp 1676037725
transform 1 0 169004 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1837
timestamp 1676037725
transform 1 0 170108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1845
timestamp 1676037725
transform 1 0 170844 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1849
timestamp 1676037725
transform 1 0 171212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1861
timestamp 1676037725
transform 1 0 172316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1873
timestamp 1676037725
transform 1 0 173420 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1881
timestamp 1676037725
transform 1 0 174156 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1893
timestamp 1676037725
transform 1 0 175260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1901
timestamp 1676037725
transform 1 0 175996 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1905
timestamp 1676037725
transform 1 0 176364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1917
timestamp 1676037725
transform 1 0 177468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1929
timestamp 1676037725
transform 1 0 178572 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1937
timestamp 1676037725
transform 1 0 179308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1949
timestamp 1676037725
transform 1 0 180412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1957
timestamp 1676037725
transform 1 0 181148 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1961
timestamp 1676037725
transform 1 0 181516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1973
timestamp 1676037725
transform 1 0 182620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1985
timestamp 1676037725
transform 1 0 183724 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1993
timestamp 1676037725
transform 1 0 184460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2005
timestamp 1676037725
transform 1 0 185564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_2013
timestamp 1676037725
transform 1 0 186300 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2017
timestamp 1676037725
transform 1 0 186668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2029
timestamp 1676037725
transform 1 0 187772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2041
timestamp 1676037725
transform 1 0 188876 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2049
timestamp 1676037725
transform 1 0 189612 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2061
timestamp 1676037725
transform 1 0 190716 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_2069
timestamp 1676037725
transform 1 0 191452 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2073
timestamp 1676037725
transform 1 0 191820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2085
timestamp 1676037725
transform 1 0 192924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2097
timestamp 1676037725
transform 1 0 194028 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2105
timestamp 1676037725
transform 1 0 194764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2117
timestamp 1676037725
transform 1 0 195868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_2125
timestamp 1676037725
transform 1 0 196604 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2129
timestamp 1676037725
transform 1 0 196972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2141
timestamp 1676037725
transform 1 0 198076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2153
timestamp 1676037725
transform 1 0 199180 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2163
timestamp 1676037725
transform 1 0 200100 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2175
timestamp 1676037725
transform 1 0 201204 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2183
timestamp 1676037725
transform 1 0 201940 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2185
timestamp 1676037725
transform 1 0 202124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2197
timestamp 1676037725
transform 1 0 203228 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2209
timestamp 1676037725
transform 1 0 204332 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2219
timestamp 1676037725
transform 1 0 205252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2231
timestamp 1676037725
transform 1 0 206356 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2239
timestamp 1676037725
transform 1 0 207092 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2241
timestamp 1676037725
transform 1 0 207276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2253
timestamp 1676037725
transform 1 0 208380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2265
timestamp 1676037725
transform 1 0 209484 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2275
timestamp 1676037725
transform 1 0 210404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2287
timestamp 1676037725
transform 1 0 211508 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2295
timestamp 1676037725
transform 1 0 212244 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2297
timestamp 1676037725
transform 1 0 212428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2309
timestamp 1676037725
transform 1 0 213532 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2321
timestamp 1676037725
transform 1 0 214636 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2331
timestamp 1676037725
transform 1 0 215556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2343
timestamp 1676037725
transform 1 0 216660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2351
timestamp 1676037725
transform 1 0 217396 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2353
timestamp 1676037725
transform 1 0 217580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2365
timestamp 1676037725
transform 1 0 218684 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2377
timestamp 1676037725
transform 1 0 219788 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2387
timestamp 1676037725
transform 1 0 220708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2399
timestamp 1676037725
transform 1 0 221812 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2407
timestamp 1676037725
transform 1 0 222548 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2409
timestamp 1676037725
transform 1 0 222732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2421
timestamp 1676037725
transform 1 0 223836 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2433
timestamp 1676037725
transform 1 0 224940 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2443
timestamp 1676037725
transform 1 0 225860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_2455
timestamp 1676037725
transform 1 0 226964 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2463
timestamp 1676037725
transform 1 0 227700 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2465
timestamp 1676037725
transform 1 0 227884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2477
timestamp 1676037725
transform 1 0 228988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2489
timestamp 1676037725
transform 1 0 230092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2501
timestamp 1676037725
transform 1 0 231196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2513
timestamp 1676037725
transform 1 0 232300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2519
timestamp 1676037725
transform 1 0 232852 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2521
timestamp 1676037725
transform 1 0 233036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2533
timestamp 1676037725
transform 1 0 234140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2545
timestamp 1676037725
transform 1 0 235244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2557
timestamp 1676037725
transform 1 0 236348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2569
timestamp 1676037725
transform 1 0 237452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2575
timestamp 1676037725
transform 1 0 238004 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2577
timestamp 1676037725
transform 1 0 238188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2589
timestamp 1676037725
transform 1 0 239292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2601
timestamp 1676037725
transform 1 0 240396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2613
timestamp 1676037725
transform 1 0 241500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2625
timestamp 1676037725
transform 1 0 242604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2631
timestamp 1676037725
transform 1 0 243156 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2633
timestamp 1676037725
transform 1 0 243340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2645
timestamp 1676037725
transform 1 0 244444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2657
timestamp 1676037725
transform 1 0 245548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2669
timestamp 1676037725
transform 1 0 246652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2681
timestamp 1676037725
transform 1 0 247756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2687
timestamp 1676037725
transform 1 0 248308 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2689
timestamp 1676037725
transform 1 0 248492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2701
timestamp 1676037725
transform 1 0 249596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2713
timestamp 1676037725
transform 1 0 250700 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2725
timestamp 1676037725
transform 1 0 251804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2737
timestamp 1676037725
transform 1 0 252908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2743
timestamp 1676037725
transform 1 0 253460 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2745
timestamp 1676037725
transform 1 0 253644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2757
timestamp 1676037725
transform 1 0 254748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2769
timestamp 1676037725
transform 1 0 255852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2781
timestamp 1676037725
transform 1 0 256956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2793
timestamp 1676037725
transform 1 0 258060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2799
timestamp 1676037725
transform 1 0 258612 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2801
timestamp 1676037725
transform 1 0 258796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2813
timestamp 1676037725
transform 1 0 259900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2825
timestamp 1676037725
transform 1 0 261004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2837
timestamp 1676037725
transform 1 0 262108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2849
timestamp 1676037725
transform 1 0 263212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2855
timestamp 1676037725
transform 1 0 263764 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2857
timestamp 1676037725
transform 1 0 263948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2869
timestamp 1676037725
transform 1 0 265052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2881
timestamp 1676037725
transform 1 0 266156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2893
timestamp 1676037725
transform 1 0 267260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2905
timestamp 1676037725
transform 1 0 268364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2911
timestamp 1676037725
transform 1 0 268916 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2913
timestamp 1676037725
transform 1 0 269100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2925
timestamp 1676037725
transform 1 0 270204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2937
timestamp 1676037725
transform 1 0 271308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2949
timestamp 1676037725
transform 1 0 272412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_2961
timestamp 1676037725
transform 1 0 273516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_2967
timestamp 1676037725
transform 1 0 274068 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2969
timestamp 1676037725
transform 1 0 274252 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2981
timestamp 1676037725
transform 1 0 275356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_2993
timestamp 1676037725
transform 1 0 276460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3005
timestamp 1676037725
transform 1 0 277564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3017
timestamp 1676037725
transform 1 0 278668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3023
timestamp 1676037725
transform 1 0 279220 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3025
timestamp 1676037725
transform 1 0 279404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3037
timestamp 1676037725
transform 1 0 280508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3049
timestamp 1676037725
transform 1 0 281612 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3061
timestamp 1676037725
transform 1 0 282716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3073
timestamp 1676037725
transform 1 0 283820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3079
timestamp 1676037725
transform 1 0 284372 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3081
timestamp 1676037725
transform 1 0 284556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3093
timestamp 1676037725
transform 1 0 285660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3105
timestamp 1676037725
transform 1 0 286764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3117
timestamp 1676037725
transform 1 0 287868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3129
timestamp 1676037725
transform 1 0 288972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3135
timestamp 1676037725
transform 1 0 289524 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3137
timestamp 1676037725
transform 1 0 289708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3149
timestamp 1676037725
transform 1 0 290812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3161
timestamp 1676037725
transform 1 0 291916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3173
timestamp 1676037725
transform 1 0 293020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3185
timestamp 1676037725
transform 1 0 294124 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3191
timestamp 1676037725
transform 1 0 294676 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3193
timestamp 1676037725
transform 1 0 294860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3205
timestamp 1676037725
transform 1 0 295964 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3217
timestamp 1676037725
transform 1 0 297068 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3229
timestamp 1676037725
transform 1 0 298172 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3241
timestamp 1676037725
transform 1 0 299276 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3247
timestamp 1676037725
transform 1 0 299828 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3249
timestamp 1676037725
transform 1 0 300012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3261
timestamp 1676037725
transform 1 0 301116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3273
timestamp 1676037725
transform 1 0 302220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3285
timestamp 1676037725
transform 1 0 303324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3297
timestamp 1676037725
transform 1 0 304428 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3303
timestamp 1676037725
transform 1 0 304980 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3305
timestamp 1676037725
transform 1 0 305164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3317
timestamp 1676037725
transform 1 0 306268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3329
timestamp 1676037725
transform 1 0 307372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3341
timestamp 1676037725
transform 1 0 308476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3353
timestamp 1676037725
transform 1 0 309580 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3359
timestamp 1676037725
transform 1 0 310132 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3361
timestamp 1676037725
transform 1 0 310316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3373
timestamp 1676037725
transform 1 0 311420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3385
timestamp 1676037725
transform 1 0 312524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3397
timestamp 1676037725
transform 1 0 313628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3409
timestamp 1676037725
transform 1 0 314732 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3415
timestamp 1676037725
transform 1 0 315284 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3417
timestamp 1676037725
transform 1 0 315468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3429
timestamp 1676037725
transform 1 0 316572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3441
timestamp 1676037725
transform 1 0 317676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3453
timestamp 1676037725
transform 1 0 318780 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3465
timestamp 1676037725
transform 1 0 319884 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3471
timestamp 1676037725
transform 1 0 320436 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3473
timestamp 1676037725
transform 1 0 320620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3485
timestamp 1676037725
transform 1 0 321724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3497
timestamp 1676037725
transform 1 0 322828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3509
timestamp 1676037725
transform 1 0 323932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3521
timestamp 1676037725
transform 1 0 325036 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3527
timestamp 1676037725
transform 1 0 325588 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3529
timestamp 1676037725
transform 1 0 325772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3541
timestamp 1676037725
transform 1 0 326876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3553
timestamp 1676037725
transform 1 0 327980 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3565
timestamp 1676037725
transform 1 0 329084 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3577
timestamp 1676037725
transform 1 0 330188 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3583
timestamp 1676037725
transform 1 0 330740 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3585
timestamp 1676037725
transform 1 0 330924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3597
timestamp 1676037725
transform 1 0 332028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3609
timestamp 1676037725
transform 1 0 333132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3621
timestamp 1676037725
transform 1 0 334236 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3633
timestamp 1676037725
transform 1 0 335340 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3639
timestamp 1676037725
transform 1 0 335892 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3641
timestamp 1676037725
transform 1 0 336076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3653
timestamp 1676037725
transform 1 0 337180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3665
timestamp 1676037725
transform 1 0 338284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3677
timestamp 1676037725
transform 1 0 339388 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3689
timestamp 1676037725
transform 1 0 340492 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3695
timestamp 1676037725
transform 1 0 341044 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3697
timestamp 1676037725
transform 1 0 341228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3709
timestamp 1676037725
transform 1 0 342332 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3721
timestamp 1676037725
transform 1 0 343436 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3733
timestamp 1676037725
transform 1 0 344540 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3745
timestamp 1676037725
transform 1 0 345644 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3751
timestamp 1676037725
transform 1 0 346196 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3753
timestamp 1676037725
transform 1 0 346380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3765
timestamp 1676037725
transform 1 0 347484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3777
timestamp 1676037725
transform 1 0 348588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3789
timestamp 1676037725
transform 1 0 349692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3801
timestamp 1676037725
transform 1 0 350796 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3807
timestamp 1676037725
transform 1 0 351348 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3809
timestamp 1676037725
transform 1 0 351532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3821
timestamp 1676037725
transform 1 0 352636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3833
timestamp 1676037725
transform 1 0 353740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3845
timestamp 1676037725
transform 1 0 354844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3857
timestamp 1676037725
transform 1 0 355948 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3863
timestamp 1676037725
transform 1 0 356500 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3865
timestamp 1676037725
transform 1 0 356684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3877
timestamp 1676037725
transform 1 0 357788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3889
timestamp 1676037725
transform 1 0 358892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3901
timestamp 1676037725
transform 1 0 359996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3913
timestamp 1676037725
transform 1 0 361100 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3919
timestamp 1676037725
transform 1 0 361652 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3921
timestamp 1676037725
transform 1 0 361836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3933
timestamp 1676037725
transform 1 0 362940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3945
timestamp 1676037725
transform 1 0 364044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3957
timestamp 1676037725
transform 1 0 365148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3969
timestamp 1676037725
transform 1 0 366252 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3975
timestamp 1676037725
transform 1 0 366804 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3977
timestamp 1676037725
transform 1 0 366988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3989
timestamp 1676037725
transform 1 0 368092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4001
timestamp 1676037725
transform 1 0 369196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4013
timestamp 1676037725
transform 1 0 370300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4025
timestamp 1676037725
transform 1 0 371404 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4031
timestamp 1676037725
transform 1 0 371956 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4033
timestamp 1676037725
transform 1 0 372140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4045
timestamp 1676037725
transform 1 0 373244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4057
timestamp 1676037725
transform 1 0 374348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4069
timestamp 1676037725
transform 1 0 375452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4081
timestamp 1676037725
transform 1 0 376556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4087
timestamp 1676037725
transform 1 0 377108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4089
timestamp 1676037725
transform 1 0 377292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4101
timestamp 1676037725
transform 1 0 378396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4113
timestamp 1676037725
transform 1 0 379500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4125
timestamp 1676037725
transform 1 0 380604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4137
timestamp 1676037725
transform 1 0 381708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4143
timestamp 1676037725
transform 1 0 382260 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4145
timestamp 1676037725
transform 1 0 382444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4157
timestamp 1676037725
transform 1 0 383548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4169
timestamp 1676037725
transform 1 0 384652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4181
timestamp 1676037725
transform 1 0 385756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4193
timestamp 1676037725
transform 1 0 386860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4199
timestamp 1676037725
transform 1 0 387412 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4201
timestamp 1676037725
transform 1 0 387596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4213
timestamp 1676037725
transform 1 0 388700 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4225
timestamp 1676037725
transform 1 0 389804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4237
timestamp 1676037725
transform 1 0 390908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4249
timestamp 1676037725
transform 1 0 392012 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4255
timestamp 1676037725
transform 1 0 392564 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4257
timestamp 1676037725
transform 1 0 392748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4269
timestamp 1676037725
transform 1 0 393852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4281
timestamp 1676037725
transform 1 0 394956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4293
timestamp 1676037725
transform 1 0 396060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4305
timestamp 1676037725
transform 1 0 397164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4311
timestamp 1676037725
transform 1 0 397716 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4313
timestamp 1676037725
transform 1 0 397900 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4325
timestamp 1676037725
transform 1 0 399004 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4337
timestamp 1676037725
transform 1 0 400108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4349
timestamp 1676037725
transform 1 0 401212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4361
timestamp 1676037725
transform 1 0 402316 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4367
timestamp 1676037725
transform 1 0 402868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4369
timestamp 1676037725
transform 1 0 403052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4381
timestamp 1676037725
transform 1 0 404156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4393
timestamp 1676037725
transform 1 0 405260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4405
timestamp 1676037725
transform 1 0 406364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4417
timestamp 1676037725
transform 1 0 407468 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4423
timestamp 1676037725
transform 1 0 408020 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4425
timestamp 1676037725
transform 1 0 408204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4437
timestamp 1676037725
transform 1 0 409308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4449
timestamp 1676037725
transform 1 0 410412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4461
timestamp 1676037725
transform 1 0 411516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4473
timestamp 1676037725
transform 1 0 412620 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4479
timestamp 1676037725
transform 1 0 413172 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4481
timestamp 1676037725
transform 1 0 413356 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4493
timestamp 1676037725
transform 1 0 414460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4505
timestamp 1676037725
transform 1 0 415564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4517
timestamp 1676037725
transform 1 0 416668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4529
timestamp 1676037725
transform 1 0 417772 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4535
timestamp 1676037725
transform 1 0 418324 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4537
timestamp 1676037725
transform 1 0 418508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4549
timestamp 1676037725
transform 1 0 419612 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4561
timestamp 1676037725
transform 1 0 420716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4573
timestamp 1676037725
transform 1 0 421820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4585
timestamp 1676037725
transform 1 0 422924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4591
timestamp 1676037725
transform 1 0 423476 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4593
timestamp 1676037725
transform 1 0 423660 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4605
timestamp 1676037725
transform 1 0 424764 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4617
timestamp 1676037725
transform 1 0 425868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4629
timestamp 1676037725
transform 1 0 426972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4641
timestamp 1676037725
transform 1 0 428076 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4647
timestamp 1676037725
transform 1 0 428628 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4649
timestamp 1676037725
transform 1 0 428812 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4661
timestamp 1676037725
transform 1 0 429916 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4673
timestamp 1676037725
transform 1 0 431020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4685
timestamp 1676037725
transform 1 0 432124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4697
timestamp 1676037725
transform 1 0 433228 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4703
timestamp 1676037725
transform 1 0 433780 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4705
timestamp 1676037725
transform 1 0 433964 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4717
timestamp 1676037725
transform 1 0 435068 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4729
timestamp 1676037725
transform 1 0 436172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4741
timestamp 1676037725
transform 1 0 437276 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4753
timestamp 1676037725
transform 1 0 438380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4759
timestamp 1676037725
transform 1 0 438932 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4761
timestamp 1676037725
transform 1 0 439116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4773
timestamp 1676037725
transform 1 0 440220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4785
timestamp 1676037725
transform 1 0 441324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4797
timestamp 1676037725
transform 1 0 442428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4809
timestamp 1676037725
transform 1 0 443532 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4815
timestamp 1676037725
transform 1 0 444084 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4817
timestamp 1676037725
transform 1 0 444268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4829
timestamp 1676037725
transform 1 0 445372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4841
timestamp 1676037725
transform 1 0 446476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4853
timestamp 1676037725
transform 1 0 447580 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4865
timestamp 1676037725
transform 1 0 448684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4871
timestamp 1676037725
transform 1 0 449236 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4873
timestamp 1676037725
transform 1 0 449420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4885
timestamp 1676037725
transform 1 0 450524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4897
timestamp 1676037725
transform 1 0 451628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4909
timestamp 1676037725
transform 1 0 452732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4921
timestamp 1676037725
transform 1 0 453836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4927
timestamp 1676037725
transform 1 0 454388 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4929
timestamp 1676037725
transform 1 0 454572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4941
timestamp 1676037725
transform 1 0 455676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4953
timestamp 1676037725
transform 1 0 456780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4965
timestamp 1676037725
transform 1 0 457884 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_4977
timestamp 1676037725
transform 1 0 458988 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_4983
timestamp 1676037725
transform 1 0 459540 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4985
timestamp 1676037725
transform 1 0 459724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_4997
timestamp 1676037725
transform 1 0 460828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5009
timestamp 1676037725
transform 1 0 461932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5021
timestamp 1676037725
transform 1 0 463036 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5033
timestamp 1676037725
transform 1 0 464140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5039
timestamp 1676037725
transform 1 0 464692 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5041
timestamp 1676037725
transform 1 0 464876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5053
timestamp 1676037725
transform 1 0 465980 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5065
timestamp 1676037725
transform 1 0 467084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5077
timestamp 1676037725
transform 1 0 468188 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5089
timestamp 1676037725
transform 1 0 469292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5095
timestamp 1676037725
transform 1 0 469844 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5097
timestamp 1676037725
transform 1 0 470028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5109
timestamp 1676037725
transform 1 0 471132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5121
timestamp 1676037725
transform 1 0 472236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5133
timestamp 1676037725
transform 1 0 473340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5145
timestamp 1676037725
transform 1 0 474444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5151
timestamp 1676037725
transform 1 0 474996 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5153
timestamp 1676037725
transform 1 0 475180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5165
timestamp 1676037725
transform 1 0 476284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5177
timestamp 1676037725
transform 1 0 477388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5189
timestamp 1676037725
transform 1 0 478492 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5201
timestamp 1676037725
transform 1 0 479596 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5207
timestamp 1676037725
transform 1 0 480148 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5209
timestamp 1676037725
transform 1 0 480332 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5221
timestamp 1676037725
transform 1 0 481436 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5233
timestamp 1676037725
transform 1 0 482540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5245
timestamp 1676037725
transform 1 0 483644 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5257
timestamp 1676037725
transform 1 0 484748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5263
timestamp 1676037725
transform 1 0 485300 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5265
timestamp 1676037725
transform 1 0 485484 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5271
timestamp 1676037725
transform 1 0 486036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5283
timestamp 1676037725
transform 1 0 487140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5295
timestamp 1676037725
transform 1 0 488244 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5299
timestamp 1676037725
transform 1 0 488612 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5311
timestamp 1676037725
transform 1 0 489716 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5319
timestamp 1676037725
transform 1 0 490452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5321
timestamp 1676037725
transform 1 0 490636 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5327
timestamp 1676037725
transform 1 0 491188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5339
timestamp 1676037725
transform 1 0 492292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5351
timestamp 1676037725
transform 1 0 493396 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5355
timestamp 1676037725
transform 1 0 493764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5367
timestamp 1676037725
transform 1 0 494868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5375
timestamp 1676037725
transform 1 0 495604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5377
timestamp 1676037725
transform 1 0 495788 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5383
timestamp 1676037725
transform 1 0 496340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5395
timestamp 1676037725
transform 1 0 497444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5407
timestamp 1676037725
transform 1 0 498548 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5411
timestamp 1676037725
transform 1 0 498916 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5423
timestamp 1676037725
transform 1 0 500020 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5431
timestamp 1676037725
transform 1 0 500756 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5433
timestamp 1676037725
transform 1 0 500940 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5439
timestamp 1676037725
transform 1 0 501492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5451
timestamp 1676037725
transform 1 0 502596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5463
timestamp 1676037725
transform 1 0 503700 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5467
timestamp 1676037725
transform 1 0 504068 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5479
timestamp 1676037725
transform 1 0 505172 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5487
timestamp 1676037725
transform 1 0 505908 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5489
timestamp 1676037725
transform 1 0 506092 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5495
timestamp 1676037725
transform 1 0 506644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5507
timestamp 1676037725
transform 1 0 507748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5519
timestamp 1676037725
transform 1 0 508852 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5523
timestamp 1676037725
transform 1 0 509220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5535
timestamp 1676037725
transform 1 0 510324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5543
timestamp 1676037725
transform 1 0 511060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5545
timestamp 1676037725
transform 1 0 511244 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5551
timestamp 1676037725
transform 1 0 511796 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5563
timestamp 1676037725
transform 1 0 512900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5575
timestamp 1676037725
transform 1 0 514004 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5579
timestamp 1676037725
transform 1 0 514372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5591
timestamp 1676037725
transform 1 0 515476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5599
timestamp 1676037725
transform 1 0 516212 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5601
timestamp 1676037725
transform 1 0 516396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5613
timestamp 1676037725
transform 1 0 517500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5625
timestamp 1676037725
transform 1 0 518604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5637
timestamp 1676037725
transform 1 0 519708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5649
timestamp 1676037725
transform 1 0 520812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5655
timestamp 1676037725
transform 1 0 521364 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5657
timestamp 1676037725
transform 1 0 521548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5669
timestamp 1676037725
transform 1 0 522652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5681
timestamp 1676037725
transform 1 0 523756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5693
timestamp 1676037725
transform 1 0 524860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_5705
timestamp 1676037725
transform 1 0 525964 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_5711
timestamp 1676037725
transform 1 0 526516 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5713
timestamp 1676037725
transform 1 0 526700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_5725
timestamp 1676037725
transform 1 0 527804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_11
timestamp 1676037725
transform 1 0 2116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1676037725
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_39
timestamp 1676037725
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1676037725
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_67
timestamp 1676037725
transform 1 0 7268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1676037725
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_95
timestamp 1676037725
transform 1 0 9844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1676037725
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_113
timestamp 1676037725
transform 1 0 11500 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_123
timestamp 1676037725
transform 1 0 12420 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1676037725
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_151
timestamp 1676037725
transform 1 0 14996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1676037725
transform 1 0 16100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_169
timestamp 1676037725
transform 1 0 16652 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1676037725
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_207
timestamp 1676037725
transform 1 0 20148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_225
timestamp 1676037725
transform 1 0 21804 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1676037725
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_263
timestamp 1676037725
transform 1 0 25300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_275
timestamp 1676037725
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_281
timestamp 1676037725
transform 1 0 26956 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_291
timestamp 1676037725
transform 1 0 27876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1676037725
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_319
timestamp 1676037725
transform 1 0 30452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_331
timestamp 1676037725
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_337
timestamp 1676037725
transform 1 0 32108 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_347
timestamp 1676037725
transform 1 0 33028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_359
timestamp 1676037725
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_375
timestamp 1676037725
transform 1 0 35604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_381
timestamp 1676037725
transform 1 0 36156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_393
timestamp 1676037725
transform 1 0 37260 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_403
timestamp 1676037725
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1676037725
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_431
timestamp 1676037725
transform 1 0 40756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_443
timestamp 1676037725
transform 1 0 41860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_459
timestamp 1676037725
transform 1 0 43332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_465
timestamp 1676037725
transform 1 0 43884 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1676037725
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_487
timestamp 1676037725
transform 1 0 45908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_499
timestamp 1676037725
transform 1 0 47012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_507
timestamp 1676037725
transform 1 0 47748 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_515
timestamp 1676037725
transform 1 0 48484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_527
timestamp 1676037725
transform 1 0 49588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1676037725
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_543
timestamp 1676037725
transform 1 0 51060 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_549
timestamp 1676037725
transform 1 0 51612 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_563
timestamp 1676037725
transform 1 0 52900 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_571
timestamp 1676037725
transform 1 0 53636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_583
timestamp 1676037725
transform 1 0 54740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1676037725
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_599
timestamp 1676037725
transform 1 0 56212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_611
timestamp 1676037725
transform 1 0 57316 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_627
timestamp 1676037725
transform 1 0 58788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_633
timestamp 1676037725
transform 1 0 59340 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_641
timestamp 1676037725
transform 1 0 60076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_645
timestamp 1676037725
transform 1 0 60444 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_655
timestamp 1676037725
transform 1 0 61364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_667
timestamp 1676037725
transform 1 0 62468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_675
timestamp 1676037725
transform 1 0 63204 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_683
timestamp 1676037725
transform 1 0 63940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_695
timestamp 1676037725
transform 1 0 65044 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1676037725
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_701
timestamp 1676037725
transform 1 0 65596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_711
timestamp 1676037725
transform 1 0 66516 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_717
timestamp 1676037725
transform 1 0 67068 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_731
timestamp 1676037725
transform 1 0 68356 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_739
timestamp 1676037725
transform 1 0 69092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_751
timestamp 1676037725
transform 1 0 70196 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1676037725
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_757
timestamp 1676037725
transform 1 0 70748 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_767
timestamp 1676037725
transform 1 0 71668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_779
timestamp 1676037725
transform 1 0 72772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_795
timestamp 1676037725
transform 1 0 74244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_801
timestamp 1676037725
transform 1 0 74796 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_809
timestamp 1676037725
transform 1 0 75532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_813
timestamp 1676037725
transform 1 0 75900 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_823
timestamp 1676037725
transform 1 0 76820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_835
timestamp 1676037725
transform 1 0 77924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_843
timestamp 1676037725
transform 1 0 78660 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_851
timestamp 1676037725
transform 1 0 79396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_863
timestamp 1676037725
transform 1 0 80500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1676037725
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_869
timestamp 1676037725
transform 1 0 81052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_879
timestamp 1676037725
transform 1 0 81972 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_885
timestamp 1676037725
transform 1 0 82524 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_899
timestamp 1676037725
transform 1 0 83812 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_907
timestamp 1676037725
transform 1 0 84548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_919
timestamp 1676037725
transform 1 0 85652 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1676037725
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_925
timestamp 1676037725
transform 1 0 86204 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_935
timestamp 1676037725
transform 1 0 87124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_947
timestamp 1676037725
transform 1 0 88228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_963
timestamp 1676037725
transform 1 0 89700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_969
timestamp 1676037725
transform 1 0 90252 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_977
timestamp 1676037725
transform 1 0 90988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_981
timestamp 1676037725
transform 1 0 91356 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_991
timestamp 1676037725
transform 1 0 92276 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1003
timestamp 1676037725
transform 1 0 93380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1011
timestamp 1676037725
transform 1 0 94116 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1019
timestamp 1676037725
transform 1 0 94852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1031
timestamp 1676037725
transform 1 0 95956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1676037725
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1037
timestamp 1676037725
transform 1 0 96508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1047
timestamp 1676037725
transform 1 0 97428 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1053
timestamp 1676037725
transform 1 0 97980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1067
timestamp 1676037725
transform 1 0 99268 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1075
timestamp 1676037725
transform 1 0 100004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1087
timestamp 1676037725
transform 1 0 101108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1676037725
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1093
timestamp 1676037725
transform 1 0 101660 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1103
timestamp 1676037725
transform 1 0 102580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1115
timestamp 1676037725
transform 1 0 103684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1131
timestamp 1676037725
transform 1 0 105156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1137
timestamp 1676037725
transform 1 0 105708 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1145
timestamp 1676037725
transform 1 0 106444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1149
timestamp 1676037725
transform 1 0 106812 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1159
timestamp 1676037725
transform 1 0 107732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1171
timestamp 1676037725
transform 1 0 108836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1179
timestamp 1676037725
transform 1 0 109572 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1187
timestamp 1676037725
transform 1 0 110308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1199
timestamp 1676037725
transform 1 0 111412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1676037725
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1205
timestamp 1676037725
transform 1 0 111964 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1215
timestamp 1676037725
transform 1 0 112884 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1221
timestamp 1676037725
transform 1 0 113436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1235
timestamp 1676037725
transform 1 0 114724 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1243
timestamp 1676037725
transform 1 0 115460 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1255
timestamp 1676037725
transform 1 0 116564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1259
timestamp 1676037725
transform 1 0 116932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1261
timestamp 1676037725
transform 1 0 117116 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1271
timestamp 1676037725
transform 1 0 118036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1283
timestamp 1676037725
transform 1 0 119140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1299
timestamp 1676037725
transform 1 0 120612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1305
timestamp 1676037725
transform 1 0 121164 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1313
timestamp 1676037725
transform 1 0 121900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1317
timestamp 1676037725
transform 1 0 122268 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1327
timestamp 1676037725
transform 1 0 123188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1339
timestamp 1676037725
transform 1 0 124292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1347
timestamp 1676037725
transform 1 0 125028 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1355
timestamp 1676037725
transform 1 0 125764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1367
timestamp 1676037725
transform 1 0 126868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1371
timestamp 1676037725
transform 1 0 127236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1373
timestamp 1676037725
transform 1 0 127420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1383
timestamp 1676037725
transform 1 0 128340 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1389
timestamp 1676037725
transform 1 0 128892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1401
timestamp 1676037725
transform 1 0 129996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1407
timestamp 1676037725
transform 1 0 130548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1411
timestamp 1676037725
transform 1 0 130916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1417
timestamp 1676037725
transform 1 0 131468 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1425
timestamp 1676037725
transform 1 0 132204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1429
timestamp 1676037725
transform 1 0 132572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1435
timestamp 1676037725
transform 1 0 133124 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1439
timestamp 1676037725
transform 1 0 133492 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1445
timestamp 1676037725
transform 1 0 134044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1457
timestamp 1676037725
transform 1 0 135148 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1467
timestamp 1676037725
transform 1 0 136068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1473
timestamp 1676037725
transform 1 0 136620 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1481
timestamp 1676037725
transform 1 0 137356 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1485
timestamp 1676037725
transform 1 0 137724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1497
timestamp 1676037725
transform 1 0 138828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1509
timestamp 1676037725
transform 1 0 139932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1521
timestamp 1676037725
transform 1 0 141036 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1533
timestamp 1676037725
transform 1 0 142140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1539
timestamp 1676037725
transform 1 0 142692 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1541
timestamp 1676037725
transform 1 0 142876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1553
timestamp 1676037725
transform 1 0 143980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1565
timestamp 1676037725
transform 1 0 145084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1577
timestamp 1676037725
transform 1 0 146188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1589
timestamp 1676037725
transform 1 0 147292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1595
timestamp 1676037725
transform 1 0 147844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1597
timestamp 1676037725
transform 1 0 148028 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1601
timestamp 1676037725
transform 1 0 148396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1613
timestamp 1676037725
transform 1 0 149500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1625
timestamp 1676037725
transform 1 0 150604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1637
timestamp 1676037725
transform 1 0 151708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1649
timestamp 1676037725
transform 1 0 152812 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1653
timestamp 1676037725
transform 1 0 153180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1665
timestamp 1676037725
transform 1 0 154284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1677
timestamp 1676037725
transform 1 0 155388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1689
timestamp 1676037725
transform 1 0 156492 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1701
timestamp 1676037725
transform 1 0 157596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1707
timestamp 1676037725
transform 1 0 158148 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1709
timestamp 1676037725
transform 1 0 158332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1721
timestamp 1676037725
transform 1 0 159436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1733
timestamp 1676037725
transform 1 0 160540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1745
timestamp 1676037725
transform 1 0 161644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1757
timestamp 1676037725
transform 1 0 162748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1763
timestamp 1676037725
transform 1 0 163300 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1765
timestamp 1676037725
transform 1 0 163484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1777
timestamp 1676037725
transform 1 0 164588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1789
timestamp 1676037725
transform 1 0 165692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1801
timestamp 1676037725
transform 1 0 166796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1813
timestamp 1676037725
transform 1 0 167900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1819
timestamp 1676037725
transform 1 0 168452 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1821
timestamp 1676037725
transform 1 0 168636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1833
timestamp 1676037725
transform 1 0 169740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1845
timestamp 1676037725
transform 1 0 170844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1857
timestamp 1676037725
transform 1 0 171948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1869
timestamp 1676037725
transform 1 0 173052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1875
timestamp 1676037725
transform 1 0 173604 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1877
timestamp 1676037725
transform 1 0 173788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1889
timestamp 1676037725
transform 1 0 174892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1901
timestamp 1676037725
transform 1 0 175996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1913
timestamp 1676037725
transform 1 0 177100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1925
timestamp 1676037725
transform 1 0 178204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1931
timestamp 1676037725
transform 1 0 178756 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1933
timestamp 1676037725
transform 1 0 178940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1945
timestamp 1676037725
transform 1 0 180044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1957
timestamp 1676037725
transform 1 0 181148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1969
timestamp 1676037725
transform 1 0 182252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1981
timestamp 1676037725
transform 1 0 183356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1987
timestamp 1676037725
transform 1 0 183908 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1989
timestamp 1676037725
transform 1 0 184092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2001
timestamp 1676037725
transform 1 0 185196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2013
timestamp 1676037725
transform 1 0 186300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2025
timestamp 1676037725
transform 1 0 187404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2037
timestamp 1676037725
transform 1 0 188508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2043
timestamp 1676037725
transform 1 0 189060 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2045
timestamp 1676037725
transform 1 0 189244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2057
timestamp 1676037725
transform 1 0 190348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2069
timestamp 1676037725
transform 1 0 191452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2081
timestamp 1676037725
transform 1 0 192556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2093
timestamp 1676037725
transform 1 0 193660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2099
timestamp 1676037725
transform 1 0 194212 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2101
timestamp 1676037725
transform 1 0 194396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2113
timestamp 1676037725
transform 1 0 195500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2125
timestamp 1676037725
transform 1 0 196604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2137
timestamp 1676037725
transform 1 0 197708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2149
timestamp 1676037725
transform 1 0 198812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2155
timestamp 1676037725
transform 1 0 199364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2157
timestamp 1676037725
transform 1 0 199548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2169
timestamp 1676037725
transform 1 0 200652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2181
timestamp 1676037725
transform 1 0 201756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2193
timestamp 1676037725
transform 1 0 202860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2205
timestamp 1676037725
transform 1 0 203964 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2211
timestamp 1676037725
transform 1 0 204516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2213
timestamp 1676037725
transform 1 0 204700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2225
timestamp 1676037725
transform 1 0 205804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2237
timestamp 1676037725
transform 1 0 206908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2249
timestamp 1676037725
transform 1 0 208012 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2261
timestamp 1676037725
transform 1 0 209116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2267
timestamp 1676037725
transform 1 0 209668 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2269
timestamp 1676037725
transform 1 0 209852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2281
timestamp 1676037725
transform 1 0 210956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2293
timestamp 1676037725
transform 1 0 212060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2305
timestamp 1676037725
transform 1 0 213164 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2317
timestamp 1676037725
transform 1 0 214268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2323
timestamp 1676037725
transform 1 0 214820 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2325
timestamp 1676037725
transform 1 0 215004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2337
timestamp 1676037725
transform 1 0 216108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2349
timestamp 1676037725
transform 1 0 217212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2361
timestamp 1676037725
transform 1 0 218316 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2373
timestamp 1676037725
transform 1 0 219420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2379
timestamp 1676037725
transform 1 0 219972 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2381
timestamp 1676037725
transform 1 0 220156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2393
timestamp 1676037725
transform 1 0 221260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2405
timestamp 1676037725
transform 1 0 222364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2417
timestamp 1676037725
transform 1 0 223468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2429
timestamp 1676037725
transform 1 0 224572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2435
timestamp 1676037725
transform 1 0 225124 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2437
timestamp 1676037725
transform 1 0 225308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2449
timestamp 1676037725
transform 1 0 226412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2461
timestamp 1676037725
transform 1 0 227516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2473
timestamp 1676037725
transform 1 0 228620 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2485
timestamp 1676037725
transform 1 0 229724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2491
timestamp 1676037725
transform 1 0 230276 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2493
timestamp 1676037725
transform 1 0 230460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2505
timestamp 1676037725
transform 1 0 231564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2517
timestamp 1676037725
transform 1 0 232668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2529
timestamp 1676037725
transform 1 0 233772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2541
timestamp 1676037725
transform 1 0 234876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2547
timestamp 1676037725
transform 1 0 235428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2549
timestamp 1676037725
transform 1 0 235612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2561
timestamp 1676037725
transform 1 0 236716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2573
timestamp 1676037725
transform 1 0 237820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2585
timestamp 1676037725
transform 1 0 238924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2597
timestamp 1676037725
transform 1 0 240028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2603
timestamp 1676037725
transform 1 0 240580 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2605
timestamp 1676037725
transform 1 0 240764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2617
timestamp 1676037725
transform 1 0 241868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2629
timestamp 1676037725
transform 1 0 242972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2641
timestamp 1676037725
transform 1 0 244076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2653
timestamp 1676037725
transform 1 0 245180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2659
timestamp 1676037725
transform 1 0 245732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2661
timestamp 1676037725
transform 1 0 245916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2673
timestamp 1676037725
transform 1 0 247020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2685
timestamp 1676037725
transform 1 0 248124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2697
timestamp 1676037725
transform 1 0 249228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2709
timestamp 1676037725
transform 1 0 250332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2715
timestamp 1676037725
transform 1 0 250884 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2717
timestamp 1676037725
transform 1 0 251068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2729
timestamp 1676037725
transform 1 0 252172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2741
timestamp 1676037725
transform 1 0 253276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2753
timestamp 1676037725
transform 1 0 254380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2765
timestamp 1676037725
transform 1 0 255484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2771
timestamp 1676037725
transform 1 0 256036 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2773
timestamp 1676037725
transform 1 0 256220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2785
timestamp 1676037725
transform 1 0 257324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2797
timestamp 1676037725
transform 1 0 258428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2809
timestamp 1676037725
transform 1 0 259532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2821
timestamp 1676037725
transform 1 0 260636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2827
timestamp 1676037725
transform 1 0 261188 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2829
timestamp 1676037725
transform 1 0 261372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2841
timestamp 1676037725
transform 1 0 262476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2853
timestamp 1676037725
transform 1 0 263580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2865
timestamp 1676037725
transform 1 0 264684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2877
timestamp 1676037725
transform 1 0 265788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2883
timestamp 1676037725
transform 1 0 266340 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2885
timestamp 1676037725
transform 1 0 266524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2897
timestamp 1676037725
transform 1 0 267628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2909
timestamp 1676037725
transform 1 0 268732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2921
timestamp 1676037725
transform 1 0 269836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2933
timestamp 1676037725
transform 1 0 270940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2939
timestamp 1676037725
transform 1 0 271492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2941
timestamp 1676037725
transform 1 0 271676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2953
timestamp 1676037725
transform 1 0 272780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2965
timestamp 1676037725
transform 1 0 273884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2977
timestamp 1676037725
transform 1 0 274988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_2989
timestamp 1676037725
transform 1 0 276092 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_2995
timestamp 1676037725
transform 1 0 276644 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_2997
timestamp 1676037725
transform 1 0 276828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3009
timestamp 1676037725
transform 1 0 277932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3021
timestamp 1676037725
transform 1 0 279036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3033
timestamp 1676037725
transform 1 0 280140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3045
timestamp 1676037725
transform 1 0 281244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3051
timestamp 1676037725
transform 1 0 281796 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3053
timestamp 1676037725
transform 1 0 281980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3065
timestamp 1676037725
transform 1 0 283084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3077
timestamp 1676037725
transform 1 0 284188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3089
timestamp 1676037725
transform 1 0 285292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3101
timestamp 1676037725
transform 1 0 286396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3107
timestamp 1676037725
transform 1 0 286948 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3109
timestamp 1676037725
transform 1 0 287132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3121
timestamp 1676037725
transform 1 0 288236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3133
timestamp 1676037725
transform 1 0 289340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3145
timestamp 1676037725
transform 1 0 290444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3157
timestamp 1676037725
transform 1 0 291548 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3163
timestamp 1676037725
transform 1 0 292100 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3165
timestamp 1676037725
transform 1 0 292284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3177
timestamp 1676037725
transform 1 0 293388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3189
timestamp 1676037725
transform 1 0 294492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3201
timestamp 1676037725
transform 1 0 295596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3213
timestamp 1676037725
transform 1 0 296700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3219
timestamp 1676037725
transform 1 0 297252 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3221
timestamp 1676037725
transform 1 0 297436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3233
timestamp 1676037725
transform 1 0 298540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3245
timestamp 1676037725
transform 1 0 299644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3257
timestamp 1676037725
transform 1 0 300748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3269
timestamp 1676037725
transform 1 0 301852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3275
timestamp 1676037725
transform 1 0 302404 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3277
timestamp 1676037725
transform 1 0 302588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3289
timestamp 1676037725
transform 1 0 303692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3301
timestamp 1676037725
transform 1 0 304796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3313
timestamp 1676037725
transform 1 0 305900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3325
timestamp 1676037725
transform 1 0 307004 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3331
timestamp 1676037725
transform 1 0 307556 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3333
timestamp 1676037725
transform 1 0 307740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3345
timestamp 1676037725
transform 1 0 308844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3357
timestamp 1676037725
transform 1 0 309948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3369
timestamp 1676037725
transform 1 0 311052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3381
timestamp 1676037725
transform 1 0 312156 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3387
timestamp 1676037725
transform 1 0 312708 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3389
timestamp 1676037725
transform 1 0 312892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3401
timestamp 1676037725
transform 1 0 313996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3413
timestamp 1676037725
transform 1 0 315100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3425
timestamp 1676037725
transform 1 0 316204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3437
timestamp 1676037725
transform 1 0 317308 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3443
timestamp 1676037725
transform 1 0 317860 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3445
timestamp 1676037725
transform 1 0 318044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3457
timestamp 1676037725
transform 1 0 319148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3469
timestamp 1676037725
transform 1 0 320252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3481
timestamp 1676037725
transform 1 0 321356 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3493
timestamp 1676037725
transform 1 0 322460 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3499
timestamp 1676037725
transform 1 0 323012 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3501
timestamp 1676037725
transform 1 0 323196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3513
timestamp 1676037725
transform 1 0 324300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3525
timestamp 1676037725
transform 1 0 325404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3537
timestamp 1676037725
transform 1 0 326508 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3549
timestamp 1676037725
transform 1 0 327612 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3555
timestamp 1676037725
transform 1 0 328164 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3557
timestamp 1676037725
transform 1 0 328348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3569
timestamp 1676037725
transform 1 0 329452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3581
timestamp 1676037725
transform 1 0 330556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3593
timestamp 1676037725
transform 1 0 331660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3605
timestamp 1676037725
transform 1 0 332764 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3611
timestamp 1676037725
transform 1 0 333316 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3613
timestamp 1676037725
transform 1 0 333500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3625
timestamp 1676037725
transform 1 0 334604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3637
timestamp 1676037725
transform 1 0 335708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3649
timestamp 1676037725
transform 1 0 336812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3661
timestamp 1676037725
transform 1 0 337916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3667
timestamp 1676037725
transform 1 0 338468 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3669
timestamp 1676037725
transform 1 0 338652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3681
timestamp 1676037725
transform 1 0 339756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3693
timestamp 1676037725
transform 1 0 340860 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3705
timestamp 1676037725
transform 1 0 341964 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3717
timestamp 1676037725
transform 1 0 343068 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3723
timestamp 1676037725
transform 1 0 343620 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3725
timestamp 1676037725
transform 1 0 343804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3737
timestamp 1676037725
transform 1 0 344908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3749
timestamp 1676037725
transform 1 0 346012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3761
timestamp 1676037725
transform 1 0 347116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3773
timestamp 1676037725
transform 1 0 348220 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3779
timestamp 1676037725
transform 1 0 348772 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3781
timestamp 1676037725
transform 1 0 348956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3793
timestamp 1676037725
transform 1 0 350060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3805
timestamp 1676037725
transform 1 0 351164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3817
timestamp 1676037725
transform 1 0 352268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3829
timestamp 1676037725
transform 1 0 353372 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3835
timestamp 1676037725
transform 1 0 353924 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3837
timestamp 1676037725
transform 1 0 354108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3849
timestamp 1676037725
transform 1 0 355212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3861
timestamp 1676037725
transform 1 0 356316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3873
timestamp 1676037725
transform 1 0 357420 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3885
timestamp 1676037725
transform 1 0 358524 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3891
timestamp 1676037725
transform 1 0 359076 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3893
timestamp 1676037725
transform 1 0 359260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3905
timestamp 1676037725
transform 1 0 360364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3917
timestamp 1676037725
transform 1 0 361468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3929
timestamp 1676037725
transform 1 0 362572 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3941
timestamp 1676037725
transform 1 0 363676 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3947
timestamp 1676037725
transform 1 0 364228 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3949
timestamp 1676037725
transform 1 0 364412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3961
timestamp 1676037725
transform 1 0 365516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3973
timestamp 1676037725
transform 1 0 366620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3985
timestamp 1676037725
transform 1 0 367724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3997
timestamp 1676037725
transform 1 0 368828 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4003
timestamp 1676037725
transform 1 0 369380 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4005
timestamp 1676037725
transform 1 0 369564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4017
timestamp 1676037725
transform 1 0 370668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4029
timestamp 1676037725
transform 1 0 371772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4041
timestamp 1676037725
transform 1 0 372876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4053
timestamp 1676037725
transform 1 0 373980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4059
timestamp 1676037725
transform 1 0 374532 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4061
timestamp 1676037725
transform 1 0 374716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4073
timestamp 1676037725
transform 1 0 375820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4085
timestamp 1676037725
transform 1 0 376924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4097
timestamp 1676037725
transform 1 0 378028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4109
timestamp 1676037725
transform 1 0 379132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4115
timestamp 1676037725
transform 1 0 379684 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4117
timestamp 1676037725
transform 1 0 379868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4129
timestamp 1676037725
transform 1 0 380972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4141
timestamp 1676037725
transform 1 0 382076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4153
timestamp 1676037725
transform 1 0 383180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4165
timestamp 1676037725
transform 1 0 384284 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4171
timestamp 1676037725
transform 1 0 384836 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4173
timestamp 1676037725
transform 1 0 385020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4185
timestamp 1676037725
transform 1 0 386124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4197
timestamp 1676037725
transform 1 0 387228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4209
timestamp 1676037725
transform 1 0 388332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4221
timestamp 1676037725
transform 1 0 389436 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4227
timestamp 1676037725
transform 1 0 389988 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4229
timestamp 1676037725
transform 1 0 390172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4241
timestamp 1676037725
transform 1 0 391276 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4253
timestamp 1676037725
transform 1 0 392380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4265
timestamp 1676037725
transform 1 0 393484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4277
timestamp 1676037725
transform 1 0 394588 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4283
timestamp 1676037725
transform 1 0 395140 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4285
timestamp 1676037725
transform 1 0 395324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4297
timestamp 1676037725
transform 1 0 396428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4309
timestamp 1676037725
transform 1 0 397532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4321
timestamp 1676037725
transform 1 0 398636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4333
timestamp 1676037725
transform 1 0 399740 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4339
timestamp 1676037725
transform 1 0 400292 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4341
timestamp 1676037725
transform 1 0 400476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4353
timestamp 1676037725
transform 1 0 401580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4365
timestamp 1676037725
transform 1 0 402684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4377
timestamp 1676037725
transform 1 0 403788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4389
timestamp 1676037725
transform 1 0 404892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4395
timestamp 1676037725
transform 1 0 405444 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4397
timestamp 1676037725
transform 1 0 405628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4409
timestamp 1676037725
transform 1 0 406732 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4421
timestamp 1676037725
transform 1 0 407836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4433
timestamp 1676037725
transform 1 0 408940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4445
timestamp 1676037725
transform 1 0 410044 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4451
timestamp 1676037725
transform 1 0 410596 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4453
timestamp 1676037725
transform 1 0 410780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4465
timestamp 1676037725
transform 1 0 411884 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4477
timestamp 1676037725
transform 1 0 412988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4489
timestamp 1676037725
transform 1 0 414092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4501
timestamp 1676037725
transform 1 0 415196 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4507
timestamp 1676037725
transform 1 0 415748 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4509
timestamp 1676037725
transform 1 0 415932 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4521
timestamp 1676037725
transform 1 0 417036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4533
timestamp 1676037725
transform 1 0 418140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4545
timestamp 1676037725
transform 1 0 419244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4557
timestamp 1676037725
transform 1 0 420348 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4563
timestamp 1676037725
transform 1 0 420900 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4565
timestamp 1676037725
transform 1 0 421084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4577
timestamp 1676037725
transform 1 0 422188 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4589
timestamp 1676037725
transform 1 0 423292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4601
timestamp 1676037725
transform 1 0 424396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4613
timestamp 1676037725
transform 1 0 425500 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4619
timestamp 1676037725
transform 1 0 426052 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4621
timestamp 1676037725
transform 1 0 426236 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4633
timestamp 1676037725
transform 1 0 427340 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4645
timestamp 1676037725
transform 1 0 428444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4657
timestamp 1676037725
transform 1 0 429548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4669
timestamp 1676037725
transform 1 0 430652 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4675
timestamp 1676037725
transform 1 0 431204 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4677
timestamp 1676037725
transform 1 0 431388 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4689
timestamp 1676037725
transform 1 0 432492 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4701
timestamp 1676037725
transform 1 0 433596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4713
timestamp 1676037725
transform 1 0 434700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4725
timestamp 1676037725
transform 1 0 435804 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4731
timestamp 1676037725
transform 1 0 436356 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4733
timestamp 1676037725
transform 1 0 436540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4745
timestamp 1676037725
transform 1 0 437644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4757
timestamp 1676037725
transform 1 0 438748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4769
timestamp 1676037725
transform 1 0 439852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4781
timestamp 1676037725
transform 1 0 440956 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4787
timestamp 1676037725
transform 1 0 441508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4789
timestamp 1676037725
transform 1 0 441692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4801
timestamp 1676037725
transform 1 0 442796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4813
timestamp 1676037725
transform 1 0 443900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4825
timestamp 1676037725
transform 1 0 445004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4837
timestamp 1676037725
transform 1 0 446108 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4843
timestamp 1676037725
transform 1 0 446660 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4845
timestamp 1676037725
transform 1 0 446844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4857
timestamp 1676037725
transform 1 0 447948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4869
timestamp 1676037725
transform 1 0 449052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4881
timestamp 1676037725
transform 1 0 450156 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4893
timestamp 1676037725
transform 1 0 451260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4899
timestamp 1676037725
transform 1 0 451812 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4901
timestamp 1676037725
transform 1 0 451996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4913
timestamp 1676037725
transform 1 0 453100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4925
timestamp 1676037725
transform 1 0 454204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4937
timestamp 1676037725
transform 1 0 455308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_4949
timestamp 1676037725
transform 1 0 456412 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_4955
timestamp 1676037725
transform 1 0 456964 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4957
timestamp 1676037725
transform 1 0 457148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4969
timestamp 1676037725
transform 1 0 458252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4981
timestamp 1676037725
transform 1 0 459356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_4993
timestamp 1676037725
transform 1 0 460460 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5005
timestamp 1676037725
transform 1 0 461564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5011
timestamp 1676037725
transform 1 0 462116 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5013
timestamp 1676037725
transform 1 0 462300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5025
timestamp 1676037725
transform 1 0 463404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5037
timestamp 1676037725
transform 1 0 464508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5049
timestamp 1676037725
transform 1 0 465612 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5061
timestamp 1676037725
transform 1 0 466716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5067
timestamp 1676037725
transform 1 0 467268 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5069
timestamp 1676037725
transform 1 0 467452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5081
timestamp 1676037725
transform 1 0 468556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5093
timestamp 1676037725
transform 1 0 469660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5105
timestamp 1676037725
transform 1 0 470764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5117
timestamp 1676037725
transform 1 0 471868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5123
timestamp 1676037725
transform 1 0 472420 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5125
timestamp 1676037725
transform 1 0 472604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5137
timestamp 1676037725
transform 1 0 473708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5149
timestamp 1676037725
transform 1 0 474812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5161
timestamp 1676037725
transform 1 0 475916 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5173
timestamp 1676037725
transform 1 0 477020 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5179
timestamp 1676037725
transform 1 0 477572 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5181
timestamp 1676037725
transform 1 0 477756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5193
timestamp 1676037725
transform 1 0 478860 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5205
timestamp 1676037725
transform 1 0 479964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5217
timestamp 1676037725
transform 1 0 481068 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5229
timestamp 1676037725
transform 1 0 482172 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5235
timestamp 1676037725
transform 1 0 482724 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5237
timestamp 1676037725
transform 1 0 482908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5249
timestamp 1676037725
transform 1 0 484012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5261
timestamp 1676037725
transform 1 0 485116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5273
timestamp 1676037725
transform 1 0 486220 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5285
timestamp 1676037725
transform 1 0 487324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5291
timestamp 1676037725
transform 1 0 487876 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5293
timestamp 1676037725
transform 1 0 488060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5305
timestamp 1676037725
transform 1 0 489164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5317
timestamp 1676037725
transform 1 0 490268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5329
timestamp 1676037725
transform 1 0 491372 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5341
timestamp 1676037725
transform 1 0 492476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5347
timestamp 1676037725
transform 1 0 493028 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5349
timestamp 1676037725
transform 1 0 493212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5361
timestamp 1676037725
transform 1 0 494316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5373
timestamp 1676037725
transform 1 0 495420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5385
timestamp 1676037725
transform 1 0 496524 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5397
timestamp 1676037725
transform 1 0 497628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5403
timestamp 1676037725
transform 1 0 498180 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5405
timestamp 1676037725
transform 1 0 498364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5417
timestamp 1676037725
transform 1 0 499468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5429
timestamp 1676037725
transform 1 0 500572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5441
timestamp 1676037725
transform 1 0 501676 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5453
timestamp 1676037725
transform 1 0 502780 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5459
timestamp 1676037725
transform 1 0 503332 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5461
timestamp 1676037725
transform 1 0 503516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5473
timestamp 1676037725
transform 1 0 504620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5485
timestamp 1676037725
transform 1 0 505724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5497
timestamp 1676037725
transform 1 0 506828 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5509
timestamp 1676037725
transform 1 0 507932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5515
timestamp 1676037725
transform 1 0 508484 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5517
timestamp 1676037725
transform 1 0 508668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5529
timestamp 1676037725
transform 1 0 509772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5541
timestamp 1676037725
transform 1 0 510876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5553
timestamp 1676037725
transform 1 0 511980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5565
timestamp 1676037725
transform 1 0 513084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5571
timestamp 1676037725
transform 1 0 513636 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5573
timestamp 1676037725
transform 1 0 513820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5585
timestamp 1676037725
transform 1 0 514924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5597
timestamp 1676037725
transform 1 0 516028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5609
timestamp 1676037725
transform 1 0 517132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5621
timestamp 1676037725
transform 1 0 518236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5627
timestamp 1676037725
transform 1 0 518788 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5629
timestamp 1676037725
transform 1 0 518972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5641
timestamp 1676037725
transform 1 0 520076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5653
timestamp 1676037725
transform 1 0 521180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5665
timestamp 1676037725
transform 1 0 522284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_5677
timestamp 1676037725
transform 1 0 523388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_5683
timestamp 1676037725
transform 1 0 523940 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5685
timestamp 1676037725
transform 1 0 524124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5697
timestamp 1676037725
transform 1 0 525228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5709
timestamp 1676037725
transform 1 0 526332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_5721
timestamp 1676037725
transform 1 0 527436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1676037725
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1676037725
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1676037725
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1676037725
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1676037725
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1676037725
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1676037725
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1676037725
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1676037725
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1676037725
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1676037725
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1676037725
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1676037725
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1676037725
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1676037725
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1676037725
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1676037725
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1676037725
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1676037725
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1676037725
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1676037725
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1676037725
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1676037725
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1676037725
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1676037725
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1676037725
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1676037725
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1676037725
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1676037725
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1676037725
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1676037725
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1676037725
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1676037725
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1676037725
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1676037725
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1676037725
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1676037725
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1676037725
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1676037725
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1676037725
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1676037725
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1676037725
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1676037725
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1676037725
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1676037725
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1676037725
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1676037725
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1676037725
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1676037725
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1676037725
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1676037725
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1676037725
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1676037725
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1676037725
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1676037725
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1676037725
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1676037725
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1676037725
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1676037725
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1676037725
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1676037725
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1676037725
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1676037725
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1676037725
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1676037725
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1676037725
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1676037725
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1676037725
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1676037725
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1676037725
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1676037725
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1676037725
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1676037725
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1676037725
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1676037725
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1676037725
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1257
timestamp 1676037725
transform 1 0 116748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1269
timestamp 1676037725
transform 1 0 117852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1281
timestamp 1676037725
transform 1 0 118956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1287
timestamp 1676037725
transform 1 0 119508 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1289
timestamp 1676037725
transform 1 0 119692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1301
timestamp 1676037725
transform 1 0 120796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1313
timestamp 1676037725
transform 1 0 121900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1325
timestamp 1676037725
transform 1 0 123004 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1337
timestamp 1676037725
transform 1 0 124108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1343
timestamp 1676037725
transform 1 0 124660 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1345
timestamp 1676037725
transform 1 0 124844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1357
timestamp 1676037725
transform 1 0 125948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1369
timestamp 1676037725
transform 1 0 127052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1381
timestamp 1676037725
transform 1 0 128156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1393
timestamp 1676037725
transform 1 0 129260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1399
timestamp 1676037725
transform 1 0 129812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1401
timestamp 1676037725
transform 1 0 129996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1413
timestamp 1676037725
transform 1 0 131100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1425
timestamp 1676037725
transform 1 0 132204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1437
timestamp 1676037725
transform 1 0 133308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1449
timestamp 1676037725
transform 1 0 134412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1455
timestamp 1676037725
transform 1 0 134964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1457
timestamp 1676037725
transform 1 0 135148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1469
timestamp 1676037725
transform 1 0 136252 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1481
timestamp 1676037725
transform 1 0 137356 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1487
timestamp 1676037725
transform 1 0 137908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1499
timestamp 1676037725
transform 1 0 139012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1511
timestamp 1676037725
transform 1 0 140116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1513
timestamp 1676037725
transform 1 0 140300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1521
timestamp 1676037725
transform 1 0 141036 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1524
timestamp 1676037725
transform 1 0 141312 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1536
timestamp 1676037725
transform 1 0 142416 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1546
timestamp 1676037725
transform 1 0 143336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1556
timestamp 1676037725
transform 1 0 144256 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1566
timestamp 1676037725
transform 1 0 145176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1569
timestamp 1676037725
transform 1 0 145452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1577
timestamp 1676037725
transform 1 0 146188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1581
timestamp 1676037725
transform 1 0 146556 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1584
timestamp 1676037725
transform 1 0 146832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1594
timestamp 1676037725
transform 1 0 147752 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1600
timestamp 1676037725
transform 1 0 148304 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1607
timestamp 1676037725
transform 1 0 148948 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1619
timestamp 1676037725
transform 1 0 150052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1623
timestamp 1676037725
transform 1 0 150420 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1625
timestamp 1676037725
transform 1 0 150604 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1633
timestamp 1676037725
transform 1 0 151340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1645
timestamp 1676037725
transform 1 0 152444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1657
timestamp 1676037725
transform 1 0 153548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1669
timestamp 1676037725
transform 1 0 154652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1677
timestamp 1676037725
transform 1 0 155388 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1681
timestamp 1676037725
transform 1 0 155756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1693
timestamp 1676037725
transform 1 0 156860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1705
timestamp 1676037725
transform 1 0 157964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1717
timestamp 1676037725
transform 1 0 159068 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1729
timestamp 1676037725
transform 1 0 160172 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1735
timestamp 1676037725
transform 1 0 160724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1737
timestamp 1676037725
transform 1 0 160908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1749
timestamp 1676037725
transform 1 0 162012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1761
timestamp 1676037725
transform 1 0 163116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1773
timestamp 1676037725
transform 1 0 164220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1785
timestamp 1676037725
transform 1 0 165324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1791
timestamp 1676037725
transform 1 0 165876 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1793
timestamp 1676037725
transform 1 0 166060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1805
timestamp 1676037725
transform 1 0 167164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1817
timestamp 1676037725
transform 1 0 168268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1829
timestamp 1676037725
transform 1 0 169372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1841
timestamp 1676037725
transform 1 0 170476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1847
timestamp 1676037725
transform 1 0 171028 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1849
timestamp 1676037725
transform 1 0 171212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1861
timestamp 1676037725
transform 1 0 172316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1873
timestamp 1676037725
transform 1 0 173420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1885
timestamp 1676037725
transform 1 0 174524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1897
timestamp 1676037725
transform 1 0 175628 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1903
timestamp 1676037725
transform 1 0 176180 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1905
timestamp 1676037725
transform 1 0 176364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1917
timestamp 1676037725
transform 1 0 177468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1929
timestamp 1676037725
transform 1 0 178572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1941
timestamp 1676037725
transform 1 0 179676 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1953
timestamp 1676037725
transform 1 0 180780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1959
timestamp 1676037725
transform 1 0 181332 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1961
timestamp 1676037725
transform 1 0 181516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1973
timestamp 1676037725
transform 1 0 182620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1985
timestamp 1676037725
transform 1 0 183724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1997
timestamp 1676037725
transform 1 0 184828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2009
timestamp 1676037725
transform 1 0 185932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2015
timestamp 1676037725
transform 1 0 186484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2017
timestamp 1676037725
transform 1 0 186668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2029
timestamp 1676037725
transform 1 0 187772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2041
timestamp 1676037725
transform 1 0 188876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2053
timestamp 1676037725
transform 1 0 189980 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2065
timestamp 1676037725
transform 1 0 191084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2071
timestamp 1676037725
transform 1 0 191636 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2073
timestamp 1676037725
transform 1 0 191820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2085
timestamp 1676037725
transform 1 0 192924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2097
timestamp 1676037725
transform 1 0 194028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2109
timestamp 1676037725
transform 1 0 195132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2121
timestamp 1676037725
transform 1 0 196236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2127
timestamp 1676037725
transform 1 0 196788 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2129
timestamp 1676037725
transform 1 0 196972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2141
timestamp 1676037725
transform 1 0 198076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2153
timestamp 1676037725
transform 1 0 199180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2165
timestamp 1676037725
transform 1 0 200284 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2177
timestamp 1676037725
transform 1 0 201388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2183
timestamp 1676037725
transform 1 0 201940 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2185
timestamp 1676037725
transform 1 0 202124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2197
timestamp 1676037725
transform 1 0 203228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2209
timestamp 1676037725
transform 1 0 204332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2221
timestamp 1676037725
transform 1 0 205436 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2233
timestamp 1676037725
transform 1 0 206540 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2239
timestamp 1676037725
transform 1 0 207092 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2241
timestamp 1676037725
transform 1 0 207276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2253
timestamp 1676037725
transform 1 0 208380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2265
timestamp 1676037725
transform 1 0 209484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2277
timestamp 1676037725
transform 1 0 210588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2289
timestamp 1676037725
transform 1 0 211692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2295
timestamp 1676037725
transform 1 0 212244 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2297
timestamp 1676037725
transform 1 0 212428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2309
timestamp 1676037725
transform 1 0 213532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2321
timestamp 1676037725
transform 1 0 214636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2333
timestamp 1676037725
transform 1 0 215740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2345
timestamp 1676037725
transform 1 0 216844 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2351
timestamp 1676037725
transform 1 0 217396 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2353
timestamp 1676037725
transform 1 0 217580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2365
timestamp 1676037725
transform 1 0 218684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2377
timestamp 1676037725
transform 1 0 219788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2389
timestamp 1676037725
transform 1 0 220892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2401
timestamp 1676037725
transform 1 0 221996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2407
timestamp 1676037725
transform 1 0 222548 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2409
timestamp 1676037725
transform 1 0 222732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2421
timestamp 1676037725
transform 1 0 223836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2433
timestamp 1676037725
transform 1 0 224940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2445
timestamp 1676037725
transform 1 0 226044 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2457
timestamp 1676037725
transform 1 0 227148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2463
timestamp 1676037725
transform 1 0 227700 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2465
timestamp 1676037725
transform 1 0 227884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2477
timestamp 1676037725
transform 1 0 228988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2489
timestamp 1676037725
transform 1 0 230092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2501
timestamp 1676037725
transform 1 0 231196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2513
timestamp 1676037725
transform 1 0 232300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2519
timestamp 1676037725
transform 1 0 232852 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2521
timestamp 1676037725
transform 1 0 233036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2533
timestamp 1676037725
transform 1 0 234140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2545
timestamp 1676037725
transform 1 0 235244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2557
timestamp 1676037725
transform 1 0 236348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2569
timestamp 1676037725
transform 1 0 237452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2575
timestamp 1676037725
transform 1 0 238004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2577
timestamp 1676037725
transform 1 0 238188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2589
timestamp 1676037725
transform 1 0 239292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2601
timestamp 1676037725
transform 1 0 240396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2613
timestamp 1676037725
transform 1 0 241500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2625
timestamp 1676037725
transform 1 0 242604 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2631
timestamp 1676037725
transform 1 0 243156 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2633
timestamp 1676037725
transform 1 0 243340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2645
timestamp 1676037725
transform 1 0 244444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2657
timestamp 1676037725
transform 1 0 245548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2669
timestamp 1676037725
transform 1 0 246652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2681
timestamp 1676037725
transform 1 0 247756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2687
timestamp 1676037725
transform 1 0 248308 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2689
timestamp 1676037725
transform 1 0 248492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2701
timestamp 1676037725
transform 1 0 249596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2713
timestamp 1676037725
transform 1 0 250700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2725
timestamp 1676037725
transform 1 0 251804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2737
timestamp 1676037725
transform 1 0 252908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2743
timestamp 1676037725
transform 1 0 253460 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2745
timestamp 1676037725
transform 1 0 253644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2757
timestamp 1676037725
transform 1 0 254748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2769
timestamp 1676037725
transform 1 0 255852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2781
timestamp 1676037725
transform 1 0 256956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2793
timestamp 1676037725
transform 1 0 258060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2799
timestamp 1676037725
transform 1 0 258612 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2801
timestamp 1676037725
transform 1 0 258796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2813
timestamp 1676037725
transform 1 0 259900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2825
timestamp 1676037725
transform 1 0 261004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2837
timestamp 1676037725
transform 1 0 262108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2849
timestamp 1676037725
transform 1 0 263212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2855
timestamp 1676037725
transform 1 0 263764 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2857
timestamp 1676037725
transform 1 0 263948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2869
timestamp 1676037725
transform 1 0 265052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2881
timestamp 1676037725
transform 1 0 266156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2893
timestamp 1676037725
transform 1 0 267260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2905
timestamp 1676037725
transform 1 0 268364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2911
timestamp 1676037725
transform 1 0 268916 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2913
timestamp 1676037725
transform 1 0 269100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2925
timestamp 1676037725
transform 1 0 270204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2937
timestamp 1676037725
transform 1 0 271308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2949
timestamp 1676037725
transform 1 0 272412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_2961
timestamp 1676037725
transform 1 0 273516 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_2967
timestamp 1676037725
transform 1 0 274068 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2969
timestamp 1676037725
transform 1 0 274252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2981
timestamp 1676037725
transform 1 0 275356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_2993
timestamp 1676037725
transform 1 0 276460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3005
timestamp 1676037725
transform 1 0 277564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3017
timestamp 1676037725
transform 1 0 278668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3023
timestamp 1676037725
transform 1 0 279220 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3025
timestamp 1676037725
transform 1 0 279404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3037
timestamp 1676037725
transform 1 0 280508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3049
timestamp 1676037725
transform 1 0 281612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3061
timestamp 1676037725
transform 1 0 282716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3073
timestamp 1676037725
transform 1 0 283820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3079
timestamp 1676037725
transform 1 0 284372 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3081
timestamp 1676037725
transform 1 0 284556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3093
timestamp 1676037725
transform 1 0 285660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3105
timestamp 1676037725
transform 1 0 286764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3117
timestamp 1676037725
transform 1 0 287868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3129
timestamp 1676037725
transform 1 0 288972 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3135
timestamp 1676037725
transform 1 0 289524 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3137
timestamp 1676037725
transform 1 0 289708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3149
timestamp 1676037725
transform 1 0 290812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3161
timestamp 1676037725
transform 1 0 291916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3173
timestamp 1676037725
transform 1 0 293020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3185
timestamp 1676037725
transform 1 0 294124 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3191
timestamp 1676037725
transform 1 0 294676 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3193
timestamp 1676037725
transform 1 0 294860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3205
timestamp 1676037725
transform 1 0 295964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3217
timestamp 1676037725
transform 1 0 297068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3229
timestamp 1676037725
transform 1 0 298172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3241
timestamp 1676037725
transform 1 0 299276 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3247
timestamp 1676037725
transform 1 0 299828 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3249
timestamp 1676037725
transform 1 0 300012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3261
timestamp 1676037725
transform 1 0 301116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3273
timestamp 1676037725
transform 1 0 302220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3285
timestamp 1676037725
transform 1 0 303324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3297
timestamp 1676037725
transform 1 0 304428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3303
timestamp 1676037725
transform 1 0 304980 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3305
timestamp 1676037725
transform 1 0 305164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3317
timestamp 1676037725
transform 1 0 306268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3329
timestamp 1676037725
transform 1 0 307372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3341
timestamp 1676037725
transform 1 0 308476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3353
timestamp 1676037725
transform 1 0 309580 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3359
timestamp 1676037725
transform 1 0 310132 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3361
timestamp 1676037725
transform 1 0 310316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3373
timestamp 1676037725
transform 1 0 311420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3385
timestamp 1676037725
transform 1 0 312524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3397
timestamp 1676037725
transform 1 0 313628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3409
timestamp 1676037725
transform 1 0 314732 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3415
timestamp 1676037725
transform 1 0 315284 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3417
timestamp 1676037725
transform 1 0 315468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3429
timestamp 1676037725
transform 1 0 316572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3441
timestamp 1676037725
transform 1 0 317676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3453
timestamp 1676037725
transform 1 0 318780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3465
timestamp 1676037725
transform 1 0 319884 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3471
timestamp 1676037725
transform 1 0 320436 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3473
timestamp 1676037725
transform 1 0 320620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3485
timestamp 1676037725
transform 1 0 321724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3497
timestamp 1676037725
transform 1 0 322828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3509
timestamp 1676037725
transform 1 0 323932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3521
timestamp 1676037725
transform 1 0 325036 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3527
timestamp 1676037725
transform 1 0 325588 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3529
timestamp 1676037725
transform 1 0 325772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3541
timestamp 1676037725
transform 1 0 326876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3553
timestamp 1676037725
transform 1 0 327980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3565
timestamp 1676037725
transform 1 0 329084 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3577
timestamp 1676037725
transform 1 0 330188 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3583
timestamp 1676037725
transform 1 0 330740 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3585
timestamp 1676037725
transform 1 0 330924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3597
timestamp 1676037725
transform 1 0 332028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3609
timestamp 1676037725
transform 1 0 333132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3621
timestamp 1676037725
transform 1 0 334236 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3633
timestamp 1676037725
transform 1 0 335340 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3639
timestamp 1676037725
transform 1 0 335892 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3641
timestamp 1676037725
transform 1 0 336076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3653
timestamp 1676037725
transform 1 0 337180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3665
timestamp 1676037725
transform 1 0 338284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3677
timestamp 1676037725
transform 1 0 339388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3689
timestamp 1676037725
transform 1 0 340492 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3695
timestamp 1676037725
transform 1 0 341044 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3697
timestamp 1676037725
transform 1 0 341228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3709
timestamp 1676037725
transform 1 0 342332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3721
timestamp 1676037725
transform 1 0 343436 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3733
timestamp 1676037725
transform 1 0 344540 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3745
timestamp 1676037725
transform 1 0 345644 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3751
timestamp 1676037725
transform 1 0 346196 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3753
timestamp 1676037725
transform 1 0 346380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3765
timestamp 1676037725
transform 1 0 347484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3777
timestamp 1676037725
transform 1 0 348588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3789
timestamp 1676037725
transform 1 0 349692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3801
timestamp 1676037725
transform 1 0 350796 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3807
timestamp 1676037725
transform 1 0 351348 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3809
timestamp 1676037725
transform 1 0 351532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3821
timestamp 1676037725
transform 1 0 352636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3833
timestamp 1676037725
transform 1 0 353740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3845
timestamp 1676037725
transform 1 0 354844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3857
timestamp 1676037725
transform 1 0 355948 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3863
timestamp 1676037725
transform 1 0 356500 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3865
timestamp 1676037725
transform 1 0 356684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3877
timestamp 1676037725
transform 1 0 357788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3889
timestamp 1676037725
transform 1 0 358892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3901
timestamp 1676037725
transform 1 0 359996 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3913
timestamp 1676037725
transform 1 0 361100 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3919
timestamp 1676037725
transform 1 0 361652 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3921
timestamp 1676037725
transform 1 0 361836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3933
timestamp 1676037725
transform 1 0 362940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3945
timestamp 1676037725
transform 1 0 364044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3957
timestamp 1676037725
transform 1 0 365148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3969
timestamp 1676037725
transform 1 0 366252 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3975
timestamp 1676037725
transform 1 0 366804 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3977
timestamp 1676037725
transform 1 0 366988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3989
timestamp 1676037725
transform 1 0 368092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4001
timestamp 1676037725
transform 1 0 369196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4013
timestamp 1676037725
transform 1 0 370300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4025
timestamp 1676037725
transform 1 0 371404 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4031
timestamp 1676037725
transform 1 0 371956 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4033
timestamp 1676037725
transform 1 0 372140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4045
timestamp 1676037725
transform 1 0 373244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4057
timestamp 1676037725
transform 1 0 374348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4069
timestamp 1676037725
transform 1 0 375452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4081
timestamp 1676037725
transform 1 0 376556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4087
timestamp 1676037725
transform 1 0 377108 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4089
timestamp 1676037725
transform 1 0 377292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4101
timestamp 1676037725
transform 1 0 378396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4113
timestamp 1676037725
transform 1 0 379500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4125
timestamp 1676037725
transform 1 0 380604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4137
timestamp 1676037725
transform 1 0 381708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4143
timestamp 1676037725
transform 1 0 382260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4145
timestamp 1676037725
transform 1 0 382444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4157
timestamp 1676037725
transform 1 0 383548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4169
timestamp 1676037725
transform 1 0 384652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4181
timestamp 1676037725
transform 1 0 385756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4193
timestamp 1676037725
transform 1 0 386860 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4199
timestamp 1676037725
transform 1 0 387412 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4201
timestamp 1676037725
transform 1 0 387596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4213
timestamp 1676037725
transform 1 0 388700 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4225
timestamp 1676037725
transform 1 0 389804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4237
timestamp 1676037725
transform 1 0 390908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4249
timestamp 1676037725
transform 1 0 392012 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4255
timestamp 1676037725
transform 1 0 392564 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4257
timestamp 1676037725
transform 1 0 392748 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4269
timestamp 1676037725
transform 1 0 393852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4281
timestamp 1676037725
transform 1 0 394956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4293
timestamp 1676037725
transform 1 0 396060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4305
timestamp 1676037725
transform 1 0 397164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4311
timestamp 1676037725
transform 1 0 397716 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4313
timestamp 1676037725
transform 1 0 397900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4325
timestamp 1676037725
transform 1 0 399004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4337
timestamp 1676037725
transform 1 0 400108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4349
timestamp 1676037725
transform 1 0 401212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4361
timestamp 1676037725
transform 1 0 402316 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4367
timestamp 1676037725
transform 1 0 402868 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4369
timestamp 1676037725
transform 1 0 403052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4381
timestamp 1676037725
transform 1 0 404156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4393
timestamp 1676037725
transform 1 0 405260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4405
timestamp 1676037725
transform 1 0 406364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4417
timestamp 1676037725
transform 1 0 407468 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4423
timestamp 1676037725
transform 1 0 408020 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4425
timestamp 1676037725
transform 1 0 408204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4437
timestamp 1676037725
transform 1 0 409308 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4449
timestamp 1676037725
transform 1 0 410412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4461
timestamp 1676037725
transform 1 0 411516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4473
timestamp 1676037725
transform 1 0 412620 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4479
timestamp 1676037725
transform 1 0 413172 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4481
timestamp 1676037725
transform 1 0 413356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4493
timestamp 1676037725
transform 1 0 414460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4505
timestamp 1676037725
transform 1 0 415564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4517
timestamp 1676037725
transform 1 0 416668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4529
timestamp 1676037725
transform 1 0 417772 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4535
timestamp 1676037725
transform 1 0 418324 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4537
timestamp 1676037725
transform 1 0 418508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4549
timestamp 1676037725
transform 1 0 419612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4561
timestamp 1676037725
transform 1 0 420716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4573
timestamp 1676037725
transform 1 0 421820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4585
timestamp 1676037725
transform 1 0 422924 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4591
timestamp 1676037725
transform 1 0 423476 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4593
timestamp 1676037725
transform 1 0 423660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4605
timestamp 1676037725
transform 1 0 424764 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4617
timestamp 1676037725
transform 1 0 425868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4629
timestamp 1676037725
transform 1 0 426972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4641
timestamp 1676037725
transform 1 0 428076 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4647
timestamp 1676037725
transform 1 0 428628 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4649
timestamp 1676037725
transform 1 0 428812 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4661
timestamp 1676037725
transform 1 0 429916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4673
timestamp 1676037725
transform 1 0 431020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4685
timestamp 1676037725
transform 1 0 432124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4697
timestamp 1676037725
transform 1 0 433228 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4703
timestamp 1676037725
transform 1 0 433780 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4705
timestamp 1676037725
transform 1 0 433964 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4717
timestamp 1676037725
transform 1 0 435068 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4729
timestamp 1676037725
transform 1 0 436172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4741
timestamp 1676037725
transform 1 0 437276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4753
timestamp 1676037725
transform 1 0 438380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4759
timestamp 1676037725
transform 1 0 438932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4761
timestamp 1676037725
transform 1 0 439116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4773
timestamp 1676037725
transform 1 0 440220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4785
timestamp 1676037725
transform 1 0 441324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4797
timestamp 1676037725
transform 1 0 442428 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4809
timestamp 1676037725
transform 1 0 443532 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4815
timestamp 1676037725
transform 1 0 444084 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4817
timestamp 1676037725
transform 1 0 444268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4829
timestamp 1676037725
transform 1 0 445372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4841
timestamp 1676037725
transform 1 0 446476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4853
timestamp 1676037725
transform 1 0 447580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4865
timestamp 1676037725
transform 1 0 448684 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4871
timestamp 1676037725
transform 1 0 449236 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4873
timestamp 1676037725
transform 1 0 449420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4885
timestamp 1676037725
transform 1 0 450524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4897
timestamp 1676037725
transform 1 0 451628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4909
timestamp 1676037725
transform 1 0 452732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4921
timestamp 1676037725
transform 1 0 453836 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4927
timestamp 1676037725
transform 1 0 454388 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4929
timestamp 1676037725
transform 1 0 454572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4941
timestamp 1676037725
transform 1 0 455676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4953
timestamp 1676037725
transform 1 0 456780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4965
timestamp 1676037725
transform 1 0 457884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_4977
timestamp 1676037725
transform 1 0 458988 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_4983
timestamp 1676037725
transform 1 0 459540 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4985
timestamp 1676037725
transform 1 0 459724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_4997
timestamp 1676037725
transform 1 0 460828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5009
timestamp 1676037725
transform 1 0 461932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5021
timestamp 1676037725
transform 1 0 463036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5033
timestamp 1676037725
transform 1 0 464140 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5039
timestamp 1676037725
transform 1 0 464692 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5041
timestamp 1676037725
transform 1 0 464876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5053
timestamp 1676037725
transform 1 0 465980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5065
timestamp 1676037725
transform 1 0 467084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5077
timestamp 1676037725
transform 1 0 468188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5089
timestamp 1676037725
transform 1 0 469292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5095
timestamp 1676037725
transform 1 0 469844 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5097
timestamp 1676037725
transform 1 0 470028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5109
timestamp 1676037725
transform 1 0 471132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5121
timestamp 1676037725
transform 1 0 472236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5133
timestamp 1676037725
transform 1 0 473340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5145
timestamp 1676037725
transform 1 0 474444 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5151
timestamp 1676037725
transform 1 0 474996 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5153
timestamp 1676037725
transform 1 0 475180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5165
timestamp 1676037725
transform 1 0 476284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5177
timestamp 1676037725
transform 1 0 477388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5189
timestamp 1676037725
transform 1 0 478492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5201
timestamp 1676037725
transform 1 0 479596 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5207
timestamp 1676037725
transform 1 0 480148 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5209
timestamp 1676037725
transform 1 0 480332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5221
timestamp 1676037725
transform 1 0 481436 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5233
timestamp 1676037725
transform 1 0 482540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5245
timestamp 1676037725
transform 1 0 483644 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5257
timestamp 1676037725
transform 1 0 484748 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5263
timestamp 1676037725
transform 1 0 485300 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5265
timestamp 1676037725
transform 1 0 485484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5277
timestamp 1676037725
transform 1 0 486588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5289
timestamp 1676037725
transform 1 0 487692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5301
timestamp 1676037725
transform 1 0 488796 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5313
timestamp 1676037725
transform 1 0 489900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5319
timestamp 1676037725
transform 1 0 490452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5321
timestamp 1676037725
transform 1 0 490636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5333
timestamp 1676037725
transform 1 0 491740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5345
timestamp 1676037725
transform 1 0 492844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5357
timestamp 1676037725
transform 1 0 493948 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5369
timestamp 1676037725
transform 1 0 495052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5375
timestamp 1676037725
transform 1 0 495604 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5377
timestamp 1676037725
transform 1 0 495788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5389
timestamp 1676037725
transform 1 0 496892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5401
timestamp 1676037725
transform 1 0 497996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5413
timestamp 1676037725
transform 1 0 499100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5425
timestamp 1676037725
transform 1 0 500204 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5431
timestamp 1676037725
transform 1 0 500756 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5433
timestamp 1676037725
transform 1 0 500940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5445
timestamp 1676037725
transform 1 0 502044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5457
timestamp 1676037725
transform 1 0 503148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5469
timestamp 1676037725
transform 1 0 504252 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5481
timestamp 1676037725
transform 1 0 505356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5487
timestamp 1676037725
transform 1 0 505908 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5489
timestamp 1676037725
transform 1 0 506092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5501
timestamp 1676037725
transform 1 0 507196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5513
timestamp 1676037725
transform 1 0 508300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5525
timestamp 1676037725
transform 1 0 509404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5537
timestamp 1676037725
transform 1 0 510508 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5543
timestamp 1676037725
transform 1 0 511060 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5545
timestamp 1676037725
transform 1 0 511244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5557
timestamp 1676037725
transform 1 0 512348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5569
timestamp 1676037725
transform 1 0 513452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5581
timestamp 1676037725
transform 1 0 514556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5593
timestamp 1676037725
transform 1 0 515660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5599
timestamp 1676037725
transform 1 0 516212 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5601
timestamp 1676037725
transform 1 0 516396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5613
timestamp 1676037725
transform 1 0 517500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5625
timestamp 1676037725
transform 1 0 518604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5637
timestamp 1676037725
transform 1 0 519708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5649
timestamp 1676037725
transform 1 0 520812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5655
timestamp 1676037725
transform 1 0 521364 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5657
timestamp 1676037725
transform 1 0 521548 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5669
timestamp 1676037725
transform 1 0 522652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5681
timestamp 1676037725
transform 1 0 523756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5693
timestamp 1676037725
transform 1 0 524860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_5705
timestamp 1676037725
transform 1 0 525964 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_5711
timestamp 1676037725
transform 1 0 526516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5713
timestamp 1676037725
transform 1 0 526700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_5725
timestamp 1676037725
transform 1 0 527804 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1676037725
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1676037725
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1676037725
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1676037725
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1676037725
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1676037725
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1676037725
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1676037725
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1676037725
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1676037725
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1676037725
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1676037725
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1676037725
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1676037725
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1676037725
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1676037725
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1676037725
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1676037725
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1676037725
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1676037725
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1676037725
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1676037725
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1676037725
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1676037725
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1676037725
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1676037725
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1676037725
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1676037725
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1676037725
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1676037725
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1676037725
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1676037725
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1676037725
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1676037725
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1676037725
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1676037725
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1676037725
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1676037725
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1676037725
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1676037725
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1676037725
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1676037725
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1676037725
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1676037725
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1676037725
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1676037725
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1676037725
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1676037725
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1676037725
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1676037725
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1676037725
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1676037725
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1676037725
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1676037725
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1676037725
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1676037725
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1676037725
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1676037725
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1676037725
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1676037725
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1676037725
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1676037725
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1676037725
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1676037725
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1676037725
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1676037725
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1676037725
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1676037725
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1676037725
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1217
timestamp 1676037725
transform 1 0 113068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1229
timestamp 1676037725
transform 1 0 114172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1241
timestamp 1676037725
transform 1 0 115276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1253
timestamp 1676037725
transform 1 0 116380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1676037725
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1261
timestamp 1676037725
transform 1 0 117116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1273
timestamp 1676037725
transform 1 0 118220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1285
timestamp 1676037725
transform 1 0 119324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1297
timestamp 1676037725
transform 1 0 120428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1309
timestamp 1676037725
transform 1 0 121532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1315
timestamp 1676037725
transform 1 0 122084 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1317
timestamp 1676037725
transform 1 0 122268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1329
timestamp 1676037725
transform 1 0 123372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1341
timestamp 1676037725
transform 1 0 124476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1353
timestamp 1676037725
transform 1 0 125580 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1365
timestamp 1676037725
transform 1 0 126684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1371
timestamp 1676037725
transform 1 0 127236 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1373
timestamp 1676037725
transform 1 0 127420 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1377
timestamp 1676037725
transform 1 0 127788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1389
timestamp 1676037725
transform 1 0 128892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1401
timestamp 1676037725
transform 1 0 129996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1413
timestamp 1676037725
transform 1 0 131100 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1416
timestamp 1676037725
transform 1 0 131376 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1429
timestamp 1676037725
transform 1 0 132572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1441
timestamp 1676037725
transform 1 0 133676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1445
timestamp 1676037725
transform 1 0 134044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1448
timestamp 1676037725
transform 1 0 134320 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1460
timestamp 1676037725
transform 1 0 135424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1470
timestamp 1676037725
transform 1 0 136344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1480
timestamp 1676037725
transform 1 0 137264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1485
timestamp 1676037725
transform 1 0 137724 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1493
timestamp 1676037725
transform 1 0 138460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1505
timestamp 1676037725
transform 1 0 139564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1508
timestamp 1676037725
transform 1 0 139840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1518
timestamp 1676037725
transform 1 0 140760 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1530
timestamp 1676037725
transform 1 0 141864 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1538
timestamp 1676037725
transform 1 0 142600 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1541
timestamp 1676037725
transform 1 0 142876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1553
timestamp 1676037725
transform 1 0 143980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1565
timestamp 1676037725
transform 1 0 145084 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1571
timestamp 1676037725
transform 1 0 145636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1583
timestamp 1676037725
transform 1 0 146740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1595
timestamp 1676037725
transform 1 0 147844 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1597
timestamp 1676037725
transform 1 0 148028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1615
timestamp 1676037725
transform 1 0 149684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1627
timestamp 1676037725
transform 1 0 150788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1639
timestamp 1676037725
transform 1 0 151892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1651
timestamp 1676037725
transform 1 0 152996 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1653
timestamp 1676037725
transform 1 0 153180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1665
timestamp 1676037725
transform 1 0 154284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1677
timestamp 1676037725
transform 1 0 155388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1689
timestamp 1676037725
transform 1 0 156492 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1701
timestamp 1676037725
transform 1 0 157596 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1707
timestamp 1676037725
transform 1 0 158148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1709
timestamp 1676037725
transform 1 0 158332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1721
timestamp 1676037725
transform 1 0 159436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1733
timestamp 1676037725
transform 1 0 160540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1745
timestamp 1676037725
transform 1 0 161644 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1757
timestamp 1676037725
transform 1 0 162748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1763
timestamp 1676037725
transform 1 0 163300 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1765
timestamp 1676037725
transform 1 0 163484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1777
timestamp 1676037725
transform 1 0 164588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1789
timestamp 1676037725
transform 1 0 165692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1801
timestamp 1676037725
transform 1 0 166796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1813
timestamp 1676037725
transform 1 0 167900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1819
timestamp 1676037725
transform 1 0 168452 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1821
timestamp 1676037725
transform 1 0 168636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1833
timestamp 1676037725
transform 1 0 169740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1845
timestamp 1676037725
transform 1 0 170844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1857
timestamp 1676037725
transform 1 0 171948 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1869
timestamp 1676037725
transform 1 0 173052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1875
timestamp 1676037725
transform 1 0 173604 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1877
timestamp 1676037725
transform 1 0 173788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1889
timestamp 1676037725
transform 1 0 174892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1901
timestamp 1676037725
transform 1 0 175996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1913
timestamp 1676037725
transform 1 0 177100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1925
timestamp 1676037725
transform 1 0 178204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1931
timestamp 1676037725
transform 1 0 178756 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1933
timestamp 1676037725
transform 1 0 178940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1945
timestamp 1676037725
transform 1 0 180044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1957
timestamp 1676037725
transform 1 0 181148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1969
timestamp 1676037725
transform 1 0 182252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1981
timestamp 1676037725
transform 1 0 183356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1987
timestamp 1676037725
transform 1 0 183908 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1989
timestamp 1676037725
transform 1 0 184092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2001
timestamp 1676037725
transform 1 0 185196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2013
timestamp 1676037725
transform 1 0 186300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2025
timestamp 1676037725
transform 1 0 187404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2037
timestamp 1676037725
transform 1 0 188508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2043
timestamp 1676037725
transform 1 0 189060 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2045
timestamp 1676037725
transform 1 0 189244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2057
timestamp 1676037725
transform 1 0 190348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2069
timestamp 1676037725
transform 1 0 191452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2081
timestamp 1676037725
transform 1 0 192556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2093
timestamp 1676037725
transform 1 0 193660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2099
timestamp 1676037725
transform 1 0 194212 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2101
timestamp 1676037725
transform 1 0 194396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2113
timestamp 1676037725
transform 1 0 195500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2125
timestamp 1676037725
transform 1 0 196604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2137
timestamp 1676037725
transform 1 0 197708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2149
timestamp 1676037725
transform 1 0 198812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2155
timestamp 1676037725
transform 1 0 199364 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2157
timestamp 1676037725
transform 1 0 199548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2169
timestamp 1676037725
transform 1 0 200652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2181
timestamp 1676037725
transform 1 0 201756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2193
timestamp 1676037725
transform 1 0 202860 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2205
timestamp 1676037725
transform 1 0 203964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2211
timestamp 1676037725
transform 1 0 204516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2213
timestamp 1676037725
transform 1 0 204700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2225
timestamp 1676037725
transform 1 0 205804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2237
timestamp 1676037725
transform 1 0 206908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2249
timestamp 1676037725
transform 1 0 208012 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2261
timestamp 1676037725
transform 1 0 209116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2267
timestamp 1676037725
transform 1 0 209668 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2269
timestamp 1676037725
transform 1 0 209852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2281
timestamp 1676037725
transform 1 0 210956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2293
timestamp 1676037725
transform 1 0 212060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2305
timestamp 1676037725
transform 1 0 213164 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2317
timestamp 1676037725
transform 1 0 214268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2323
timestamp 1676037725
transform 1 0 214820 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2325
timestamp 1676037725
transform 1 0 215004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2337
timestamp 1676037725
transform 1 0 216108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2349
timestamp 1676037725
transform 1 0 217212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2361
timestamp 1676037725
transform 1 0 218316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2373
timestamp 1676037725
transform 1 0 219420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2379
timestamp 1676037725
transform 1 0 219972 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2381
timestamp 1676037725
transform 1 0 220156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2393
timestamp 1676037725
transform 1 0 221260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2405
timestamp 1676037725
transform 1 0 222364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2417
timestamp 1676037725
transform 1 0 223468 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2429
timestamp 1676037725
transform 1 0 224572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2435
timestamp 1676037725
transform 1 0 225124 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2437
timestamp 1676037725
transform 1 0 225308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2449
timestamp 1676037725
transform 1 0 226412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2461
timestamp 1676037725
transform 1 0 227516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2473
timestamp 1676037725
transform 1 0 228620 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2485
timestamp 1676037725
transform 1 0 229724 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2491
timestamp 1676037725
transform 1 0 230276 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2493
timestamp 1676037725
transform 1 0 230460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2505
timestamp 1676037725
transform 1 0 231564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2517
timestamp 1676037725
transform 1 0 232668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2529
timestamp 1676037725
transform 1 0 233772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2541
timestamp 1676037725
transform 1 0 234876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2547
timestamp 1676037725
transform 1 0 235428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2549
timestamp 1676037725
transform 1 0 235612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2561
timestamp 1676037725
transform 1 0 236716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2573
timestamp 1676037725
transform 1 0 237820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2585
timestamp 1676037725
transform 1 0 238924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2597
timestamp 1676037725
transform 1 0 240028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2603
timestamp 1676037725
transform 1 0 240580 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2605
timestamp 1676037725
transform 1 0 240764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2617
timestamp 1676037725
transform 1 0 241868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2629
timestamp 1676037725
transform 1 0 242972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2641
timestamp 1676037725
transform 1 0 244076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2653
timestamp 1676037725
transform 1 0 245180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2659
timestamp 1676037725
transform 1 0 245732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2661
timestamp 1676037725
transform 1 0 245916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2673
timestamp 1676037725
transform 1 0 247020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2685
timestamp 1676037725
transform 1 0 248124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2697
timestamp 1676037725
transform 1 0 249228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2709
timestamp 1676037725
transform 1 0 250332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2715
timestamp 1676037725
transform 1 0 250884 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2717
timestamp 1676037725
transform 1 0 251068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2729
timestamp 1676037725
transform 1 0 252172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2741
timestamp 1676037725
transform 1 0 253276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2753
timestamp 1676037725
transform 1 0 254380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2765
timestamp 1676037725
transform 1 0 255484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2771
timestamp 1676037725
transform 1 0 256036 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2773
timestamp 1676037725
transform 1 0 256220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2785
timestamp 1676037725
transform 1 0 257324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2797
timestamp 1676037725
transform 1 0 258428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2809
timestamp 1676037725
transform 1 0 259532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2821
timestamp 1676037725
transform 1 0 260636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2827
timestamp 1676037725
transform 1 0 261188 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2829
timestamp 1676037725
transform 1 0 261372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2841
timestamp 1676037725
transform 1 0 262476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2853
timestamp 1676037725
transform 1 0 263580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2865
timestamp 1676037725
transform 1 0 264684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2877
timestamp 1676037725
transform 1 0 265788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2883
timestamp 1676037725
transform 1 0 266340 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2885
timestamp 1676037725
transform 1 0 266524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2897
timestamp 1676037725
transform 1 0 267628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2909
timestamp 1676037725
transform 1 0 268732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2921
timestamp 1676037725
transform 1 0 269836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2933
timestamp 1676037725
transform 1 0 270940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2939
timestamp 1676037725
transform 1 0 271492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2941
timestamp 1676037725
transform 1 0 271676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2953
timestamp 1676037725
transform 1 0 272780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2965
timestamp 1676037725
transform 1 0 273884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2977
timestamp 1676037725
transform 1 0 274988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_2989
timestamp 1676037725
transform 1 0 276092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_2995
timestamp 1676037725
transform 1 0 276644 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_2997
timestamp 1676037725
transform 1 0 276828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3009
timestamp 1676037725
transform 1 0 277932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3021
timestamp 1676037725
transform 1 0 279036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3033
timestamp 1676037725
transform 1 0 280140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3045
timestamp 1676037725
transform 1 0 281244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3051
timestamp 1676037725
transform 1 0 281796 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3053
timestamp 1676037725
transform 1 0 281980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3065
timestamp 1676037725
transform 1 0 283084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3077
timestamp 1676037725
transform 1 0 284188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3089
timestamp 1676037725
transform 1 0 285292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3101
timestamp 1676037725
transform 1 0 286396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3107
timestamp 1676037725
transform 1 0 286948 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3109
timestamp 1676037725
transform 1 0 287132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3121
timestamp 1676037725
transform 1 0 288236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3133
timestamp 1676037725
transform 1 0 289340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3145
timestamp 1676037725
transform 1 0 290444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3157
timestamp 1676037725
transform 1 0 291548 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3163
timestamp 1676037725
transform 1 0 292100 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3165
timestamp 1676037725
transform 1 0 292284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3177
timestamp 1676037725
transform 1 0 293388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3189
timestamp 1676037725
transform 1 0 294492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3201
timestamp 1676037725
transform 1 0 295596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3213
timestamp 1676037725
transform 1 0 296700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3219
timestamp 1676037725
transform 1 0 297252 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3221
timestamp 1676037725
transform 1 0 297436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3233
timestamp 1676037725
transform 1 0 298540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3245
timestamp 1676037725
transform 1 0 299644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3257
timestamp 1676037725
transform 1 0 300748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3269
timestamp 1676037725
transform 1 0 301852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3275
timestamp 1676037725
transform 1 0 302404 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3277
timestamp 1676037725
transform 1 0 302588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3289
timestamp 1676037725
transform 1 0 303692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3301
timestamp 1676037725
transform 1 0 304796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3313
timestamp 1676037725
transform 1 0 305900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3325
timestamp 1676037725
transform 1 0 307004 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3331
timestamp 1676037725
transform 1 0 307556 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3333
timestamp 1676037725
transform 1 0 307740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3345
timestamp 1676037725
transform 1 0 308844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3357
timestamp 1676037725
transform 1 0 309948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3369
timestamp 1676037725
transform 1 0 311052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3381
timestamp 1676037725
transform 1 0 312156 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3387
timestamp 1676037725
transform 1 0 312708 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3389
timestamp 1676037725
transform 1 0 312892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3401
timestamp 1676037725
transform 1 0 313996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3413
timestamp 1676037725
transform 1 0 315100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3425
timestamp 1676037725
transform 1 0 316204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3437
timestamp 1676037725
transform 1 0 317308 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3443
timestamp 1676037725
transform 1 0 317860 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3445
timestamp 1676037725
transform 1 0 318044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3457
timestamp 1676037725
transform 1 0 319148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3469
timestamp 1676037725
transform 1 0 320252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3481
timestamp 1676037725
transform 1 0 321356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3493
timestamp 1676037725
transform 1 0 322460 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3499
timestamp 1676037725
transform 1 0 323012 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3501
timestamp 1676037725
transform 1 0 323196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3513
timestamp 1676037725
transform 1 0 324300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3525
timestamp 1676037725
transform 1 0 325404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3537
timestamp 1676037725
transform 1 0 326508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3549
timestamp 1676037725
transform 1 0 327612 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3555
timestamp 1676037725
transform 1 0 328164 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3557
timestamp 1676037725
transform 1 0 328348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3569
timestamp 1676037725
transform 1 0 329452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3581
timestamp 1676037725
transform 1 0 330556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3593
timestamp 1676037725
transform 1 0 331660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3605
timestamp 1676037725
transform 1 0 332764 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3611
timestamp 1676037725
transform 1 0 333316 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3613
timestamp 1676037725
transform 1 0 333500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3625
timestamp 1676037725
transform 1 0 334604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3637
timestamp 1676037725
transform 1 0 335708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3649
timestamp 1676037725
transform 1 0 336812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3661
timestamp 1676037725
transform 1 0 337916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3667
timestamp 1676037725
transform 1 0 338468 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3669
timestamp 1676037725
transform 1 0 338652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3681
timestamp 1676037725
transform 1 0 339756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3693
timestamp 1676037725
transform 1 0 340860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3705
timestamp 1676037725
transform 1 0 341964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3717
timestamp 1676037725
transform 1 0 343068 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3723
timestamp 1676037725
transform 1 0 343620 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3725
timestamp 1676037725
transform 1 0 343804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3737
timestamp 1676037725
transform 1 0 344908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3749
timestamp 1676037725
transform 1 0 346012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3761
timestamp 1676037725
transform 1 0 347116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3773
timestamp 1676037725
transform 1 0 348220 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3779
timestamp 1676037725
transform 1 0 348772 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3781
timestamp 1676037725
transform 1 0 348956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3793
timestamp 1676037725
transform 1 0 350060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3805
timestamp 1676037725
transform 1 0 351164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3817
timestamp 1676037725
transform 1 0 352268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3829
timestamp 1676037725
transform 1 0 353372 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3835
timestamp 1676037725
transform 1 0 353924 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3837
timestamp 1676037725
transform 1 0 354108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3849
timestamp 1676037725
transform 1 0 355212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3861
timestamp 1676037725
transform 1 0 356316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3873
timestamp 1676037725
transform 1 0 357420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3885
timestamp 1676037725
transform 1 0 358524 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3891
timestamp 1676037725
transform 1 0 359076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3893
timestamp 1676037725
transform 1 0 359260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3905
timestamp 1676037725
transform 1 0 360364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3917
timestamp 1676037725
transform 1 0 361468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3929
timestamp 1676037725
transform 1 0 362572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3941
timestamp 1676037725
transform 1 0 363676 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3947
timestamp 1676037725
transform 1 0 364228 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3949
timestamp 1676037725
transform 1 0 364412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3961
timestamp 1676037725
transform 1 0 365516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3973
timestamp 1676037725
transform 1 0 366620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3985
timestamp 1676037725
transform 1 0 367724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3997
timestamp 1676037725
transform 1 0 368828 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4003
timestamp 1676037725
transform 1 0 369380 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4005
timestamp 1676037725
transform 1 0 369564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4017
timestamp 1676037725
transform 1 0 370668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4029
timestamp 1676037725
transform 1 0 371772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4041
timestamp 1676037725
transform 1 0 372876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4053
timestamp 1676037725
transform 1 0 373980 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4059
timestamp 1676037725
transform 1 0 374532 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4061
timestamp 1676037725
transform 1 0 374716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4073
timestamp 1676037725
transform 1 0 375820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4085
timestamp 1676037725
transform 1 0 376924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4097
timestamp 1676037725
transform 1 0 378028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4109
timestamp 1676037725
transform 1 0 379132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4115
timestamp 1676037725
transform 1 0 379684 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4117
timestamp 1676037725
transform 1 0 379868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4129
timestamp 1676037725
transform 1 0 380972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4141
timestamp 1676037725
transform 1 0 382076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4153
timestamp 1676037725
transform 1 0 383180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4165
timestamp 1676037725
transform 1 0 384284 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4171
timestamp 1676037725
transform 1 0 384836 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4173
timestamp 1676037725
transform 1 0 385020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4185
timestamp 1676037725
transform 1 0 386124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4197
timestamp 1676037725
transform 1 0 387228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4209
timestamp 1676037725
transform 1 0 388332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4221
timestamp 1676037725
transform 1 0 389436 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4227
timestamp 1676037725
transform 1 0 389988 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4229
timestamp 1676037725
transform 1 0 390172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4241
timestamp 1676037725
transform 1 0 391276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4253
timestamp 1676037725
transform 1 0 392380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4265
timestamp 1676037725
transform 1 0 393484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4277
timestamp 1676037725
transform 1 0 394588 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4283
timestamp 1676037725
transform 1 0 395140 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4285
timestamp 1676037725
transform 1 0 395324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4297
timestamp 1676037725
transform 1 0 396428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4309
timestamp 1676037725
transform 1 0 397532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4321
timestamp 1676037725
transform 1 0 398636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4333
timestamp 1676037725
transform 1 0 399740 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4339
timestamp 1676037725
transform 1 0 400292 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4341
timestamp 1676037725
transform 1 0 400476 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4353
timestamp 1676037725
transform 1 0 401580 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4365
timestamp 1676037725
transform 1 0 402684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4377
timestamp 1676037725
transform 1 0 403788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4389
timestamp 1676037725
transform 1 0 404892 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4395
timestamp 1676037725
transform 1 0 405444 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4397
timestamp 1676037725
transform 1 0 405628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4409
timestamp 1676037725
transform 1 0 406732 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4421
timestamp 1676037725
transform 1 0 407836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4433
timestamp 1676037725
transform 1 0 408940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4445
timestamp 1676037725
transform 1 0 410044 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4451
timestamp 1676037725
transform 1 0 410596 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4453
timestamp 1676037725
transform 1 0 410780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4465
timestamp 1676037725
transform 1 0 411884 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4477
timestamp 1676037725
transform 1 0 412988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4489
timestamp 1676037725
transform 1 0 414092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4501
timestamp 1676037725
transform 1 0 415196 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4507
timestamp 1676037725
transform 1 0 415748 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4509
timestamp 1676037725
transform 1 0 415932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4521
timestamp 1676037725
transform 1 0 417036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4533
timestamp 1676037725
transform 1 0 418140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4545
timestamp 1676037725
transform 1 0 419244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4557
timestamp 1676037725
transform 1 0 420348 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4563
timestamp 1676037725
transform 1 0 420900 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4565
timestamp 1676037725
transform 1 0 421084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4577
timestamp 1676037725
transform 1 0 422188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4589
timestamp 1676037725
transform 1 0 423292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4601
timestamp 1676037725
transform 1 0 424396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4613
timestamp 1676037725
transform 1 0 425500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4619
timestamp 1676037725
transform 1 0 426052 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4621
timestamp 1676037725
transform 1 0 426236 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4633
timestamp 1676037725
transform 1 0 427340 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4645
timestamp 1676037725
transform 1 0 428444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4657
timestamp 1676037725
transform 1 0 429548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4669
timestamp 1676037725
transform 1 0 430652 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4675
timestamp 1676037725
transform 1 0 431204 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4677
timestamp 1676037725
transform 1 0 431388 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4689
timestamp 1676037725
transform 1 0 432492 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4701
timestamp 1676037725
transform 1 0 433596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4713
timestamp 1676037725
transform 1 0 434700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4725
timestamp 1676037725
transform 1 0 435804 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4731
timestamp 1676037725
transform 1 0 436356 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4733
timestamp 1676037725
transform 1 0 436540 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4745
timestamp 1676037725
transform 1 0 437644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4757
timestamp 1676037725
transform 1 0 438748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4769
timestamp 1676037725
transform 1 0 439852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4781
timestamp 1676037725
transform 1 0 440956 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4787
timestamp 1676037725
transform 1 0 441508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4789
timestamp 1676037725
transform 1 0 441692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4801
timestamp 1676037725
transform 1 0 442796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4813
timestamp 1676037725
transform 1 0 443900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4825
timestamp 1676037725
transform 1 0 445004 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4837
timestamp 1676037725
transform 1 0 446108 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4843
timestamp 1676037725
transform 1 0 446660 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4845
timestamp 1676037725
transform 1 0 446844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4857
timestamp 1676037725
transform 1 0 447948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4869
timestamp 1676037725
transform 1 0 449052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4881
timestamp 1676037725
transform 1 0 450156 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4893
timestamp 1676037725
transform 1 0 451260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4899
timestamp 1676037725
transform 1 0 451812 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4901
timestamp 1676037725
transform 1 0 451996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4913
timestamp 1676037725
transform 1 0 453100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4925
timestamp 1676037725
transform 1 0 454204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4937
timestamp 1676037725
transform 1 0 455308 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_4949
timestamp 1676037725
transform 1 0 456412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_4955
timestamp 1676037725
transform 1 0 456964 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4957
timestamp 1676037725
transform 1 0 457148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4969
timestamp 1676037725
transform 1 0 458252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4981
timestamp 1676037725
transform 1 0 459356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_4993
timestamp 1676037725
transform 1 0 460460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5005
timestamp 1676037725
transform 1 0 461564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5011
timestamp 1676037725
transform 1 0 462116 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5013
timestamp 1676037725
transform 1 0 462300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5025
timestamp 1676037725
transform 1 0 463404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5037
timestamp 1676037725
transform 1 0 464508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5049
timestamp 1676037725
transform 1 0 465612 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5061
timestamp 1676037725
transform 1 0 466716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5067
timestamp 1676037725
transform 1 0 467268 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5069
timestamp 1676037725
transform 1 0 467452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5081
timestamp 1676037725
transform 1 0 468556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5093
timestamp 1676037725
transform 1 0 469660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5105
timestamp 1676037725
transform 1 0 470764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5117
timestamp 1676037725
transform 1 0 471868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5123
timestamp 1676037725
transform 1 0 472420 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5125
timestamp 1676037725
transform 1 0 472604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5137
timestamp 1676037725
transform 1 0 473708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5149
timestamp 1676037725
transform 1 0 474812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5161
timestamp 1676037725
transform 1 0 475916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5173
timestamp 1676037725
transform 1 0 477020 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5179
timestamp 1676037725
transform 1 0 477572 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5181
timestamp 1676037725
transform 1 0 477756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5193
timestamp 1676037725
transform 1 0 478860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5205
timestamp 1676037725
transform 1 0 479964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5217
timestamp 1676037725
transform 1 0 481068 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5229
timestamp 1676037725
transform 1 0 482172 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5235
timestamp 1676037725
transform 1 0 482724 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5237
timestamp 1676037725
transform 1 0 482908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5249
timestamp 1676037725
transform 1 0 484012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5261
timestamp 1676037725
transform 1 0 485116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5273
timestamp 1676037725
transform 1 0 486220 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5285
timestamp 1676037725
transform 1 0 487324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5291
timestamp 1676037725
transform 1 0 487876 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5293
timestamp 1676037725
transform 1 0 488060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5305
timestamp 1676037725
transform 1 0 489164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5317
timestamp 1676037725
transform 1 0 490268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5329
timestamp 1676037725
transform 1 0 491372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5341
timestamp 1676037725
transform 1 0 492476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5347
timestamp 1676037725
transform 1 0 493028 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5349
timestamp 1676037725
transform 1 0 493212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5361
timestamp 1676037725
transform 1 0 494316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5373
timestamp 1676037725
transform 1 0 495420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5385
timestamp 1676037725
transform 1 0 496524 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5397
timestamp 1676037725
transform 1 0 497628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5403
timestamp 1676037725
transform 1 0 498180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5405
timestamp 1676037725
transform 1 0 498364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5417
timestamp 1676037725
transform 1 0 499468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5429
timestamp 1676037725
transform 1 0 500572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5441
timestamp 1676037725
transform 1 0 501676 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5453
timestamp 1676037725
transform 1 0 502780 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5459
timestamp 1676037725
transform 1 0 503332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5461
timestamp 1676037725
transform 1 0 503516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5473
timestamp 1676037725
transform 1 0 504620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5485
timestamp 1676037725
transform 1 0 505724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5497
timestamp 1676037725
transform 1 0 506828 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5509
timestamp 1676037725
transform 1 0 507932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5515
timestamp 1676037725
transform 1 0 508484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5517
timestamp 1676037725
transform 1 0 508668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5529
timestamp 1676037725
transform 1 0 509772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5541
timestamp 1676037725
transform 1 0 510876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5553
timestamp 1676037725
transform 1 0 511980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5565
timestamp 1676037725
transform 1 0 513084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5571
timestamp 1676037725
transform 1 0 513636 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5573
timestamp 1676037725
transform 1 0 513820 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5585
timestamp 1676037725
transform 1 0 514924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5597
timestamp 1676037725
transform 1 0 516028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5609
timestamp 1676037725
transform 1 0 517132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5621
timestamp 1676037725
transform 1 0 518236 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5627
timestamp 1676037725
transform 1 0 518788 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5629
timestamp 1676037725
transform 1 0 518972 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5641
timestamp 1676037725
transform 1 0 520076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5653
timestamp 1676037725
transform 1 0 521180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5665
timestamp 1676037725
transform 1 0 522284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_5677
timestamp 1676037725
transform 1 0 523388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_5683
timestamp 1676037725
transform 1 0 523940 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5685
timestamp 1676037725
transform 1 0 524124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5697
timestamp 1676037725
transform 1 0 525228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5709
timestamp 1676037725
transform 1 0 526332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5721
timestamp 1676037725
transform 1 0 527436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1676037725
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1676037725
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1676037725
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1676037725
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1676037725
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1676037725
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1676037725
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1676037725
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1676037725
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1676037725
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1676037725
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1676037725
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1676037725
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1676037725
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1676037725
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1676037725
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1676037725
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1676037725
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1676037725
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1676037725
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1676037725
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1676037725
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1676037725
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1676037725
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1676037725
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1676037725
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1676037725
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1676037725
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1676037725
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1676037725
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1676037725
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1676037725
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1676037725
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1676037725
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1676037725
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1676037725
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1676037725
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1676037725
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1676037725
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1676037725
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1676037725
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1676037725
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1676037725
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1676037725
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1676037725
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1676037725
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1676037725
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1676037725
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1676037725
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1676037725
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1676037725
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1676037725
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1676037725
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1676037725
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1676037725
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1676037725
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1676037725
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1676037725
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1676037725
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1676037725
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1676037725
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1676037725
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1676037725
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1676037725
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1676037725
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1676037725
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1676037725
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1676037725
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1676037725
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1676037725
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1676037725
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1676037725
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1676037725
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1245
timestamp 1676037725
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1257
timestamp 1676037725
transform 1 0 116748 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1263
timestamp 1676037725
transform 1 0 117300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1275
timestamp 1676037725
transform 1 0 118404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1287
timestamp 1676037725
transform 1 0 119508 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1289
timestamp 1676037725
transform 1 0 119692 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1299
timestamp 1676037725
transform 1 0 120612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1311
timestamp 1676037725
transform 1 0 121716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1319
timestamp 1676037725
transform 1 0 122452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1323
timestamp 1676037725
transform 1 0 122820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1331
timestamp 1676037725
transform 1 0 123556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1336
timestamp 1676037725
transform 1 0 124016 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1345
timestamp 1676037725
transform 1 0 124844 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1353
timestamp 1676037725
transform 1 0 125580 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1356
timestamp 1676037725
transform 1 0 125856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1369
timestamp 1676037725
transform 1 0 127052 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1382
timestamp 1676037725
transform 1 0 128248 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1394
timestamp 1676037725
transform 1 0 129352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1398
timestamp 1676037725
transform 1 0 129720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1401
timestamp 1676037725
transform 1 0 129996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1412
timestamp 1676037725
transform 1 0 131008 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1422
timestamp 1676037725
transform 1 0 131928 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1432
timestamp 1676037725
transform 1 0 132848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1442
timestamp 1676037725
transform 1 0 133768 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1454
timestamp 1676037725
transform 1 0 134872 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1457
timestamp 1676037725
transform 1 0 135148 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1461
timestamp 1676037725
transform 1 0 135516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1473
timestamp 1676037725
transform 1 0 136620 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1479
timestamp 1676037725
transform 1 0 137172 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1489
timestamp 1676037725
transform 1 0 138092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1501
timestamp 1676037725
transform 1 0 139196 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1509
timestamp 1676037725
transform 1 0 139932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1513
timestamp 1676037725
transform 1 0 140300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1517
timestamp 1676037725
transform 1 0 140668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1527
timestamp 1676037725
transform 1 0 141588 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1539
timestamp 1676037725
transform 1 0 142692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1551
timestamp 1676037725
transform 1 0 143796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1555
timestamp 1676037725
transform 1 0 144164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1565
timestamp 1676037725
transform 1 0 145084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1569
timestamp 1676037725
transform 1 0 145452 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1577
timestamp 1676037725
transform 1 0 146188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1589
timestamp 1676037725
transform 1 0 147292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1593
timestamp 1676037725
transform 1 0 147660 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1603
timestamp 1676037725
transform 1 0 148580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1615
timestamp 1676037725
transform 1 0 149684 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1623
timestamp 1676037725
transform 1 0 150420 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1625
timestamp 1676037725
transform 1 0 150604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1637
timestamp 1676037725
transform 1 0 151708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1649
timestamp 1676037725
transform 1 0 152812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1661
timestamp 1676037725
transform 1 0 153916 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1673
timestamp 1676037725
transform 1 0 155020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1679
timestamp 1676037725
transform 1 0 155572 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1681
timestamp 1676037725
transform 1 0 155756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1693
timestamp 1676037725
transform 1 0 156860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1705
timestamp 1676037725
transform 1 0 157964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1717
timestamp 1676037725
transform 1 0 159068 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1729
timestamp 1676037725
transform 1 0 160172 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1735
timestamp 1676037725
transform 1 0 160724 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1737
timestamp 1676037725
transform 1 0 160908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1749
timestamp 1676037725
transform 1 0 162012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1761
timestamp 1676037725
transform 1 0 163116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1773
timestamp 1676037725
transform 1 0 164220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1785
timestamp 1676037725
transform 1 0 165324 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1791
timestamp 1676037725
transform 1 0 165876 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1793
timestamp 1676037725
transform 1 0 166060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1805
timestamp 1676037725
transform 1 0 167164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1817
timestamp 1676037725
transform 1 0 168268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1829
timestamp 1676037725
transform 1 0 169372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1841
timestamp 1676037725
transform 1 0 170476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1847
timestamp 1676037725
transform 1 0 171028 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1849
timestamp 1676037725
transform 1 0 171212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1861
timestamp 1676037725
transform 1 0 172316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1873
timestamp 1676037725
transform 1 0 173420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1885
timestamp 1676037725
transform 1 0 174524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1897
timestamp 1676037725
transform 1 0 175628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1903
timestamp 1676037725
transform 1 0 176180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1905
timestamp 1676037725
transform 1 0 176364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1917
timestamp 1676037725
transform 1 0 177468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1929
timestamp 1676037725
transform 1 0 178572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1941
timestamp 1676037725
transform 1 0 179676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1953
timestamp 1676037725
transform 1 0 180780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1959
timestamp 1676037725
transform 1 0 181332 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1961
timestamp 1676037725
transform 1 0 181516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1973
timestamp 1676037725
transform 1 0 182620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1985
timestamp 1676037725
transform 1 0 183724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1997
timestamp 1676037725
transform 1 0 184828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2009
timestamp 1676037725
transform 1 0 185932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2015
timestamp 1676037725
transform 1 0 186484 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2017
timestamp 1676037725
transform 1 0 186668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2029
timestamp 1676037725
transform 1 0 187772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2041
timestamp 1676037725
transform 1 0 188876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2053
timestamp 1676037725
transform 1 0 189980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2065
timestamp 1676037725
transform 1 0 191084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2071
timestamp 1676037725
transform 1 0 191636 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2073
timestamp 1676037725
transform 1 0 191820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2085
timestamp 1676037725
transform 1 0 192924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2097
timestamp 1676037725
transform 1 0 194028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2109
timestamp 1676037725
transform 1 0 195132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2121
timestamp 1676037725
transform 1 0 196236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2127
timestamp 1676037725
transform 1 0 196788 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2129
timestamp 1676037725
transform 1 0 196972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2141
timestamp 1676037725
transform 1 0 198076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2153
timestamp 1676037725
transform 1 0 199180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2165
timestamp 1676037725
transform 1 0 200284 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2177
timestamp 1676037725
transform 1 0 201388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2183
timestamp 1676037725
transform 1 0 201940 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2185
timestamp 1676037725
transform 1 0 202124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2197
timestamp 1676037725
transform 1 0 203228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2209
timestamp 1676037725
transform 1 0 204332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2221
timestamp 1676037725
transform 1 0 205436 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2233
timestamp 1676037725
transform 1 0 206540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2239
timestamp 1676037725
transform 1 0 207092 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2241
timestamp 1676037725
transform 1 0 207276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2253
timestamp 1676037725
transform 1 0 208380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2265
timestamp 1676037725
transform 1 0 209484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2277
timestamp 1676037725
transform 1 0 210588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2289
timestamp 1676037725
transform 1 0 211692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2295
timestamp 1676037725
transform 1 0 212244 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2297
timestamp 1676037725
transform 1 0 212428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2309
timestamp 1676037725
transform 1 0 213532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2321
timestamp 1676037725
transform 1 0 214636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2333
timestamp 1676037725
transform 1 0 215740 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2345
timestamp 1676037725
transform 1 0 216844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2351
timestamp 1676037725
transform 1 0 217396 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2353
timestamp 1676037725
transform 1 0 217580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2365
timestamp 1676037725
transform 1 0 218684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2377
timestamp 1676037725
transform 1 0 219788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2389
timestamp 1676037725
transform 1 0 220892 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2401
timestamp 1676037725
transform 1 0 221996 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2407
timestamp 1676037725
transform 1 0 222548 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2409
timestamp 1676037725
transform 1 0 222732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2421
timestamp 1676037725
transform 1 0 223836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2433
timestamp 1676037725
transform 1 0 224940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2445
timestamp 1676037725
transform 1 0 226044 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2457
timestamp 1676037725
transform 1 0 227148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2463
timestamp 1676037725
transform 1 0 227700 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2465
timestamp 1676037725
transform 1 0 227884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2477
timestamp 1676037725
transform 1 0 228988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2489
timestamp 1676037725
transform 1 0 230092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2501
timestamp 1676037725
transform 1 0 231196 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2513
timestamp 1676037725
transform 1 0 232300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2519
timestamp 1676037725
transform 1 0 232852 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2521
timestamp 1676037725
transform 1 0 233036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2533
timestamp 1676037725
transform 1 0 234140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2545
timestamp 1676037725
transform 1 0 235244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2557
timestamp 1676037725
transform 1 0 236348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2569
timestamp 1676037725
transform 1 0 237452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2575
timestamp 1676037725
transform 1 0 238004 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2577
timestamp 1676037725
transform 1 0 238188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2589
timestamp 1676037725
transform 1 0 239292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2601
timestamp 1676037725
transform 1 0 240396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2613
timestamp 1676037725
transform 1 0 241500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2625
timestamp 1676037725
transform 1 0 242604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2631
timestamp 1676037725
transform 1 0 243156 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2633
timestamp 1676037725
transform 1 0 243340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2645
timestamp 1676037725
transform 1 0 244444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2657
timestamp 1676037725
transform 1 0 245548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2669
timestamp 1676037725
transform 1 0 246652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2681
timestamp 1676037725
transform 1 0 247756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2687
timestamp 1676037725
transform 1 0 248308 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2689
timestamp 1676037725
transform 1 0 248492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2701
timestamp 1676037725
transform 1 0 249596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2713
timestamp 1676037725
transform 1 0 250700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2725
timestamp 1676037725
transform 1 0 251804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2737
timestamp 1676037725
transform 1 0 252908 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2743
timestamp 1676037725
transform 1 0 253460 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2745
timestamp 1676037725
transform 1 0 253644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2757
timestamp 1676037725
transform 1 0 254748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2769
timestamp 1676037725
transform 1 0 255852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2781
timestamp 1676037725
transform 1 0 256956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2793
timestamp 1676037725
transform 1 0 258060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2799
timestamp 1676037725
transform 1 0 258612 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2801
timestamp 1676037725
transform 1 0 258796 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2813
timestamp 1676037725
transform 1 0 259900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2825
timestamp 1676037725
transform 1 0 261004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2837
timestamp 1676037725
transform 1 0 262108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2849
timestamp 1676037725
transform 1 0 263212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2855
timestamp 1676037725
transform 1 0 263764 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2857
timestamp 1676037725
transform 1 0 263948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2869
timestamp 1676037725
transform 1 0 265052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2881
timestamp 1676037725
transform 1 0 266156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2893
timestamp 1676037725
transform 1 0 267260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2907
timestamp 1676037725
transform 1 0 268548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2911
timestamp 1676037725
transform 1 0 268916 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2913
timestamp 1676037725
transform 1 0 269100 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_2921
timestamp 1676037725
transform 1 0 269836 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2927
timestamp 1676037725
transform 1 0 270388 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_2930
timestamp 1676037725
transform 1 0 270664 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2943
timestamp 1676037725
transform 1 0 271860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2955
timestamp 1676037725
transform 1 0 272964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_2967
timestamp 1676037725
transform 1 0 274068 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2969
timestamp 1676037725
transform 1 0 274252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2981
timestamp 1676037725
transform 1 0 275356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_2993
timestamp 1676037725
transform 1 0 276460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3005
timestamp 1676037725
transform 1 0 277564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3017
timestamp 1676037725
transform 1 0 278668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3023
timestamp 1676037725
transform 1 0 279220 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3025
timestamp 1676037725
transform 1 0 279404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3037
timestamp 1676037725
transform 1 0 280508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3049
timestamp 1676037725
transform 1 0 281612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3061
timestamp 1676037725
transform 1 0 282716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3073
timestamp 1676037725
transform 1 0 283820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3079
timestamp 1676037725
transform 1 0 284372 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3081
timestamp 1676037725
transform 1 0 284556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3093
timestamp 1676037725
transform 1 0 285660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3105
timestamp 1676037725
transform 1 0 286764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3117
timestamp 1676037725
transform 1 0 287868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3129
timestamp 1676037725
transform 1 0 288972 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3135
timestamp 1676037725
transform 1 0 289524 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3137
timestamp 1676037725
transform 1 0 289708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3149
timestamp 1676037725
transform 1 0 290812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3161
timestamp 1676037725
transform 1 0 291916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3173
timestamp 1676037725
transform 1 0 293020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3185
timestamp 1676037725
transform 1 0 294124 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3191
timestamp 1676037725
transform 1 0 294676 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3193
timestamp 1676037725
transform 1 0 294860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3205
timestamp 1676037725
transform 1 0 295964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3217
timestamp 1676037725
transform 1 0 297068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3229
timestamp 1676037725
transform 1 0 298172 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3241
timestamp 1676037725
transform 1 0 299276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3247
timestamp 1676037725
transform 1 0 299828 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3249
timestamp 1676037725
transform 1 0 300012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3261
timestamp 1676037725
transform 1 0 301116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3273
timestamp 1676037725
transform 1 0 302220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3285
timestamp 1676037725
transform 1 0 303324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3297
timestamp 1676037725
transform 1 0 304428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3303
timestamp 1676037725
transform 1 0 304980 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3305
timestamp 1676037725
transform 1 0 305164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3317
timestamp 1676037725
transform 1 0 306268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3329
timestamp 1676037725
transform 1 0 307372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3341
timestamp 1676037725
transform 1 0 308476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3353
timestamp 1676037725
transform 1 0 309580 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3359
timestamp 1676037725
transform 1 0 310132 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3361
timestamp 1676037725
transform 1 0 310316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3373
timestamp 1676037725
transform 1 0 311420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3385
timestamp 1676037725
transform 1 0 312524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3397
timestamp 1676037725
transform 1 0 313628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3409
timestamp 1676037725
transform 1 0 314732 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3415
timestamp 1676037725
transform 1 0 315284 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3417
timestamp 1676037725
transform 1 0 315468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3429
timestamp 1676037725
transform 1 0 316572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3441
timestamp 1676037725
transform 1 0 317676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3453
timestamp 1676037725
transform 1 0 318780 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3465
timestamp 1676037725
transform 1 0 319884 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3471
timestamp 1676037725
transform 1 0 320436 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3473
timestamp 1676037725
transform 1 0 320620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3485
timestamp 1676037725
transform 1 0 321724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3497
timestamp 1676037725
transform 1 0 322828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3509
timestamp 1676037725
transform 1 0 323932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3521
timestamp 1676037725
transform 1 0 325036 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3527
timestamp 1676037725
transform 1 0 325588 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3529
timestamp 1676037725
transform 1 0 325772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3541
timestamp 1676037725
transform 1 0 326876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3553
timestamp 1676037725
transform 1 0 327980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3565
timestamp 1676037725
transform 1 0 329084 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3577
timestamp 1676037725
transform 1 0 330188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3583
timestamp 1676037725
transform 1 0 330740 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3585
timestamp 1676037725
transform 1 0 330924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3597
timestamp 1676037725
transform 1 0 332028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3609
timestamp 1676037725
transform 1 0 333132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3621
timestamp 1676037725
transform 1 0 334236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3633
timestamp 1676037725
transform 1 0 335340 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3639
timestamp 1676037725
transform 1 0 335892 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3641
timestamp 1676037725
transform 1 0 336076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3653
timestamp 1676037725
transform 1 0 337180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3665
timestamp 1676037725
transform 1 0 338284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3677
timestamp 1676037725
transform 1 0 339388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3689
timestamp 1676037725
transform 1 0 340492 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3695
timestamp 1676037725
transform 1 0 341044 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3697
timestamp 1676037725
transform 1 0 341228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3709
timestamp 1676037725
transform 1 0 342332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3721
timestamp 1676037725
transform 1 0 343436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3733
timestamp 1676037725
transform 1 0 344540 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3745
timestamp 1676037725
transform 1 0 345644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3751
timestamp 1676037725
transform 1 0 346196 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3753
timestamp 1676037725
transform 1 0 346380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3765
timestamp 1676037725
transform 1 0 347484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3777
timestamp 1676037725
transform 1 0 348588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3789
timestamp 1676037725
transform 1 0 349692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3801
timestamp 1676037725
transform 1 0 350796 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3807
timestamp 1676037725
transform 1 0 351348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3809
timestamp 1676037725
transform 1 0 351532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3821
timestamp 1676037725
transform 1 0 352636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3833
timestamp 1676037725
transform 1 0 353740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3845
timestamp 1676037725
transform 1 0 354844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3857
timestamp 1676037725
transform 1 0 355948 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3863
timestamp 1676037725
transform 1 0 356500 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3865
timestamp 1676037725
transform 1 0 356684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3877
timestamp 1676037725
transform 1 0 357788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3889
timestamp 1676037725
transform 1 0 358892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3901
timestamp 1676037725
transform 1 0 359996 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3913
timestamp 1676037725
transform 1 0 361100 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3919
timestamp 1676037725
transform 1 0 361652 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3921
timestamp 1676037725
transform 1 0 361836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3933
timestamp 1676037725
transform 1 0 362940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3945
timestamp 1676037725
transform 1 0 364044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3957
timestamp 1676037725
transform 1 0 365148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3969
timestamp 1676037725
transform 1 0 366252 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3975
timestamp 1676037725
transform 1 0 366804 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3977
timestamp 1676037725
transform 1 0 366988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3989
timestamp 1676037725
transform 1 0 368092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4001
timestamp 1676037725
transform 1 0 369196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4013
timestamp 1676037725
transform 1 0 370300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4025
timestamp 1676037725
transform 1 0 371404 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4031
timestamp 1676037725
transform 1 0 371956 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4033
timestamp 1676037725
transform 1 0 372140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4045
timestamp 1676037725
transform 1 0 373244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4057
timestamp 1676037725
transform 1 0 374348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4069
timestamp 1676037725
transform 1 0 375452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4081
timestamp 1676037725
transform 1 0 376556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4087
timestamp 1676037725
transform 1 0 377108 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4089
timestamp 1676037725
transform 1 0 377292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4101
timestamp 1676037725
transform 1 0 378396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4113
timestamp 1676037725
transform 1 0 379500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4125
timestamp 1676037725
transform 1 0 380604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4137
timestamp 1676037725
transform 1 0 381708 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4143
timestamp 1676037725
transform 1 0 382260 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4145
timestamp 1676037725
transform 1 0 382444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4157
timestamp 1676037725
transform 1 0 383548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4169
timestamp 1676037725
transform 1 0 384652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4181
timestamp 1676037725
transform 1 0 385756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4193
timestamp 1676037725
transform 1 0 386860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4199
timestamp 1676037725
transform 1 0 387412 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4201
timestamp 1676037725
transform 1 0 387596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4213
timestamp 1676037725
transform 1 0 388700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4225
timestamp 1676037725
transform 1 0 389804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4237
timestamp 1676037725
transform 1 0 390908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4249
timestamp 1676037725
transform 1 0 392012 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4255
timestamp 1676037725
transform 1 0 392564 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4257
timestamp 1676037725
transform 1 0 392748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4269
timestamp 1676037725
transform 1 0 393852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4281
timestamp 1676037725
transform 1 0 394956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4293
timestamp 1676037725
transform 1 0 396060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4305
timestamp 1676037725
transform 1 0 397164 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4311
timestamp 1676037725
transform 1 0 397716 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4313
timestamp 1676037725
transform 1 0 397900 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4325
timestamp 1676037725
transform 1 0 399004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4337
timestamp 1676037725
transform 1 0 400108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4349
timestamp 1676037725
transform 1 0 401212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4361
timestamp 1676037725
transform 1 0 402316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4367
timestamp 1676037725
transform 1 0 402868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4369
timestamp 1676037725
transform 1 0 403052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4381
timestamp 1676037725
transform 1 0 404156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4393
timestamp 1676037725
transform 1 0 405260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4405
timestamp 1676037725
transform 1 0 406364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4417
timestamp 1676037725
transform 1 0 407468 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4423
timestamp 1676037725
transform 1 0 408020 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4425
timestamp 1676037725
transform 1 0 408204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4437
timestamp 1676037725
transform 1 0 409308 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4449
timestamp 1676037725
transform 1 0 410412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4461
timestamp 1676037725
transform 1 0 411516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4473
timestamp 1676037725
transform 1 0 412620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4479
timestamp 1676037725
transform 1 0 413172 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4481
timestamp 1676037725
transform 1 0 413356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4493
timestamp 1676037725
transform 1 0 414460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4505
timestamp 1676037725
transform 1 0 415564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4517
timestamp 1676037725
transform 1 0 416668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4529
timestamp 1676037725
transform 1 0 417772 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4535
timestamp 1676037725
transform 1 0 418324 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4537
timestamp 1676037725
transform 1 0 418508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4549
timestamp 1676037725
transform 1 0 419612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4561
timestamp 1676037725
transform 1 0 420716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4573
timestamp 1676037725
transform 1 0 421820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4585
timestamp 1676037725
transform 1 0 422924 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4591
timestamp 1676037725
transform 1 0 423476 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4593
timestamp 1676037725
transform 1 0 423660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4605
timestamp 1676037725
transform 1 0 424764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4617
timestamp 1676037725
transform 1 0 425868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4629
timestamp 1676037725
transform 1 0 426972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4641
timestamp 1676037725
transform 1 0 428076 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4647
timestamp 1676037725
transform 1 0 428628 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4649
timestamp 1676037725
transform 1 0 428812 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4661
timestamp 1676037725
transform 1 0 429916 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4673
timestamp 1676037725
transform 1 0 431020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4685
timestamp 1676037725
transform 1 0 432124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4697
timestamp 1676037725
transform 1 0 433228 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4703
timestamp 1676037725
transform 1 0 433780 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4705
timestamp 1676037725
transform 1 0 433964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4717
timestamp 1676037725
transform 1 0 435068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4729
timestamp 1676037725
transform 1 0 436172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4741
timestamp 1676037725
transform 1 0 437276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4753
timestamp 1676037725
transform 1 0 438380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4759
timestamp 1676037725
transform 1 0 438932 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4761
timestamp 1676037725
transform 1 0 439116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4773
timestamp 1676037725
transform 1 0 440220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4785
timestamp 1676037725
transform 1 0 441324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4797
timestamp 1676037725
transform 1 0 442428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4809
timestamp 1676037725
transform 1 0 443532 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4815
timestamp 1676037725
transform 1 0 444084 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4817
timestamp 1676037725
transform 1 0 444268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4829
timestamp 1676037725
transform 1 0 445372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4841
timestamp 1676037725
transform 1 0 446476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4853
timestamp 1676037725
transform 1 0 447580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4865
timestamp 1676037725
transform 1 0 448684 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4871
timestamp 1676037725
transform 1 0 449236 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4873
timestamp 1676037725
transform 1 0 449420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4885
timestamp 1676037725
transform 1 0 450524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4897
timestamp 1676037725
transform 1 0 451628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4909
timestamp 1676037725
transform 1 0 452732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4921
timestamp 1676037725
transform 1 0 453836 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4927
timestamp 1676037725
transform 1 0 454388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4929
timestamp 1676037725
transform 1 0 454572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4941
timestamp 1676037725
transform 1 0 455676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4953
timestamp 1676037725
transform 1 0 456780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4965
timestamp 1676037725
transform 1 0 457884 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_4977
timestamp 1676037725
transform 1 0 458988 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_4983
timestamp 1676037725
transform 1 0 459540 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4985
timestamp 1676037725
transform 1 0 459724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_4997
timestamp 1676037725
transform 1 0 460828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5009
timestamp 1676037725
transform 1 0 461932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5021
timestamp 1676037725
transform 1 0 463036 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5033
timestamp 1676037725
transform 1 0 464140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5039
timestamp 1676037725
transform 1 0 464692 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5041
timestamp 1676037725
transform 1 0 464876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5053
timestamp 1676037725
transform 1 0 465980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5065
timestamp 1676037725
transform 1 0 467084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5077
timestamp 1676037725
transform 1 0 468188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5089
timestamp 1676037725
transform 1 0 469292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5095
timestamp 1676037725
transform 1 0 469844 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5097
timestamp 1676037725
transform 1 0 470028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5109
timestamp 1676037725
transform 1 0 471132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5121
timestamp 1676037725
transform 1 0 472236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5133
timestamp 1676037725
transform 1 0 473340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5145
timestamp 1676037725
transform 1 0 474444 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5151
timestamp 1676037725
transform 1 0 474996 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5153
timestamp 1676037725
transform 1 0 475180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5165
timestamp 1676037725
transform 1 0 476284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5177
timestamp 1676037725
transform 1 0 477388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5189
timestamp 1676037725
transform 1 0 478492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5201
timestamp 1676037725
transform 1 0 479596 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5207
timestamp 1676037725
transform 1 0 480148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5209
timestamp 1676037725
transform 1 0 480332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5221
timestamp 1676037725
transform 1 0 481436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5233
timestamp 1676037725
transform 1 0 482540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5245
timestamp 1676037725
transform 1 0 483644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5257
timestamp 1676037725
transform 1 0 484748 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5263
timestamp 1676037725
transform 1 0 485300 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5265
timestamp 1676037725
transform 1 0 485484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5277
timestamp 1676037725
transform 1 0 486588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5289
timestamp 1676037725
transform 1 0 487692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5301
timestamp 1676037725
transform 1 0 488796 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5313
timestamp 1676037725
transform 1 0 489900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5319
timestamp 1676037725
transform 1 0 490452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5321
timestamp 1676037725
transform 1 0 490636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5333
timestamp 1676037725
transform 1 0 491740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5345
timestamp 1676037725
transform 1 0 492844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5357
timestamp 1676037725
transform 1 0 493948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5369
timestamp 1676037725
transform 1 0 495052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5375
timestamp 1676037725
transform 1 0 495604 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5377
timestamp 1676037725
transform 1 0 495788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5389
timestamp 1676037725
transform 1 0 496892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5401
timestamp 1676037725
transform 1 0 497996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5413
timestamp 1676037725
transform 1 0 499100 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5425
timestamp 1676037725
transform 1 0 500204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5431
timestamp 1676037725
transform 1 0 500756 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5433
timestamp 1676037725
transform 1 0 500940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5445
timestamp 1676037725
transform 1 0 502044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5457
timestamp 1676037725
transform 1 0 503148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5469
timestamp 1676037725
transform 1 0 504252 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5481
timestamp 1676037725
transform 1 0 505356 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5487
timestamp 1676037725
transform 1 0 505908 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5489
timestamp 1676037725
transform 1 0 506092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5501
timestamp 1676037725
transform 1 0 507196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5513
timestamp 1676037725
transform 1 0 508300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5525
timestamp 1676037725
transform 1 0 509404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5537
timestamp 1676037725
transform 1 0 510508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5543
timestamp 1676037725
transform 1 0 511060 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5545
timestamp 1676037725
transform 1 0 511244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5557
timestamp 1676037725
transform 1 0 512348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5569
timestamp 1676037725
transform 1 0 513452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5581
timestamp 1676037725
transform 1 0 514556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5593
timestamp 1676037725
transform 1 0 515660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5599
timestamp 1676037725
transform 1 0 516212 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5601
timestamp 1676037725
transform 1 0 516396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5613
timestamp 1676037725
transform 1 0 517500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5625
timestamp 1676037725
transform 1 0 518604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5637
timestamp 1676037725
transform 1 0 519708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5649
timestamp 1676037725
transform 1 0 520812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5655
timestamp 1676037725
transform 1 0 521364 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5657
timestamp 1676037725
transform 1 0 521548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5669
timestamp 1676037725
transform 1 0 522652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5681
timestamp 1676037725
transform 1 0 523756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5693
timestamp 1676037725
transform 1 0 524860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_5705
timestamp 1676037725
transform 1 0 525964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_5711
timestamp 1676037725
transform 1 0 526516 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5713
timestamp 1676037725
transform 1 0 526700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_5725
timestamp 1676037725
transform 1 0 527804 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1676037725
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1676037725
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1676037725
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1676037725
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1676037725
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1676037725
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1676037725
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1676037725
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1676037725
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1676037725
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1676037725
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1676037725
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1676037725
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1676037725
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1676037725
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1676037725
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1676037725
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1676037725
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1676037725
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1676037725
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1676037725
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1676037725
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1676037725
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1676037725
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1676037725
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1676037725
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1676037725
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1676037725
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1676037725
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1676037725
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1676037725
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1676037725
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1676037725
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1676037725
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1676037725
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1676037725
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1676037725
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1676037725
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1676037725
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1676037725
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1676037725
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1676037725
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1676037725
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1676037725
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1676037725
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1676037725
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1676037725
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1676037725
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1676037725
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1676037725
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1676037725
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1676037725
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1676037725
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1676037725
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1676037725
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1676037725
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1676037725
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1676037725
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1141
timestamp 1676037725
transform 1 0 106076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1146
timestamp 1676037725
transform 1 0 106536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1149
timestamp 1676037725
transform 1 0 106812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1160
timestamp 1676037725
transform 1 0 107824 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1168
timestamp 1676037725
transform 1 0 108560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1171
timestamp 1676037725
transform 1 0 108836 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1184
timestamp 1676037725
transform 1 0 110032 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1196
timestamp 1676037725
transform 1 0 111136 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1676037725
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1217
timestamp 1676037725
transform 1 0 113068 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1221
timestamp 1676037725
transform 1 0 113436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1233
timestamp 1676037725
transform 1 0 114540 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1241
timestamp 1676037725
transform 1 0 115276 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1245
timestamp 1676037725
transform 1 0 115644 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1258
timestamp 1676037725
transform 1 0 116840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1261
timestamp 1676037725
transform 1 0 117116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1272
timestamp 1676037725
transform 1 0 118128 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1282
timestamp 1676037725
transform 1 0 119048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1295
timestamp 1676037725
transform 1 0 120244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1308
timestamp 1676037725
transform 1 0 121440 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1317
timestamp 1676037725
transform 1 0 122268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1332
timestamp 1676037725
transform 1 0 123648 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1345
timestamp 1676037725
transform 1 0 124844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1357
timestamp 1676037725
transform 1 0 125948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1369
timestamp 1676037725
transform 1 0 127052 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1373
timestamp 1676037725
transform 1 0 127420 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1383
timestamp 1676037725
transform 1 0 128340 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1395
timestamp 1676037725
transform 1 0 129444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1401
timestamp 1676037725
transform 1 0 129996 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1404
timestamp 1676037725
transform 1 0 130272 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1414
timestamp 1676037725
transform 1 0 131192 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1426
timestamp 1676037725
transform 1 0 132296 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1429
timestamp 1676037725
transform 1 0 132572 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1437
timestamp 1676037725
transform 1 0 133308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1442
timestamp 1676037725
transform 1 0 133768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1452
timestamp 1676037725
transform 1 0 134688 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1464
timestamp 1676037725
transform 1 0 135792 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1476
timestamp 1676037725
transform 1 0 136896 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1485
timestamp 1676037725
transform 1 0 137724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1489
timestamp 1676037725
transform 1 0 138092 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1492
timestamp 1676037725
transform 1 0 138368 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1502
timestamp 1676037725
transform 1 0 139288 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1514
timestamp 1676037725
transform 1 0 140392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1526
timestamp 1676037725
transform 1 0 141496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1530
timestamp 1676037725
transform 1 0 141864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1533
timestamp 1676037725
transform 1 0 142140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1539
timestamp 1676037725
transform 1 0 142692 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1541
timestamp 1676037725
transform 1 0 142876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1553
timestamp 1676037725
transform 1 0 143980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1565
timestamp 1676037725
transform 1 0 145084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1577
timestamp 1676037725
transform 1 0 146188 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1589
timestamp 1676037725
transform 1 0 147292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1595
timestamp 1676037725
transform 1 0 147844 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1597
timestamp 1676037725
transform 1 0 148028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1609
timestamp 1676037725
transform 1 0 149132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1621
timestamp 1676037725
transform 1 0 150236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1633
timestamp 1676037725
transform 1 0 151340 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1645
timestamp 1676037725
transform 1 0 152444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1651
timestamp 1676037725
transform 1 0 152996 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1653
timestamp 1676037725
transform 1 0 153180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1665
timestamp 1676037725
transform 1 0 154284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1677
timestamp 1676037725
transform 1 0 155388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1689
timestamp 1676037725
transform 1 0 156492 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1701
timestamp 1676037725
transform 1 0 157596 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1707
timestamp 1676037725
transform 1 0 158148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1709
timestamp 1676037725
transform 1 0 158332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1721
timestamp 1676037725
transform 1 0 159436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1733
timestamp 1676037725
transform 1 0 160540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1745
timestamp 1676037725
transform 1 0 161644 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1757
timestamp 1676037725
transform 1 0 162748 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1763
timestamp 1676037725
transform 1 0 163300 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1765
timestamp 1676037725
transform 1 0 163484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1777
timestamp 1676037725
transform 1 0 164588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1789
timestamp 1676037725
transform 1 0 165692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1801
timestamp 1676037725
transform 1 0 166796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1813
timestamp 1676037725
transform 1 0 167900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1819
timestamp 1676037725
transform 1 0 168452 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1821
timestamp 1676037725
transform 1 0 168636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1833
timestamp 1676037725
transform 1 0 169740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1845
timestamp 1676037725
transform 1 0 170844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1857
timestamp 1676037725
transform 1 0 171948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1869
timestamp 1676037725
transform 1 0 173052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1875
timestamp 1676037725
transform 1 0 173604 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1877
timestamp 1676037725
transform 1 0 173788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1889
timestamp 1676037725
transform 1 0 174892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1901
timestamp 1676037725
transform 1 0 175996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1913
timestamp 1676037725
transform 1 0 177100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1925
timestamp 1676037725
transform 1 0 178204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1931
timestamp 1676037725
transform 1 0 178756 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1933
timestamp 1676037725
transform 1 0 178940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1945
timestamp 1676037725
transform 1 0 180044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1957
timestamp 1676037725
transform 1 0 181148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1969
timestamp 1676037725
transform 1 0 182252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1981
timestamp 1676037725
transform 1 0 183356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1987
timestamp 1676037725
transform 1 0 183908 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1989
timestamp 1676037725
transform 1 0 184092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2001
timestamp 1676037725
transform 1 0 185196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2013
timestamp 1676037725
transform 1 0 186300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2025
timestamp 1676037725
transform 1 0 187404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2037
timestamp 1676037725
transform 1 0 188508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2043
timestamp 1676037725
transform 1 0 189060 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2045
timestamp 1676037725
transform 1 0 189244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2057
timestamp 1676037725
transform 1 0 190348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2069
timestamp 1676037725
transform 1 0 191452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2081
timestamp 1676037725
transform 1 0 192556 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2093
timestamp 1676037725
transform 1 0 193660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2099
timestamp 1676037725
transform 1 0 194212 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2101
timestamp 1676037725
transform 1 0 194396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2113
timestamp 1676037725
transform 1 0 195500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2125
timestamp 1676037725
transform 1 0 196604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2137
timestamp 1676037725
transform 1 0 197708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2149
timestamp 1676037725
transform 1 0 198812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2155
timestamp 1676037725
transform 1 0 199364 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2157
timestamp 1676037725
transform 1 0 199548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2169
timestamp 1676037725
transform 1 0 200652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2181
timestamp 1676037725
transform 1 0 201756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2193
timestamp 1676037725
transform 1 0 202860 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2205
timestamp 1676037725
transform 1 0 203964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2211
timestamp 1676037725
transform 1 0 204516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2213
timestamp 1676037725
transform 1 0 204700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2225
timestamp 1676037725
transform 1 0 205804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2237
timestamp 1676037725
transform 1 0 206908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2249
timestamp 1676037725
transform 1 0 208012 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2261
timestamp 1676037725
transform 1 0 209116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2267
timestamp 1676037725
transform 1 0 209668 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2269
timestamp 1676037725
transform 1 0 209852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2281
timestamp 1676037725
transform 1 0 210956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2293
timestamp 1676037725
transform 1 0 212060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2305
timestamp 1676037725
transform 1 0 213164 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2317
timestamp 1676037725
transform 1 0 214268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2323
timestamp 1676037725
transform 1 0 214820 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2325
timestamp 1676037725
transform 1 0 215004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2337
timestamp 1676037725
transform 1 0 216108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2349
timestamp 1676037725
transform 1 0 217212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2361
timestamp 1676037725
transform 1 0 218316 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2373
timestamp 1676037725
transform 1 0 219420 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2379
timestamp 1676037725
transform 1 0 219972 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2381
timestamp 1676037725
transform 1 0 220156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2393
timestamp 1676037725
transform 1 0 221260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2405
timestamp 1676037725
transform 1 0 222364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2417
timestamp 1676037725
transform 1 0 223468 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2429
timestamp 1676037725
transform 1 0 224572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2435
timestamp 1676037725
transform 1 0 225124 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2437
timestamp 1676037725
transform 1 0 225308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2449
timestamp 1676037725
transform 1 0 226412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2461
timestamp 1676037725
transform 1 0 227516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2473
timestamp 1676037725
transform 1 0 228620 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2485
timestamp 1676037725
transform 1 0 229724 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2491
timestamp 1676037725
transform 1 0 230276 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2493
timestamp 1676037725
transform 1 0 230460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2505
timestamp 1676037725
transform 1 0 231564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2517
timestamp 1676037725
transform 1 0 232668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2529
timestamp 1676037725
transform 1 0 233772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2541
timestamp 1676037725
transform 1 0 234876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2547
timestamp 1676037725
transform 1 0 235428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2549
timestamp 1676037725
transform 1 0 235612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2561
timestamp 1676037725
transform 1 0 236716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2573
timestamp 1676037725
transform 1 0 237820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2585
timestamp 1676037725
transform 1 0 238924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2597
timestamp 1676037725
transform 1 0 240028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2603
timestamp 1676037725
transform 1 0 240580 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2605
timestamp 1676037725
transform 1 0 240764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2617
timestamp 1676037725
transform 1 0 241868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2629
timestamp 1676037725
transform 1 0 242972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2641
timestamp 1676037725
transform 1 0 244076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2653
timestamp 1676037725
transform 1 0 245180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2659
timestamp 1676037725
transform 1 0 245732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2661
timestamp 1676037725
transform 1 0 245916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2673
timestamp 1676037725
transform 1 0 247020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2685
timestamp 1676037725
transform 1 0 248124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2697
timestamp 1676037725
transform 1 0 249228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2709
timestamp 1676037725
transform 1 0 250332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2715
timestamp 1676037725
transform 1 0 250884 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2717
timestamp 1676037725
transform 1 0 251068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2729
timestamp 1676037725
transform 1 0 252172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2741
timestamp 1676037725
transform 1 0 253276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2753
timestamp 1676037725
transform 1 0 254380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2765
timestamp 1676037725
transform 1 0 255484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2771
timestamp 1676037725
transform 1 0 256036 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2773
timestamp 1676037725
transform 1 0 256220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2785
timestamp 1676037725
transform 1 0 257324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2797
timestamp 1676037725
transform 1 0 258428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2809
timestamp 1676037725
transform 1 0 259532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2821
timestamp 1676037725
transform 1 0 260636 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2827
timestamp 1676037725
transform 1 0 261188 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_2829
timestamp 1676037725
transform 1 0 261372 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_2837
timestamp 1676037725
transform 1 0 262108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2841
timestamp 1676037725
transform 1 0 262476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2847
timestamp 1676037725
transform 1 0 263028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2850
timestamp 1676037725
transform 1 0 263304 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2863
timestamp 1676037725
transform 1 0 264500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2875
timestamp 1676037725
transform 1 0 265604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_2881
timestamp 1676037725
transform 1 0 266156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_2885
timestamp 1676037725
transform 1 0 266524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2890
timestamp 1676037725
transform 1 0 266984 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2903
timestamp 1676037725
transform 1 0 268180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_2916
timestamp 1676037725
transform 1 0 269376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2920
timestamp 1676037725
transform 1 0 269744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_2930
timestamp 1676037725
transform 1 0 270664 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_2938
timestamp 1676037725
transform 1 0 271400 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2941
timestamp 1676037725
transform 1 0 271676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2953
timestamp 1676037725
transform 1 0 272780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2965
timestamp 1676037725
transform 1 0 273884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2977
timestamp 1676037725
transform 1 0 274988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_2989
timestamp 1676037725
transform 1 0 276092 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_2995
timestamp 1676037725
transform 1 0 276644 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_2997
timestamp 1676037725
transform 1 0 276828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3009
timestamp 1676037725
transform 1 0 277932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3021
timestamp 1676037725
transform 1 0 279036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3033
timestamp 1676037725
transform 1 0 280140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3045
timestamp 1676037725
transform 1 0 281244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3051
timestamp 1676037725
transform 1 0 281796 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3053
timestamp 1676037725
transform 1 0 281980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3065
timestamp 1676037725
transform 1 0 283084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3077
timestamp 1676037725
transform 1 0 284188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3089
timestamp 1676037725
transform 1 0 285292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3101
timestamp 1676037725
transform 1 0 286396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3107
timestamp 1676037725
transform 1 0 286948 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3109
timestamp 1676037725
transform 1 0 287132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3121
timestamp 1676037725
transform 1 0 288236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3133
timestamp 1676037725
transform 1 0 289340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3145
timestamp 1676037725
transform 1 0 290444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3157
timestamp 1676037725
transform 1 0 291548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3163
timestamp 1676037725
transform 1 0 292100 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3165
timestamp 1676037725
transform 1 0 292284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3177
timestamp 1676037725
transform 1 0 293388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3189
timestamp 1676037725
transform 1 0 294492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3201
timestamp 1676037725
transform 1 0 295596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3213
timestamp 1676037725
transform 1 0 296700 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3219
timestamp 1676037725
transform 1 0 297252 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3221
timestamp 1676037725
transform 1 0 297436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3233
timestamp 1676037725
transform 1 0 298540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3245
timestamp 1676037725
transform 1 0 299644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3257
timestamp 1676037725
transform 1 0 300748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3269
timestamp 1676037725
transform 1 0 301852 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3275
timestamp 1676037725
transform 1 0 302404 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3277
timestamp 1676037725
transform 1 0 302588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3289
timestamp 1676037725
transform 1 0 303692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3301
timestamp 1676037725
transform 1 0 304796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3313
timestamp 1676037725
transform 1 0 305900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3325
timestamp 1676037725
transform 1 0 307004 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3331
timestamp 1676037725
transform 1 0 307556 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3333
timestamp 1676037725
transform 1 0 307740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3345
timestamp 1676037725
transform 1 0 308844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3357
timestamp 1676037725
transform 1 0 309948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3369
timestamp 1676037725
transform 1 0 311052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3381
timestamp 1676037725
transform 1 0 312156 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3387
timestamp 1676037725
transform 1 0 312708 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3389
timestamp 1676037725
transform 1 0 312892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3401
timestamp 1676037725
transform 1 0 313996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3413
timestamp 1676037725
transform 1 0 315100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3425
timestamp 1676037725
transform 1 0 316204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3437
timestamp 1676037725
transform 1 0 317308 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3443
timestamp 1676037725
transform 1 0 317860 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3445
timestamp 1676037725
transform 1 0 318044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3457
timestamp 1676037725
transform 1 0 319148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3469
timestamp 1676037725
transform 1 0 320252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3481
timestamp 1676037725
transform 1 0 321356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3493
timestamp 1676037725
transform 1 0 322460 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3499
timestamp 1676037725
transform 1 0 323012 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3501
timestamp 1676037725
transform 1 0 323196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3513
timestamp 1676037725
transform 1 0 324300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3525
timestamp 1676037725
transform 1 0 325404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3537
timestamp 1676037725
transform 1 0 326508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3549
timestamp 1676037725
transform 1 0 327612 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3555
timestamp 1676037725
transform 1 0 328164 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3557
timestamp 1676037725
transform 1 0 328348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3569
timestamp 1676037725
transform 1 0 329452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3581
timestamp 1676037725
transform 1 0 330556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3593
timestamp 1676037725
transform 1 0 331660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3605
timestamp 1676037725
transform 1 0 332764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3611
timestamp 1676037725
transform 1 0 333316 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3613
timestamp 1676037725
transform 1 0 333500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3625
timestamp 1676037725
transform 1 0 334604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3637
timestamp 1676037725
transform 1 0 335708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3649
timestamp 1676037725
transform 1 0 336812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3661
timestamp 1676037725
transform 1 0 337916 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3667
timestamp 1676037725
transform 1 0 338468 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3669
timestamp 1676037725
transform 1 0 338652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3681
timestamp 1676037725
transform 1 0 339756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3693
timestamp 1676037725
transform 1 0 340860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3705
timestamp 1676037725
transform 1 0 341964 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3717
timestamp 1676037725
transform 1 0 343068 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3723
timestamp 1676037725
transform 1 0 343620 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3725
timestamp 1676037725
transform 1 0 343804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3737
timestamp 1676037725
transform 1 0 344908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3749
timestamp 1676037725
transform 1 0 346012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3761
timestamp 1676037725
transform 1 0 347116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3773
timestamp 1676037725
transform 1 0 348220 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3779
timestamp 1676037725
transform 1 0 348772 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3781
timestamp 1676037725
transform 1 0 348956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3793
timestamp 1676037725
transform 1 0 350060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3805
timestamp 1676037725
transform 1 0 351164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3817
timestamp 1676037725
transform 1 0 352268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3829
timestamp 1676037725
transform 1 0 353372 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3835
timestamp 1676037725
transform 1 0 353924 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3837
timestamp 1676037725
transform 1 0 354108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3849
timestamp 1676037725
transform 1 0 355212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3861
timestamp 1676037725
transform 1 0 356316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3873
timestamp 1676037725
transform 1 0 357420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3885
timestamp 1676037725
transform 1 0 358524 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3891
timestamp 1676037725
transform 1 0 359076 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3893
timestamp 1676037725
transform 1 0 359260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3905
timestamp 1676037725
transform 1 0 360364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3917
timestamp 1676037725
transform 1 0 361468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3929
timestamp 1676037725
transform 1 0 362572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3941
timestamp 1676037725
transform 1 0 363676 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3947
timestamp 1676037725
transform 1 0 364228 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3949
timestamp 1676037725
transform 1 0 364412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3961
timestamp 1676037725
transform 1 0 365516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3973
timestamp 1676037725
transform 1 0 366620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3985
timestamp 1676037725
transform 1 0 367724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3997
timestamp 1676037725
transform 1 0 368828 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4003
timestamp 1676037725
transform 1 0 369380 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4005
timestamp 1676037725
transform 1 0 369564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4017
timestamp 1676037725
transform 1 0 370668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4029
timestamp 1676037725
transform 1 0 371772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4041
timestamp 1676037725
transform 1 0 372876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4053
timestamp 1676037725
transform 1 0 373980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4059
timestamp 1676037725
transform 1 0 374532 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4061
timestamp 1676037725
transform 1 0 374716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4073
timestamp 1676037725
transform 1 0 375820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4085
timestamp 1676037725
transform 1 0 376924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4097
timestamp 1676037725
transform 1 0 378028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4109
timestamp 1676037725
transform 1 0 379132 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4115
timestamp 1676037725
transform 1 0 379684 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4117
timestamp 1676037725
transform 1 0 379868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4129
timestamp 1676037725
transform 1 0 380972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4141
timestamp 1676037725
transform 1 0 382076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4153
timestamp 1676037725
transform 1 0 383180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4165
timestamp 1676037725
transform 1 0 384284 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4171
timestamp 1676037725
transform 1 0 384836 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4173
timestamp 1676037725
transform 1 0 385020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4185
timestamp 1676037725
transform 1 0 386124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4197
timestamp 1676037725
transform 1 0 387228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4209
timestamp 1676037725
transform 1 0 388332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4221
timestamp 1676037725
transform 1 0 389436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4227
timestamp 1676037725
transform 1 0 389988 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4229
timestamp 1676037725
transform 1 0 390172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4241
timestamp 1676037725
transform 1 0 391276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4253
timestamp 1676037725
transform 1 0 392380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4265
timestamp 1676037725
transform 1 0 393484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4277
timestamp 1676037725
transform 1 0 394588 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4283
timestamp 1676037725
transform 1 0 395140 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4285
timestamp 1676037725
transform 1 0 395324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4297
timestamp 1676037725
transform 1 0 396428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4309
timestamp 1676037725
transform 1 0 397532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4321
timestamp 1676037725
transform 1 0 398636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4333
timestamp 1676037725
transform 1 0 399740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4339
timestamp 1676037725
transform 1 0 400292 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4341
timestamp 1676037725
transform 1 0 400476 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4353
timestamp 1676037725
transform 1 0 401580 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4365
timestamp 1676037725
transform 1 0 402684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4377
timestamp 1676037725
transform 1 0 403788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4389
timestamp 1676037725
transform 1 0 404892 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4395
timestamp 1676037725
transform 1 0 405444 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4397
timestamp 1676037725
transform 1 0 405628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4409
timestamp 1676037725
transform 1 0 406732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4421
timestamp 1676037725
transform 1 0 407836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4433
timestamp 1676037725
transform 1 0 408940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4445
timestamp 1676037725
transform 1 0 410044 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4451
timestamp 1676037725
transform 1 0 410596 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4453
timestamp 1676037725
transform 1 0 410780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4465
timestamp 1676037725
transform 1 0 411884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4477
timestamp 1676037725
transform 1 0 412988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4489
timestamp 1676037725
transform 1 0 414092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4501
timestamp 1676037725
transform 1 0 415196 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4507
timestamp 1676037725
transform 1 0 415748 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4509
timestamp 1676037725
transform 1 0 415932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4521
timestamp 1676037725
transform 1 0 417036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4533
timestamp 1676037725
transform 1 0 418140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4545
timestamp 1676037725
transform 1 0 419244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4557
timestamp 1676037725
transform 1 0 420348 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4563
timestamp 1676037725
transform 1 0 420900 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4565
timestamp 1676037725
transform 1 0 421084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4577
timestamp 1676037725
transform 1 0 422188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4589
timestamp 1676037725
transform 1 0 423292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4601
timestamp 1676037725
transform 1 0 424396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4613
timestamp 1676037725
transform 1 0 425500 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4619
timestamp 1676037725
transform 1 0 426052 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4621
timestamp 1676037725
transform 1 0 426236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4633
timestamp 1676037725
transform 1 0 427340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4645
timestamp 1676037725
transform 1 0 428444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4657
timestamp 1676037725
transform 1 0 429548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4669
timestamp 1676037725
transform 1 0 430652 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4675
timestamp 1676037725
transform 1 0 431204 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4677
timestamp 1676037725
transform 1 0 431388 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4689
timestamp 1676037725
transform 1 0 432492 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4701
timestamp 1676037725
transform 1 0 433596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4713
timestamp 1676037725
transform 1 0 434700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4725
timestamp 1676037725
transform 1 0 435804 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4731
timestamp 1676037725
transform 1 0 436356 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4733
timestamp 1676037725
transform 1 0 436540 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4745
timestamp 1676037725
transform 1 0 437644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4757
timestamp 1676037725
transform 1 0 438748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4769
timestamp 1676037725
transform 1 0 439852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4781
timestamp 1676037725
transform 1 0 440956 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4787
timestamp 1676037725
transform 1 0 441508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4789
timestamp 1676037725
transform 1 0 441692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4801
timestamp 1676037725
transform 1 0 442796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4813
timestamp 1676037725
transform 1 0 443900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4825
timestamp 1676037725
transform 1 0 445004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4837
timestamp 1676037725
transform 1 0 446108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4843
timestamp 1676037725
transform 1 0 446660 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4845
timestamp 1676037725
transform 1 0 446844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4857
timestamp 1676037725
transform 1 0 447948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4869
timestamp 1676037725
transform 1 0 449052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4881
timestamp 1676037725
transform 1 0 450156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4893
timestamp 1676037725
transform 1 0 451260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4899
timestamp 1676037725
transform 1 0 451812 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4901
timestamp 1676037725
transform 1 0 451996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4913
timestamp 1676037725
transform 1 0 453100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4925
timestamp 1676037725
transform 1 0 454204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4937
timestamp 1676037725
transform 1 0 455308 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_4949
timestamp 1676037725
transform 1 0 456412 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_4955
timestamp 1676037725
transform 1 0 456964 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4957
timestamp 1676037725
transform 1 0 457148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4969
timestamp 1676037725
transform 1 0 458252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4981
timestamp 1676037725
transform 1 0 459356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_4993
timestamp 1676037725
transform 1 0 460460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5005
timestamp 1676037725
transform 1 0 461564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5011
timestamp 1676037725
transform 1 0 462116 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5013
timestamp 1676037725
transform 1 0 462300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5025
timestamp 1676037725
transform 1 0 463404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5037
timestamp 1676037725
transform 1 0 464508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5049
timestamp 1676037725
transform 1 0 465612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5061
timestamp 1676037725
transform 1 0 466716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5067
timestamp 1676037725
transform 1 0 467268 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5069
timestamp 1676037725
transform 1 0 467452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5081
timestamp 1676037725
transform 1 0 468556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5093
timestamp 1676037725
transform 1 0 469660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5105
timestamp 1676037725
transform 1 0 470764 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5117
timestamp 1676037725
transform 1 0 471868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5123
timestamp 1676037725
transform 1 0 472420 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5125
timestamp 1676037725
transform 1 0 472604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5137
timestamp 1676037725
transform 1 0 473708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5149
timestamp 1676037725
transform 1 0 474812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5161
timestamp 1676037725
transform 1 0 475916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5173
timestamp 1676037725
transform 1 0 477020 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5179
timestamp 1676037725
transform 1 0 477572 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5181
timestamp 1676037725
transform 1 0 477756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5193
timestamp 1676037725
transform 1 0 478860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5205
timestamp 1676037725
transform 1 0 479964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5217
timestamp 1676037725
transform 1 0 481068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5229
timestamp 1676037725
transform 1 0 482172 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5235
timestamp 1676037725
transform 1 0 482724 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5237
timestamp 1676037725
transform 1 0 482908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5249
timestamp 1676037725
transform 1 0 484012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5261
timestamp 1676037725
transform 1 0 485116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5273
timestamp 1676037725
transform 1 0 486220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5285
timestamp 1676037725
transform 1 0 487324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5291
timestamp 1676037725
transform 1 0 487876 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5293
timestamp 1676037725
transform 1 0 488060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5305
timestamp 1676037725
transform 1 0 489164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5317
timestamp 1676037725
transform 1 0 490268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5329
timestamp 1676037725
transform 1 0 491372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5341
timestamp 1676037725
transform 1 0 492476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5347
timestamp 1676037725
transform 1 0 493028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5349
timestamp 1676037725
transform 1 0 493212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5361
timestamp 1676037725
transform 1 0 494316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5373
timestamp 1676037725
transform 1 0 495420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5385
timestamp 1676037725
transform 1 0 496524 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5397
timestamp 1676037725
transform 1 0 497628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5403
timestamp 1676037725
transform 1 0 498180 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5405
timestamp 1676037725
transform 1 0 498364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5417
timestamp 1676037725
transform 1 0 499468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5429
timestamp 1676037725
transform 1 0 500572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5441
timestamp 1676037725
transform 1 0 501676 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5453
timestamp 1676037725
transform 1 0 502780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5459
timestamp 1676037725
transform 1 0 503332 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5461
timestamp 1676037725
transform 1 0 503516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5473
timestamp 1676037725
transform 1 0 504620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5485
timestamp 1676037725
transform 1 0 505724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5497
timestamp 1676037725
transform 1 0 506828 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5509
timestamp 1676037725
transform 1 0 507932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5515
timestamp 1676037725
transform 1 0 508484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5517
timestamp 1676037725
transform 1 0 508668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5529
timestamp 1676037725
transform 1 0 509772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5541
timestamp 1676037725
transform 1 0 510876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5553
timestamp 1676037725
transform 1 0 511980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5565
timestamp 1676037725
transform 1 0 513084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5571
timestamp 1676037725
transform 1 0 513636 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5573
timestamp 1676037725
transform 1 0 513820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5585
timestamp 1676037725
transform 1 0 514924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5597
timestamp 1676037725
transform 1 0 516028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5609
timestamp 1676037725
transform 1 0 517132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5621
timestamp 1676037725
transform 1 0 518236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5627
timestamp 1676037725
transform 1 0 518788 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5629
timestamp 1676037725
transform 1 0 518972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5641
timestamp 1676037725
transform 1 0 520076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5653
timestamp 1676037725
transform 1 0 521180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5665
timestamp 1676037725
transform 1 0 522284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_5677
timestamp 1676037725
transform 1 0 523388 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5683
timestamp 1676037725
transform 1 0 523940 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5685
timestamp 1676037725
transform 1 0 524124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5697
timestamp 1676037725
transform 1 0 525228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5709
timestamp 1676037725
transform 1 0 526332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5721
timestamp 1676037725
transform 1 0 527436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1676037725
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1676037725
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1676037725
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1676037725
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1676037725
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1676037725
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1676037725
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1676037725
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1676037725
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1676037725
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1676037725
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1676037725
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1676037725
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1676037725
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1676037725
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1676037725
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1676037725
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1676037725
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1676037725
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1676037725
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1676037725
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1676037725
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1676037725
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1676037725
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1676037725
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1676037725
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1676037725
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1676037725
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1676037725
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1676037725
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1676037725
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1676037725
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1676037725
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1676037725
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1676037725
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1676037725
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1676037725
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1676037725
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1676037725
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1676037725
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1676037725
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1676037725
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1676037725
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1676037725
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1009
timestamp 1676037725
transform 1 0 93932 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1015
timestamp 1676037725
transform 1 0 94484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1027
timestamp 1676037725
transform 1 0 95588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1035
timestamp 1676037725
transform 1 0 96324 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1040
timestamp 1676037725
transform 1 0 96784 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1052
timestamp 1676037725
transform 1 0 97888 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1062
timestamp 1676037725
transform 1 0 98808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1065
timestamp 1676037725
transform 1 0 99084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1076
timestamp 1676037725
transform 1 0 100096 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1082
timestamp 1676037725
transform 1 0 100648 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1085
timestamp 1676037725
transform 1 0 100924 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1098
timestamp 1676037725
transform 1 0 102120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1102
timestamp 1676037725
transform 1 0 102488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1105
timestamp 1676037725
transform 1 0 102764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1118
timestamp 1676037725
transform 1 0 103960 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1121
timestamp 1676037725
transform 1 0 104236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1125
timestamp 1676037725
transform 1 0 104604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1129
timestamp 1676037725
transform 1 0 104972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1132
timestamp 1676037725
transform 1 0 105248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1145
timestamp 1676037725
transform 1 0 106444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1158
timestamp 1676037725
transform 1 0 107640 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1164
timestamp 1676037725
transform 1 0 108192 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1177
timestamp 1676037725
transform 1 0 109388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1183
timestamp 1676037725
transform 1 0 109940 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1196
timestamp 1676037725
transform 1 0 111136 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1204
timestamp 1676037725
transform 1 0 111872 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1217
timestamp 1676037725
transform 1 0 113068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1230
timestamp 1676037725
transform 1 0 114264 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1233
timestamp 1676037725
transform 1 0 114540 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1237
timestamp 1676037725
transform 1 0 114908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1249
timestamp 1676037725
transform 1 0 116012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1261
timestamp 1676037725
transform 1 0 117116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1265
timestamp 1676037725
transform 1 0 117484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1268
timestamp 1676037725
transform 1 0 117760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1281
timestamp 1676037725
transform 1 0 118956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1287
timestamp 1676037725
transform 1 0 119508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1289
timestamp 1676037725
transform 1 0 119692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1295
timestamp 1676037725
transform 1 0 120244 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1305
timestamp 1676037725
transform 1 0 121164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1318
timestamp 1676037725
transform 1 0 122360 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1326
timestamp 1676037725
transform 1 0 123096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1329
timestamp 1676037725
transform 1 0 123372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1342
timestamp 1676037725
transform 1 0 124568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1345
timestamp 1676037725
transform 1 0 124844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1356
timestamp 1676037725
transform 1 0 125856 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1366
timestamp 1676037725
transform 1 0 126776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1379
timestamp 1676037725
transform 1 0 127972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1392
timestamp 1676037725
transform 1 0 129168 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1401
timestamp 1676037725
transform 1 0 129996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1413
timestamp 1676037725
transform 1 0 131100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1417
timestamp 1676037725
transform 1 0 131468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1420
timestamp 1676037725
transform 1 0 131744 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1432
timestamp 1676037725
transform 1 0 132848 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1444
timestamp 1676037725
transform 1 0 133952 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1457
timestamp 1676037725
transform 1 0 135148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1469
timestamp 1676037725
transform 1 0 136252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1481
timestamp 1676037725
transform 1 0 137356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1493
timestamp 1676037725
transform 1 0 138460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1505
timestamp 1676037725
transform 1 0 139564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1511
timestamp 1676037725
transform 1 0 140116 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1513
timestamp 1676037725
transform 1 0 140300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1525
timestamp 1676037725
transform 1 0 141404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1537
timestamp 1676037725
transform 1 0 142508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1549
timestamp 1676037725
transform 1 0 143612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1561
timestamp 1676037725
transform 1 0 144716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1567
timestamp 1676037725
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1569
timestamp 1676037725
transform 1 0 145452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1581
timestamp 1676037725
transform 1 0 146556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1593
timestamp 1676037725
transform 1 0 147660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1605
timestamp 1676037725
transform 1 0 148764 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1617
timestamp 1676037725
transform 1 0 149868 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1623
timestamp 1676037725
transform 1 0 150420 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1625
timestamp 1676037725
transform 1 0 150604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1637
timestamp 1676037725
transform 1 0 151708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1649
timestamp 1676037725
transform 1 0 152812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1661
timestamp 1676037725
transform 1 0 153916 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1673
timestamp 1676037725
transform 1 0 155020 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1679
timestamp 1676037725
transform 1 0 155572 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1681
timestamp 1676037725
transform 1 0 155756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1693
timestamp 1676037725
transform 1 0 156860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1705
timestamp 1676037725
transform 1 0 157964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1717
timestamp 1676037725
transform 1 0 159068 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1729
timestamp 1676037725
transform 1 0 160172 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1735
timestamp 1676037725
transform 1 0 160724 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1737
timestamp 1676037725
transform 1 0 160908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1749
timestamp 1676037725
transform 1 0 162012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1761
timestamp 1676037725
transform 1 0 163116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1773
timestamp 1676037725
transform 1 0 164220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1785
timestamp 1676037725
transform 1 0 165324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1791
timestamp 1676037725
transform 1 0 165876 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1793
timestamp 1676037725
transform 1 0 166060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1805
timestamp 1676037725
transform 1 0 167164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1817
timestamp 1676037725
transform 1 0 168268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1829
timestamp 1676037725
transform 1 0 169372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1841
timestamp 1676037725
transform 1 0 170476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1847
timestamp 1676037725
transform 1 0 171028 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1849
timestamp 1676037725
transform 1 0 171212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1861
timestamp 1676037725
transform 1 0 172316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1873
timestamp 1676037725
transform 1 0 173420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1885
timestamp 1676037725
transform 1 0 174524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1897
timestamp 1676037725
transform 1 0 175628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1903
timestamp 1676037725
transform 1 0 176180 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1905
timestamp 1676037725
transform 1 0 176364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1917
timestamp 1676037725
transform 1 0 177468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1929
timestamp 1676037725
transform 1 0 178572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1941
timestamp 1676037725
transform 1 0 179676 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1953
timestamp 1676037725
transform 1 0 180780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1959
timestamp 1676037725
transform 1 0 181332 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1961
timestamp 1676037725
transform 1 0 181516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1973
timestamp 1676037725
transform 1 0 182620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1985
timestamp 1676037725
transform 1 0 183724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1997
timestamp 1676037725
transform 1 0 184828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2009
timestamp 1676037725
transform 1 0 185932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2015
timestamp 1676037725
transform 1 0 186484 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2017
timestamp 1676037725
transform 1 0 186668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2029
timestamp 1676037725
transform 1 0 187772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2041
timestamp 1676037725
transform 1 0 188876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2053
timestamp 1676037725
transform 1 0 189980 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2065
timestamp 1676037725
transform 1 0 191084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2071
timestamp 1676037725
transform 1 0 191636 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2073
timestamp 1676037725
transform 1 0 191820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2085
timestamp 1676037725
transform 1 0 192924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2097
timestamp 1676037725
transform 1 0 194028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2109
timestamp 1676037725
transform 1 0 195132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2121
timestamp 1676037725
transform 1 0 196236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2127
timestamp 1676037725
transform 1 0 196788 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2129
timestamp 1676037725
transform 1 0 196972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2141
timestamp 1676037725
transform 1 0 198076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2153
timestamp 1676037725
transform 1 0 199180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2165
timestamp 1676037725
transform 1 0 200284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2177
timestamp 1676037725
transform 1 0 201388 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2183
timestamp 1676037725
transform 1 0 201940 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2185
timestamp 1676037725
transform 1 0 202124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2197
timestamp 1676037725
transform 1 0 203228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2209
timestamp 1676037725
transform 1 0 204332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2221
timestamp 1676037725
transform 1 0 205436 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2233
timestamp 1676037725
transform 1 0 206540 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2239
timestamp 1676037725
transform 1 0 207092 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2241
timestamp 1676037725
transform 1 0 207276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2253
timestamp 1676037725
transform 1 0 208380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2265
timestamp 1676037725
transform 1 0 209484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2277
timestamp 1676037725
transform 1 0 210588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2289
timestamp 1676037725
transform 1 0 211692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2295
timestamp 1676037725
transform 1 0 212244 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2297
timestamp 1676037725
transform 1 0 212428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2309
timestamp 1676037725
transform 1 0 213532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2321
timestamp 1676037725
transform 1 0 214636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2333
timestamp 1676037725
transform 1 0 215740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2345
timestamp 1676037725
transform 1 0 216844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2351
timestamp 1676037725
transform 1 0 217396 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2353
timestamp 1676037725
transform 1 0 217580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2365
timestamp 1676037725
transform 1 0 218684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2377
timestamp 1676037725
transform 1 0 219788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2389
timestamp 1676037725
transform 1 0 220892 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2401
timestamp 1676037725
transform 1 0 221996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2407
timestamp 1676037725
transform 1 0 222548 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2409
timestamp 1676037725
transform 1 0 222732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2421
timestamp 1676037725
transform 1 0 223836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2433
timestamp 1676037725
transform 1 0 224940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2445
timestamp 1676037725
transform 1 0 226044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2457
timestamp 1676037725
transform 1 0 227148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2463
timestamp 1676037725
transform 1 0 227700 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2465
timestamp 1676037725
transform 1 0 227884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2477
timestamp 1676037725
transform 1 0 228988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2489
timestamp 1676037725
transform 1 0 230092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2501
timestamp 1676037725
transform 1 0 231196 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2513
timestamp 1676037725
transform 1 0 232300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2519
timestamp 1676037725
transform 1 0 232852 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2521
timestamp 1676037725
transform 1 0 233036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2533
timestamp 1676037725
transform 1 0 234140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2545
timestamp 1676037725
transform 1 0 235244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2557
timestamp 1676037725
transform 1 0 236348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2569
timestamp 1676037725
transform 1 0 237452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2575
timestamp 1676037725
transform 1 0 238004 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2577
timestamp 1676037725
transform 1 0 238188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2589
timestamp 1676037725
transform 1 0 239292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2601
timestamp 1676037725
transform 1 0 240396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2613
timestamp 1676037725
transform 1 0 241500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2625
timestamp 1676037725
transform 1 0 242604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2631
timestamp 1676037725
transform 1 0 243156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2633
timestamp 1676037725
transform 1 0 243340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2645
timestamp 1676037725
transform 1 0 244444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2657
timestamp 1676037725
transform 1 0 245548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2669
timestamp 1676037725
transform 1 0 246652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2681
timestamp 1676037725
transform 1 0 247756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2687
timestamp 1676037725
transform 1 0 248308 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2689
timestamp 1676037725
transform 1 0 248492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2701
timestamp 1676037725
transform 1 0 249596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2713
timestamp 1676037725
transform 1 0 250700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2725
timestamp 1676037725
transform 1 0 251804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2737
timestamp 1676037725
transform 1 0 252908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2743
timestamp 1676037725
transform 1 0 253460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2745
timestamp 1676037725
transform 1 0 253644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2757
timestamp 1676037725
transform 1 0 254748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2769
timestamp 1676037725
transform 1 0 255852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2773
timestamp 1676037725
transform 1 0 256220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_2776
timestamp 1676037725
transform 1 0 256496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_2784
timestamp 1676037725
transform 1 0 257232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_2789
timestamp 1676037725
transform 1 0 257692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_2797
timestamp 1676037725
transform 1 0 258428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_2801
timestamp 1676037725
transform 1 0 258796 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_2805
timestamp 1676037725
transform 1 0 259164 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2815
timestamp 1676037725
transform 1 0 260084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2821
timestamp 1676037725
transform 1 0 260636 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2824
timestamp 1676037725
transform 1 0 260912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2837
timestamp 1676037725
transform 1 0 262108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2850
timestamp 1676037725
transform 1 0 263304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2857
timestamp 1676037725
transform 1 0 263948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2863
timestamp 1676037725
transform 1 0 264500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_2876
timestamp 1676037725
transform 1 0 265696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2880
timestamp 1676037725
transform 1 0 266064 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2890
timestamp 1676037725
transform 1 0 266984 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_2902
timestamp 1676037725
transform 1 0 268088 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_2910
timestamp 1676037725
transform 1 0 268824 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2913
timestamp 1676037725
transform 1 0 269100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2925
timestamp 1676037725
transform 1 0 270204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2937
timestamp 1676037725
transform 1 0 271308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2949
timestamp 1676037725
transform 1 0 272412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_2961
timestamp 1676037725
transform 1 0 273516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_2967
timestamp 1676037725
transform 1 0 274068 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2969
timestamp 1676037725
transform 1 0 274252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2981
timestamp 1676037725
transform 1 0 275356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_2993
timestamp 1676037725
transform 1 0 276460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3005
timestamp 1676037725
transform 1 0 277564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3017
timestamp 1676037725
transform 1 0 278668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3023
timestamp 1676037725
transform 1 0 279220 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3025
timestamp 1676037725
transform 1 0 279404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3037
timestamp 1676037725
transform 1 0 280508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3049
timestamp 1676037725
transform 1 0 281612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3061
timestamp 1676037725
transform 1 0 282716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3073
timestamp 1676037725
transform 1 0 283820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3079
timestamp 1676037725
transform 1 0 284372 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3081
timestamp 1676037725
transform 1 0 284556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3093
timestamp 1676037725
transform 1 0 285660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3105
timestamp 1676037725
transform 1 0 286764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3117
timestamp 1676037725
transform 1 0 287868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3129
timestamp 1676037725
transform 1 0 288972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3135
timestamp 1676037725
transform 1 0 289524 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3137
timestamp 1676037725
transform 1 0 289708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3149
timestamp 1676037725
transform 1 0 290812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3161
timestamp 1676037725
transform 1 0 291916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3173
timestamp 1676037725
transform 1 0 293020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3185
timestamp 1676037725
transform 1 0 294124 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3191
timestamp 1676037725
transform 1 0 294676 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3193
timestamp 1676037725
transform 1 0 294860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3205
timestamp 1676037725
transform 1 0 295964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3217
timestamp 1676037725
transform 1 0 297068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3229
timestamp 1676037725
transform 1 0 298172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3241
timestamp 1676037725
transform 1 0 299276 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3247
timestamp 1676037725
transform 1 0 299828 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3249
timestamp 1676037725
transform 1 0 300012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3261
timestamp 1676037725
transform 1 0 301116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3273
timestamp 1676037725
transform 1 0 302220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3285
timestamp 1676037725
transform 1 0 303324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3297
timestamp 1676037725
transform 1 0 304428 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3303
timestamp 1676037725
transform 1 0 304980 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3305
timestamp 1676037725
transform 1 0 305164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3317
timestamp 1676037725
transform 1 0 306268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3329
timestamp 1676037725
transform 1 0 307372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3341
timestamp 1676037725
transform 1 0 308476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3353
timestamp 1676037725
transform 1 0 309580 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3359
timestamp 1676037725
transform 1 0 310132 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3361
timestamp 1676037725
transform 1 0 310316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3373
timestamp 1676037725
transform 1 0 311420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3385
timestamp 1676037725
transform 1 0 312524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3397
timestamp 1676037725
transform 1 0 313628 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3409
timestamp 1676037725
transform 1 0 314732 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3415
timestamp 1676037725
transform 1 0 315284 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3417
timestamp 1676037725
transform 1 0 315468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3429
timestamp 1676037725
transform 1 0 316572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3441
timestamp 1676037725
transform 1 0 317676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3453
timestamp 1676037725
transform 1 0 318780 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3465
timestamp 1676037725
transform 1 0 319884 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3471
timestamp 1676037725
transform 1 0 320436 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3473
timestamp 1676037725
transform 1 0 320620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3485
timestamp 1676037725
transform 1 0 321724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3497
timestamp 1676037725
transform 1 0 322828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3509
timestamp 1676037725
transform 1 0 323932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3521
timestamp 1676037725
transform 1 0 325036 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3527
timestamp 1676037725
transform 1 0 325588 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3529
timestamp 1676037725
transform 1 0 325772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3541
timestamp 1676037725
transform 1 0 326876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3553
timestamp 1676037725
transform 1 0 327980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3565
timestamp 1676037725
transform 1 0 329084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3577
timestamp 1676037725
transform 1 0 330188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3583
timestamp 1676037725
transform 1 0 330740 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3585
timestamp 1676037725
transform 1 0 330924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3597
timestamp 1676037725
transform 1 0 332028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3609
timestamp 1676037725
transform 1 0 333132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3621
timestamp 1676037725
transform 1 0 334236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3633
timestamp 1676037725
transform 1 0 335340 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3639
timestamp 1676037725
transform 1 0 335892 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3641
timestamp 1676037725
transform 1 0 336076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3653
timestamp 1676037725
transform 1 0 337180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3665
timestamp 1676037725
transform 1 0 338284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3677
timestamp 1676037725
transform 1 0 339388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3689
timestamp 1676037725
transform 1 0 340492 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3695
timestamp 1676037725
transform 1 0 341044 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3697
timestamp 1676037725
transform 1 0 341228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3709
timestamp 1676037725
transform 1 0 342332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3721
timestamp 1676037725
transform 1 0 343436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3733
timestamp 1676037725
transform 1 0 344540 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3745
timestamp 1676037725
transform 1 0 345644 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3751
timestamp 1676037725
transform 1 0 346196 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3753
timestamp 1676037725
transform 1 0 346380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3765
timestamp 1676037725
transform 1 0 347484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3777
timestamp 1676037725
transform 1 0 348588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3789
timestamp 1676037725
transform 1 0 349692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3801
timestamp 1676037725
transform 1 0 350796 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3807
timestamp 1676037725
transform 1 0 351348 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3809
timestamp 1676037725
transform 1 0 351532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3821
timestamp 1676037725
transform 1 0 352636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3833
timestamp 1676037725
transform 1 0 353740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3845
timestamp 1676037725
transform 1 0 354844 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3857
timestamp 1676037725
transform 1 0 355948 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3863
timestamp 1676037725
transform 1 0 356500 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3865
timestamp 1676037725
transform 1 0 356684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3877
timestamp 1676037725
transform 1 0 357788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3889
timestamp 1676037725
transform 1 0 358892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3901
timestamp 1676037725
transform 1 0 359996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3913
timestamp 1676037725
transform 1 0 361100 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3919
timestamp 1676037725
transform 1 0 361652 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3921
timestamp 1676037725
transform 1 0 361836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3933
timestamp 1676037725
transform 1 0 362940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3945
timestamp 1676037725
transform 1 0 364044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3957
timestamp 1676037725
transform 1 0 365148 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3969
timestamp 1676037725
transform 1 0 366252 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3975
timestamp 1676037725
transform 1 0 366804 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3977
timestamp 1676037725
transform 1 0 366988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3989
timestamp 1676037725
transform 1 0 368092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4001
timestamp 1676037725
transform 1 0 369196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4013
timestamp 1676037725
transform 1 0 370300 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4025
timestamp 1676037725
transform 1 0 371404 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4031
timestamp 1676037725
transform 1 0 371956 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4033
timestamp 1676037725
transform 1 0 372140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4045
timestamp 1676037725
transform 1 0 373244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4057
timestamp 1676037725
transform 1 0 374348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4069
timestamp 1676037725
transform 1 0 375452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4081
timestamp 1676037725
transform 1 0 376556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4087
timestamp 1676037725
transform 1 0 377108 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4089
timestamp 1676037725
transform 1 0 377292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4101
timestamp 1676037725
transform 1 0 378396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4113
timestamp 1676037725
transform 1 0 379500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4125
timestamp 1676037725
transform 1 0 380604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4137
timestamp 1676037725
transform 1 0 381708 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4143
timestamp 1676037725
transform 1 0 382260 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4145
timestamp 1676037725
transform 1 0 382444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4157
timestamp 1676037725
transform 1 0 383548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4169
timestamp 1676037725
transform 1 0 384652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4181
timestamp 1676037725
transform 1 0 385756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4193
timestamp 1676037725
transform 1 0 386860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4199
timestamp 1676037725
transform 1 0 387412 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4201
timestamp 1676037725
transform 1 0 387596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4213
timestamp 1676037725
transform 1 0 388700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4225
timestamp 1676037725
transform 1 0 389804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4237
timestamp 1676037725
transform 1 0 390908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4249
timestamp 1676037725
transform 1 0 392012 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4255
timestamp 1676037725
transform 1 0 392564 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4257
timestamp 1676037725
transform 1 0 392748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4269
timestamp 1676037725
transform 1 0 393852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4281
timestamp 1676037725
transform 1 0 394956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4293
timestamp 1676037725
transform 1 0 396060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4305
timestamp 1676037725
transform 1 0 397164 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4311
timestamp 1676037725
transform 1 0 397716 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4313
timestamp 1676037725
transform 1 0 397900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4325
timestamp 1676037725
transform 1 0 399004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4337
timestamp 1676037725
transform 1 0 400108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4349
timestamp 1676037725
transform 1 0 401212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4361
timestamp 1676037725
transform 1 0 402316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4367
timestamp 1676037725
transform 1 0 402868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4369
timestamp 1676037725
transform 1 0 403052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4381
timestamp 1676037725
transform 1 0 404156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4393
timestamp 1676037725
transform 1 0 405260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4405
timestamp 1676037725
transform 1 0 406364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4417
timestamp 1676037725
transform 1 0 407468 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4423
timestamp 1676037725
transform 1 0 408020 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4425
timestamp 1676037725
transform 1 0 408204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4437
timestamp 1676037725
transform 1 0 409308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4449
timestamp 1676037725
transform 1 0 410412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4461
timestamp 1676037725
transform 1 0 411516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4473
timestamp 1676037725
transform 1 0 412620 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4479
timestamp 1676037725
transform 1 0 413172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4481
timestamp 1676037725
transform 1 0 413356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4493
timestamp 1676037725
transform 1 0 414460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4505
timestamp 1676037725
transform 1 0 415564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4517
timestamp 1676037725
transform 1 0 416668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4529
timestamp 1676037725
transform 1 0 417772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4535
timestamp 1676037725
transform 1 0 418324 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4537
timestamp 1676037725
transform 1 0 418508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4549
timestamp 1676037725
transform 1 0 419612 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4561
timestamp 1676037725
transform 1 0 420716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4573
timestamp 1676037725
transform 1 0 421820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4585
timestamp 1676037725
transform 1 0 422924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4591
timestamp 1676037725
transform 1 0 423476 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4593
timestamp 1676037725
transform 1 0 423660 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4605
timestamp 1676037725
transform 1 0 424764 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4617
timestamp 1676037725
transform 1 0 425868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4629
timestamp 1676037725
transform 1 0 426972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4641
timestamp 1676037725
transform 1 0 428076 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4647
timestamp 1676037725
transform 1 0 428628 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4649
timestamp 1676037725
transform 1 0 428812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4661
timestamp 1676037725
transform 1 0 429916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4673
timestamp 1676037725
transform 1 0 431020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4685
timestamp 1676037725
transform 1 0 432124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4697
timestamp 1676037725
transform 1 0 433228 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4703
timestamp 1676037725
transform 1 0 433780 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4705
timestamp 1676037725
transform 1 0 433964 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4717
timestamp 1676037725
transform 1 0 435068 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4729
timestamp 1676037725
transform 1 0 436172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4741
timestamp 1676037725
transform 1 0 437276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4753
timestamp 1676037725
transform 1 0 438380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4759
timestamp 1676037725
transform 1 0 438932 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4761
timestamp 1676037725
transform 1 0 439116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4773
timestamp 1676037725
transform 1 0 440220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4785
timestamp 1676037725
transform 1 0 441324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4797
timestamp 1676037725
transform 1 0 442428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4809
timestamp 1676037725
transform 1 0 443532 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4815
timestamp 1676037725
transform 1 0 444084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4817
timestamp 1676037725
transform 1 0 444268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4829
timestamp 1676037725
transform 1 0 445372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4841
timestamp 1676037725
transform 1 0 446476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4853
timestamp 1676037725
transform 1 0 447580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4865
timestamp 1676037725
transform 1 0 448684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4871
timestamp 1676037725
transform 1 0 449236 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4873
timestamp 1676037725
transform 1 0 449420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4885
timestamp 1676037725
transform 1 0 450524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4897
timestamp 1676037725
transform 1 0 451628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4909
timestamp 1676037725
transform 1 0 452732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4921
timestamp 1676037725
transform 1 0 453836 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4927
timestamp 1676037725
transform 1 0 454388 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4929
timestamp 1676037725
transform 1 0 454572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4941
timestamp 1676037725
transform 1 0 455676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4953
timestamp 1676037725
transform 1 0 456780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4965
timestamp 1676037725
transform 1 0 457884 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_4977
timestamp 1676037725
transform 1 0 458988 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_4983
timestamp 1676037725
transform 1 0 459540 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4985
timestamp 1676037725
transform 1 0 459724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_4997
timestamp 1676037725
transform 1 0 460828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5009
timestamp 1676037725
transform 1 0 461932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5021
timestamp 1676037725
transform 1 0 463036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5033
timestamp 1676037725
transform 1 0 464140 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5039
timestamp 1676037725
transform 1 0 464692 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5041
timestamp 1676037725
transform 1 0 464876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5053
timestamp 1676037725
transform 1 0 465980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5065
timestamp 1676037725
transform 1 0 467084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5077
timestamp 1676037725
transform 1 0 468188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5089
timestamp 1676037725
transform 1 0 469292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5095
timestamp 1676037725
transform 1 0 469844 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5097
timestamp 1676037725
transform 1 0 470028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5109
timestamp 1676037725
transform 1 0 471132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5121
timestamp 1676037725
transform 1 0 472236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5133
timestamp 1676037725
transform 1 0 473340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5145
timestamp 1676037725
transform 1 0 474444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5151
timestamp 1676037725
transform 1 0 474996 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5153
timestamp 1676037725
transform 1 0 475180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5165
timestamp 1676037725
transform 1 0 476284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5177
timestamp 1676037725
transform 1 0 477388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5189
timestamp 1676037725
transform 1 0 478492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5201
timestamp 1676037725
transform 1 0 479596 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5207
timestamp 1676037725
transform 1 0 480148 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5209
timestamp 1676037725
transform 1 0 480332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5221
timestamp 1676037725
transform 1 0 481436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5233
timestamp 1676037725
transform 1 0 482540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5245
timestamp 1676037725
transform 1 0 483644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5257
timestamp 1676037725
transform 1 0 484748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5263
timestamp 1676037725
transform 1 0 485300 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5265
timestamp 1676037725
transform 1 0 485484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5277
timestamp 1676037725
transform 1 0 486588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5289
timestamp 1676037725
transform 1 0 487692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5301
timestamp 1676037725
transform 1 0 488796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5313
timestamp 1676037725
transform 1 0 489900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5319
timestamp 1676037725
transform 1 0 490452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5321
timestamp 1676037725
transform 1 0 490636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5333
timestamp 1676037725
transform 1 0 491740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5345
timestamp 1676037725
transform 1 0 492844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5357
timestamp 1676037725
transform 1 0 493948 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5369
timestamp 1676037725
transform 1 0 495052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5375
timestamp 1676037725
transform 1 0 495604 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5377
timestamp 1676037725
transform 1 0 495788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5389
timestamp 1676037725
transform 1 0 496892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5401
timestamp 1676037725
transform 1 0 497996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5413
timestamp 1676037725
transform 1 0 499100 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5425
timestamp 1676037725
transform 1 0 500204 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5431
timestamp 1676037725
transform 1 0 500756 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5433
timestamp 1676037725
transform 1 0 500940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5445
timestamp 1676037725
transform 1 0 502044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5457
timestamp 1676037725
transform 1 0 503148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5469
timestamp 1676037725
transform 1 0 504252 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5481
timestamp 1676037725
transform 1 0 505356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5487
timestamp 1676037725
transform 1 0 505908 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5489
timestamp 1676037725
transform 1 0 506092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5501
timestamp 1676037725
transform 1 0 507196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5513
timestamp 1676037725
transform 1 0 508300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5525
timestamp 1676037725
transform 1 0 509404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5537
timestamp 1676037725
transform 1 0 510508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5543
timestamp 1676037725
transform 1 0 511060 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5545
timestamp 1676037725
transform 1 0 511244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5557
timestamp 1676037725
transform 1 0 512348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5569
timestamp 1676037725
transform 1 0 513452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5581
timestamp 1676037725
transform 1 0 514556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5593
timestamp 1676037725
transform 1 0 515660 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5599
timestamp 1676037725
transform 1 0 516212 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5601
timestamp 1676037725
transform 1 0 516396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5613
timestamp 1676037725
transform 1 0 517500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5625
timestamp 1676037725
transform 1 0 518604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5637
timestamp 1676037725
transform 1 0 519708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5649
timestamp 1676037725
transform 1 0 520812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5655
timestamp 1676037725
transform 1 0 521364 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5657
timestamp 1676037725
transform 1 0 521548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5669
timestamp 1676037725
transform 1 0 522652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5681
timestamp 1676037725
transform 1 0 523756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5693
timestamp 1676037725
transform 1 0 524860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_5705
timestamp 1676037725
transform 1 0 525964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_5711
timestamp 1676037725
transform 1 0 526516 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_5713
timestamp 1676037725
transform 1 0 526700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_5725
timestamp 1676037725
transform 1 0 527804 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1676037725
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1676037725
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1676037725
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1676037725
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1676037725
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1676037725
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1676037725
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1676037725
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1676037725
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1676037725
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1676037725
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1676037725
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1676037725
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1676037725
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1676037725
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1676037725
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1676037725
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1676037725
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1676037725
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1676037725
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1676037725
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1676037725
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1676037725
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1676037725
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1676037725
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1676037725
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1676037725
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1676037725
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1676037725
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1676037725
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1676037725
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1676037725
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1676037725
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1676037725
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1676037725
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1676037725
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1676037725
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1676037725
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1676037725
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_973
timestamp 1676037725
transform 1 0 90620 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_978
timestamp 1676037725
transform 1 0 91080 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_981
timestamp 1676037725
transform 1 0 91356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_992
timestamp 1676037725
transform 1 0 92368 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_998
timestamp 1676037725
transform 1 0 92920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1011
timestamp 1676037725
transform 1 0 94116 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1024
timestamp 1676037725
transform 1 0 95312 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1037
timestamp 1676037725
transform 1 0 96508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1049
timestamp 1676037725
transform 1 0 97612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1059
timestamp 1676037725
transform 1 0 98532 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1072
timestamp 1676037725
transform 1 0 99728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1084
timestamp 1676037725
transform 1 0 100832 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1090
timestamp 1676037725
transform 1 0 101384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1093
timestamp 1676037725
transform 1 0 101660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1108
timestamp 1676037725
transform 1 0 103040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1121
timestamp 1676037725
transform 1 0 104236 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1134
timestamp 1676037725
transform 1 0 105432 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1146
timestamp 1676037725
transform 1 0 106536 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1149
timestamp 1676037725
transform 1 0 106812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1157
timestamp 1676037725
transform 1 0 107548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1170
timestamp 1676037725
transform 1 0 108744 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1178
timestamp 1676037725
transform 1 0 109480 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1182
timestamp 1676037725
transform 1 0 109848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1195
timestamp 1676037725
transform 1 0 111044 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1199
timestamp 1676037725
transform 1 0 111412 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1202
timestamp 1676037725
transform 1 0 111688 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1205
timestamp 1676037725
transform 1 0 111964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1216
timestamp 1676037725
transform 1 0 112976 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1231
timestamp 1676037725
transform 1 0 114356 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1244
timestamp 1676037725
transform 1 0 115552 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1258
timestamp 1676037725
transform 1 0 116840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1261
timestamp 1676037725
transform 1 0 117116 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1272
timestamp 1676037725
transform 1 0 118128 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1284
timestamp 1676037725
transform 1 0 119232 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_1292
timestamp 1676037725
transform 1 0 119968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1296
timestamp 1676037725
transform 1 0 120336 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1304
timestamp 1676037725
transform 1 0 121072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1309
timestamp 1676037725
transform 1 0 121532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1315
timestamp 1676037725
transform 1 0 122084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1317
timestamp 1676037725
transform 1 0 122268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1329
timestamp 1676037725
transform 1 0 123372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1341
timestamp 1676037725
transform 1 0 124476 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1347
timestamp 1676037725
transform 1 0 125028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1359
timestamp 1676037725
transform 1 0 126132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1371
timestamp 1676037725
transform 1 0 127236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1373
timestamp 1676037725
transform 1 0 127420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1385
timestamp 1676037725
transform 1 0 128524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1397
timestamp 1676037725
transform 1 0 129628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1409
timestamp 1676037725
transform 1 0 130732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1421
timestamp 1676037725
transform 1 0 131836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1427
timestamp 1676037725
transform 1 0 132388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1429
timestamp 1676037725
transform 1 0 132572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1441
timestamp 1676037725
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1453
timestamp 1676037725
transform 1 0 134780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1465
timestamp 1676037725
transform 1 0 135884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1477
timestamp 1676037725
transform 1 0 136988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1483
timestamp 1676037725
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1485
timestamp 1676037725
transform 1 0 137724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1497
timestamp 1676037725
transform 1 0 138828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1509
timestamp 1676037725
transform 1 0 139932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1521
timestamp 1676037725
transform 1 0 141036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1533
timestamp 1676037725
transform 1 0 142140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1539
timestamp 1676037725
transform 1 0 142692 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1541
timestamp 1676037725
transform 1 0 142876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1553
timestamp 1676037725
transform 1 0 143980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1565
timestamp 1676037725
transform 1 0 145084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1577
timestamp 1676037725
transform 1 0 146188 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1589
timestamp 1676037725
transform 1 0 147292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1595
timestamp 1676037725
transform 1 0 147844 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1597
timestamp 1676037725
transform 1 0 148028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1609
timestamp 1676037725
transform 1 0 149132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1621
timestamp 1676037725
transform 1 0 150236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1633
timestamp 1676037725
transform 1 0 151340 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1645
timestamp 1676037725
transform 1 0 152444 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1651
timestamp 1676037725
transform 1 0 152996 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1653
timestamp 1676037725
transform 1 0 153180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1665
timestamp 1676037725
transform 1 0 154284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1677
timestamp 1676037725
transform 1 0 155388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1689
timestamp 1676037725
transform 1 0 156492 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1701
timestamp 1676037725
transform 1 0 157596 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1707
timestamp 1676037725
transform 1 0 158148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1709
timestamp 1676037725
transform 1 0 158332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1721
timestamp 1676037725
transform 1 0 159436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1733
timestamp 1676037725
transform 1 0 160540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1745
timestamp 1676037725
transform 1 0 161644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1757
timestamp 1676037725
transform 1 0 162748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1763
timestamp 1676037725
transform 1 0 163300 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1765
timestamp 1676037725
transform 1 0 163484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1777
timestamp 1676037725
transform 1 0 164588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1789
timestamp 1676037725
transform 1 0 165692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1801
timestamp 1676037725
transform 1 0 166796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1813
timestamp 1676037725
transform 1 0 167900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1819
timestamp 1676037725
transform 1 0 168452 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1821
timestamp 1676037725
transform 1 0 168636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1833
timestamp 1676037725
transform 1 0 169740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1845
timestamp 1676037725
transform 1 0 170844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1857
timestamp 1676037725
transform 1 0 171948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1869
timestamp 1676037725
transform 1 0 173052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1875
timestamp 1676037725
transform 1 0 173604 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1877
timestamp 1676037725
transform 1 0 173788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1889
timestamp 1676037725
transform 1 0 174892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1901
timestamp 1676037725
transform 1 0 175996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1913
timestamp 1676037725
transform 1 0 177100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1925
timestamp 1676037725
transform 1 0 178204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1931
timestamp 1676037725
transform 1 0 178756 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1933
timestamp 1676037725
transform 1 0 178940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1945
timestamp 1676037725
transform 1 0 180044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1957
timestamp 1676037725
transform 1 0 181148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1969
timestamp 1676037725
transform 1 0 182252 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1981
timestamp 1676037725
transform 1 0 183356 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1987
timestamp 1676037725
transform 1 0 183908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1989
timestamp 1676037725
transform 1 0 184092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2001
timestamp 1676037725
transform 1 0 185196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2013
timestamp 1676037725
transform 1 0 186300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2025
timestamp 1676037725
transform 1 0 187404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2037
timestamp 1676037725
transform 1 0 188508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2043
timestamp 1676037725
transform 1 0 189060 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2045
timestamp 1676037725
transform 1 0 189244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2057
timestamp 1676037725
transform 1 0 190348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2069
timestamp 1676037725
transform 1 0 191452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2081
timestamp 1676037725
transform 1 0 192556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2093
timestamp 1676037725
transform 1 0 193660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2099
timestamp 1676037725
transform 1 0 194212 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2101
timestamp 1676037725
transform 1 0 194396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2113
timestamp 1676037725
transform 1 0 195500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2125
timestamp 1676037725
transform 1 0 196604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2137
timestamp 1676037725
transform 1 0 197708 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2149
timestamp 1676037725
transform 1 0 198812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2155
timestamp 1676037725
transform 1 0 199364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2157
timestamp 1676037725
transform 1 0 199548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2169
timestamp 1676037725
transform 1 0 200652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2181
timestamp 1676037725
transform 1 0 201756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2193
timestamp 1676037725
transform 1 0 202860 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2205
timestamp 1676037725
transform 1 0 203964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2211
timestamp 1676037725
transform 1 0 204516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2213
timestamp 1676037725
transform 1 0 204700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2225
timestamp 1676037725
transform 1 0 205804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2237
timestamp 1676037725
transform 1 0 206908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2249
timestamp 1676037725
transform 1 0 208012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2261
timestamp 1676037725
transform 1 0 209116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2267
timestamp 1676037725
transform 1 0 209668 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2269
timestamp 1676037725
transform 1 0 209852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2281
timestamp 1676037725
transform 1 0 210956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2293
timestamp 1676037725
transform 1 0 212060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2305
timestamp 1676037725
transform 1 0 213164 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2317
timestamp 1676037725
transform 1 0 214268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2323
timestamp 1676037725
transform 1 0 214820 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2325
timestamp 1676037725
transform 1 0 215004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2337
timestamp 1676037725
transform 1 0 216108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2349
timestamp 1676037725
transform 1 0 217212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2361
timestamp 1676037725
transform 1 0 218316 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2373
timestamp 1676037725
transform 1 0 219420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2379
timestamp 1676037725
transform 1 0 219972 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2381
timestamp 1676037725
transform 1 0 220156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2393
timestamp 1676037725
transform 1 0 221260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2405
timestamp 1676037725
transform 1 0 222364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2417
timestamp 1676037725
transform 1 0 223468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2429
timestamp 1676037725
transform 1 0 224572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2435
timestamp 1676037725
transform 1 0 225124 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2437
timestamp 1676037725
transform 1 0 225308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2449
timestamp 1676037725
transform 1 0 226412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2461
timestamp 1676037725
transform 1 0 227516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2473
timestamp 1676037725
transform 1 0 228620 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2485
timestamp 1676037725
transform 1 0 229724 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2491
timestamp 1676037725
transform 1 0 230276 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2493
timestamp 1676037725
transform 1 0 230460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2505
timestamp 1676037725
transform 1 0 231564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2517
timestamp 1676037725
transform 1 0 232668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2529
timestamp 1676037725
transform 1 0 233772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2541
timestamp 1676037725
transform 1 0 234876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2547
timestamp 1676037725
transform 1 0 235428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2549
timestamp 1676037725
transform 1 0 235612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2561
timestamp 1676037725
transform 1 0 236716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2573
timestamp 1676037725
transform 1 0 237820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2585
timestamp 1676037725
transform 1 0 238924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2597
timestamp 1676037725
transform 1 0 240028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2603
timestamp 1676037725
transform 1 0 240580 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2605
timestamp 1676037725
transform 1 0 240764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2617
timestamp 1676037725
transform 1 0 241868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2629
timestamp 1676037725
transform 1 0 242972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2641
timestamp 1676037725
transform 1 0 244076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2653
timestamp 1676037725
transform 1 0 245180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2659
timestamp 1676037725
transform 1 0 245732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2661
timestamp 1676037725
transform 1 0 245916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2673
timestamp 1676037725
transform 1 0 247020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2685
timestamp 1676037725
transform 1 0 248124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2697
timestamp 1676037725
transform 1 0 249228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2709
timestamp 1676037725
transform 1 0 250332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2715
timestamp 1676037725
transform 1 0 250884 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_2717
timestamp 1676037725
transform 1 0 251068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2728
timestamp 1676037725
transform 1 0 252080 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2734
timestamp 1676037725
transform 1 0 252632 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_2746
timestamp 1676037725
transform 1 0 253736 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2750
timestamp 1676037725
transform 1 0 254104 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2754
timestamp 1676037725
transform 1 0 254472 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2757
timestamp 1676037725
transform 1 0 254748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_2770
timestamp 1676037725
transform 1 0 255944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_2773
timestamp 1676037725
transform 1 0 256220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2785
timestamp 1676037725
transform 1 0 257324 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2798
timestamp 1676037725
transform 1 0 258520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2811
timestamp 1676037725
transform 1 0 259716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_2824
timestamp 1676037725
transform 1 0 260912 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2829
timestamp 1676037725
transform 1 0 261372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2841
timestamp 1676037725
transform 1 0 262476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2853
timestamp 1676037725
transform 1 0 263580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2865
timestamp 1676037725
transform 1 0 264684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2877
timestamp 1676037725
transform 1 0 265788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2883
timestamp 1676037725
transform 1 0 266340 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2885
timestamp 1676037725
transform 1 0 266524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2897
timestamp 1676037725
transform 1 0 267628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2909
timestamp 1676037725
transform 1 0 268732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2921
timestamp 1676037725
transform 1 0 269836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2933
timestamp 1676037725
transform 1 0 270940 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2939
timestamp 1676037725
transform 1 0 271492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2941
timestamp 1676037725
transform 1 0 271676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2953
timestamp 1676037725
transform 1 0 272780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2965
timestamp 1676037725
transform 1 0 273884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2977
timestamp 1676037725
transform 1 0 274988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_2989
timestamp 1676037725
transform 1 0 276092 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_2995
timestamp 1676037725
transform 1 0 276644 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_2997
timestamp 1676037725
transform 1 0 276828 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3009
timestamp 1676037725
transform 1 0 277932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3021
timestamp 1676037725
transform 1 0 279036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3033
timestamp 1676037725
transform 1 0 280140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3045
timestamp 1676037725
transform 1 0 281244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3051
timestamp 1676037725
transform 1 0 281796 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3053
timestamp 1676037725
transform 1 0 281980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3065
timestamp 1676037725
transform 1 0 283084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3077
timestamp 1676037725
transform 1 0 284188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3089
timestamp 1676037725
transform 1 0 285292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3101
timestamp 1676037725
transform 1 0 286396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3107
timestamp 1676037725
transform 1 0 286948 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3109
timestamp 1676037725
transform 1 0 287132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3121
timestamp 1676037725
transform 1 0 288236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3133
timestamp 1676037725
transform 1 0 289340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3145
timestamp 1676037725
transform 1 0 290444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3157
timestamp 1676037725
transform 1 0 291548 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3163
timestamp 1676037725
transform 1 0 292100 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3165
timestamp 1676037725
transform 1 0 292284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3177
timestamp 1676037725
transform 1 0 293388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3189
timestamp 1676037725
transform 1 0 294492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3201
timestamp 1676037725
transform 1 0 295596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3213
timestamp 1676037725
transform 1 0 296700 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3219
timestamp 1676037725
transform 1 0 297252 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3221
timestamp 1676037725
transform 1 0 297436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3233
timestamp 1676037725
transform 1 0 298540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3245
timestamp 1676037725
transform 1 0 299644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3257
timestamp 1676037725
transform 1 0 300748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3269
timestamp 1676037725
transform 1 0 301852 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3275
timestamp 1676037725
transform 1 0 302404 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3277
timestamp 1676037725
transform 1 0 302588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3289
timestamp 1676037725
transform 1 0 303692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3301
timestamp 1676037725
transform 1 0 304796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3313
timestamp 1676037725
transform 1 0 305900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3325
timestamp 1676037725
transform 1 0 307004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3331
timestamp 1676037725
transform 1 0 307556 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3333
timestamp 1676037725
transform 1 0 307740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3345
timestamp 1676037725
transform 1 0 308844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3357
timestamp 1676037725
transform 1 0 309948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3369
timestamp 1676037725
transform 1 0 311052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3381
timestamp 1676037725
transform 1 0 312156 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3387
timestamp 1676037725
transform 1 0 312708 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3389
timestamp 1676037725
transform 1 0 312892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3401
timestamp 1676037725
transform 1 0 313996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3413
timestamp 1676037725
transform 1 0 315100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3425
timestamp 1676037725
transform 1 0 316204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3437
timestamp 1676037725
transform 1 0 317308 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3443
timestamp 1676037725
transform 1 0 317860 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3445
timestamp 1676037725
transform 1 0 318044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3457
timestamp 1676037725
transform 1 0 319148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3469
timestamp 1676037725
transform 1 0 320252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3481
timestamp 1676037725
transform 1 0 321356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3493
timestamp 1676037725
transform 1 0 322460 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3499
timestamp 1676037725
transform 1 0 323012 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3501
timestamp 1676037725
transform 1 0 323196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3513
timestamp 1676037725
transform 1 0 324300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3525
timestamp 1676037725
transform 1 0 325404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3537
timestamp 1676037725
transform 1 0 326508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3549
timestamp 1676037725
transform 1 0 327612 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3555
timestamp 1676037725
transform 1 0 328164 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3557
timestamp 1676037725
transform 1 0 328348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3569
timestamp 1676037725
transform 1 0 329452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3581
timestamp 1676037725
transform 1 0 330556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3593
timestamp 1676037725
transform 1 0 331660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3605
timestamp 1676037725
transform 1 0 332764 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3611
timestamp 1676037725
transform 1 0 333316 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3613
timestamp 1676037725
transform 1 0 333500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3625
timestamp 1676037725
transform 1 0 334604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3637
timestamp 1676037725
transform 1 0 335708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3649
timestamp 1676037725
transform 1 0 336812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3661
timestamp 1676037725
transform 1 0 337916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3667
timestamp 1676037725
transform 1 0 338468 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3669
timestamp 1676037725
transform 1 0 338652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3681
timestamp 1676037725
transform 1 0 339756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3693
timestamp 1676037725
transform 1 0 340860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3705
timestamp 1676037725
transform 1 0 341964 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3717
timestamp 1676037725
transform 1 0 343068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3723
timestamp 1676037725
transform 1 0 343620 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3725
timestamp 1676037725
transform 1 0 343804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3737
timestamp 1676037725
transform 1 0 344908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3749
timestamp 1676037725
transform 1 0 346012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3761
timestamp 1676037725
transform 1 0 347116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3773
timestamp 1676037725
transform 1 0 348220 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3779
timestamp 1676037725
transform 1 0 348772 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3781
timestamp 1676037725
transform 1 0 348956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3793
timestamp 1676037725
transform 1 0 350060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3805
timestamp 1676037725
transform 1 0 351164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3817
timestamp 1676037725
transform 1 0 352268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3829
timestamp 1676037725
transform 1 0 353372 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3835
timestamp 1676037725
transform 1 0 353924 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3837
timestamp 1676037725
transform 1 0 354108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3849
timestamp 1676037725
transform 1 0 355212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3861
timestamp 1676037725
transform 1 0 356316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3873
timestamp 1676037725
transform 1 0 357420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3885
timestamp 1676037725
transform 1 0 358524 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3891
timestamp 1676037725
transform 1 0 359076 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3893
timestamp 1676037725
transform 1 0 359260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3905
timestamp 1676037725
transform 1 0 360364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3917
timestamp 1676037725
transform 1 0 361468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3929
timestamp 1676037725
transform 1 0 362572 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3941
timestamp 1676037725
transform 1 0 363676 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3947
timestamp 1676037725
transform 1 0 364228 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3949
timestamp 1676037725
transform 1 0 364412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3961
timestamp 1676037725
transform 1 0 365516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3973
timestamp 1676037725
transform 1 0 366620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3985
timestamp 1676037725
transform 1 0 367724 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3997
timestamp 1676037725
transform 1 0 368828 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4003
timestamp 1676037725
transform 1 0 369380 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4005
timestamp 1676037725
transform 1 0 369564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4017
timestamp 1676037725
transform 1 0 370668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4029
timestamp 1676037725
transform 1 0 371772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4041
timestamp 1676037725
transform 1 0 372876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4053
timestamp 1676037725
transform 1 0 373980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4059
timestamp 1676037725
transform 1 0 374532 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4061
timestamp 1676037725
transform 1 0 374716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4073
timestamp 1676037725
transform 1 0 375820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4085
timestamp 1676037725
transform 1 0 376924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4097
timestamp 1676037725
transform 1 0 378028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4109
timestamp 1676037725
transform 1 0 379132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4115
timestamp 1676037725
transform 1 0 379684 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4117
timestamp 1676037725
transform 1 0 379868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4129
timestamp 1676037725
transform 1 0 380972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4141
timestamp 1676037725
transform 1 0 382076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4153
timestamp 1676037725
transform 1 0 383180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4165
timestamp 1676037725
transform 1 0 384284 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4171
timestamp 1676037725
transform 1 0 384836 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4173
timestamp 1676037725
transform 1 0 385020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4185
timestamp 1676037725
transform 1 0 386124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4197
timestamp 1676037725
transform 1 0 387228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4209
timestamp 1676037725
transform 1 0 388332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4221
timestamp 1676037725
transform 1 0 389436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4227
timestamp 1676037725
transform 1 0 389988 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4229
timestamp 1676037725
transform 1 0 390172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4241
timestamp 1676037725
transform 1 0 391276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4253
timestamp 1676037725
transform 1 0 392380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4265
timestamp 1676037725
transform 1 0 393484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4277
timestamp 1676037725
transform 1 0 394588 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4283
timestamp 1676037725
transform 1 0 395140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4285
timestamp 1676037725
transform 1 0 395324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4297
timestamp 1676037725
transform 1 0 396428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4309
timestamp 1676037725
transform 1 0 397532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4321
timestamp 1676037725
transform 1 0 398636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4333
timestamp 1676037725
transform 1 0 399740 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4339
timestamp 1676037725
transform 1 0 400292 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4341
timestamp 1676037725
transform 1 0 400476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4353
timestamp 1676037725
transform 1 0 401580 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4365
timestamp 1676037725
transform 1 0 402684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4377
timestamp 1676037725
transform 1 0 403788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4389
timestamp 1676037725
transform 1 0 404892 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4395
timestamp 1676037725
transform 1 0 405444 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4397
timestamp 1676037725
transform 1 0 405628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4409
timestamp 1676037725
transform 1 0 406732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4421
timestamp 1676037725
transform 1 0 407836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4433
timestamp 1676037725
transform 1 0 408940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4445
timestamp 1676037725
transform 1 0 410044 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4451
timestamp 1676037725
transform 1 0 410596 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4453
timestamp 1676037725
transform 1 0 410780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4465
timestamp 1676037725
transform 1 0 411884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4477
timestamp 1676037725
transform 1 0 412988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4489
timestamp 1676037725
transform 1 0 414092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4501
timestamp 1676037725
transform 1 0 415196 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4507
timestamp 1676037725
transform 1 0 415748 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4509
timestamp 1676037725
transform 1 0 415932 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4521
timestamp 1676037725
transform 1 0 417036 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4533
timestamp 1676037725
transform 1 0 418140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4545
timestamp 1676037725
transform 1 0 419244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4557
timestamp 1676037725
transform 1 0 420348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4563
timestamp 1676037725
transform 1 0 420900 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4565
timestamp 1676037725
transform 1 0 421084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4577
timestamp 1676037725
transform 1 0 422188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4589
timestamp 1676037725
transform 1 0 423292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4601
timestamp 1676037725
transform 1 0 424396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4613
timestamp 1676037725
transform 1 0 425500 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4619
timestamp 1676037725
transform 1 0 426052 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4621
timestamp 1676037725
transform 1 0 426236 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4633
timestamp 1676037725
transform 1 0 427340 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4645
timestamp 1676037725
transform 1 0 428444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4657
timestamp 1676037725
transform 1 0 429548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4669
timestamp 1676037725
transform 1 0 430652 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4675
timestamp 1676037725
transform 1 0 431204 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4677
timestamp 1676037725
transform 1 0 431388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4689
timestamp 1676037725
transform 1 0 432492 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4701
timestamp 1676037725
transform 1 0 433596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4713
timestamp 1676037725
transform 1 0 434700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4725
timestamp 1676037725
transform 1 0 435804 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4731
timestamp 1676037725
transform 1 0 436356 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4733
timestamp 1676037725
transform 1 0 436540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4745
timestamp 1676037725
transform 1 0 437644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4757
timestamp 1676037725
transform 1 0 438748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4769
timestamp 1676037725
transform 1 0 439852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4781
timestamp 1676037725
transform 1 0 440956 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4787
timestamp 1676037725
transform 1 0 441508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4789
timestamp 1676037725
transform 1 0 441692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4801
timestamp 1676037725
transform 1 0 442796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4813
timestamp 1676037725
transform 1 0 443900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4825
timestamp 1676037725
transform 1 0 445004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4837
timestamp 1676037725
transform 1 0 446108 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4843
timestamp 1676037725
transform 1 0 446660 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4845
timestamp 1676037725
transform 1 0 446844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4857
timestamp 1676037725
transform 1 0 447948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4869
timestamp 1676037725
transform 1 0 449052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4881
timestamp 1676037725
transform 1 0 450156 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4893
timestamp 1676037725
transform 1 0 451260 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4899
timestamp 1676037725
transform 1 0 451812 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4901
timestamp 1676037725
transform 1 0 451996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4913
timestamp 1676037725
transform 1 0 453100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4925
timestamp 1676037725
transform 1 0 454204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4937
timestamp 1676037725
transform 1 0 455308 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_4949
timestamp 1676037725
transform 1 0 456412 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_4955
timestamp 1676037725
transform 1 0 456964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4957
timestamp 1676037725
transform 1 0 457148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4969
timestamp 1676037725
transform 1 0 458252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4981
timestamp 1676037725
transform 1 0 459356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_4993
timestamp 1676037725
transform 1 0 460460 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5005
timestamp 1676037725
transform 1 0 461564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5011
timestamp 1676037725
transform 1 0 462116 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5013
timestamp 1676037725
transform 1 0 462300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5025
timestamp 1676037725
transform 1 0 463404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5037
timestamp 1676037725
transform 1 0 464508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5049
timestamp 1676037725
transform 1 0 465612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5061
timestamp 1676037725
transform 1 0 466716 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5067
timestamp 1676037725
transform 1 0 467268 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5069
timestamp 1676037725
transform 1 0 467452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5081
timestamp 1676037725
transform 1 0 468556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5093
timestamp 1676037725
transform 1 0 469660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5105
timestamp 1676037725
transform 1 0 470764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5117
timestamp 1676037725
transform 1 0 471868 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5123
timestamp 1676037725
transform 1 0 472420 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5125
timestamp 1676037725
transform 1 0 472604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5137
timestamp 1676037725
transform 1 0 473708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5149
timestamp 1676037725
transform 1 0 474812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5161
timestamp 1676037725
transform 1 0 475916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5173
timestamp 1676037725
transform 1 0 477020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5179
timestamp 1676037725
transform 1 0 477572 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5181
timestamp 1676037725
transform 1 0 477756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5193
timestamp 1676037725
transform 1 0 478860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5205
timestamp 1676037725
transform 1 0 479964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5217
timestamp 1676037725
transform 1 0 481068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5229
timestamp 1676037725
transform 1 0 482172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5235
timestamp 1676037725
transform 1 0 482724 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5237
timestamp 1676037725
transform 1 0 482908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5249
timestamp 1676037725
transform 1 0 484012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5261
timestamp 1676037725
transform 1 0 485116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5273
timestamp 1676037725
transform 1 0 486220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5285
timestamp 1676037725
transform 1 0 487324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5291
timestamp 1676037725
transform 1 0 487876 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5293
timestamp 1676037725
transform 1 0 488060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5305
timestamp 1676037725
transform 1 0 489164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5317
timestamp 1676037725
transform 1 0 490268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5329
timestamp 1676037725
transform 1 0 491372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5341
timestamp 1676037725
transform 1 0 492476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5347
timestamp 1676037725
transform 1 0 493028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5349
timestamp 1676037725
transform 1 0 493212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5361
timestamp 1676037725
transform 1 0 494316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5373
timestamp 1676037725
transform 1 0 495420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5385
timestamp 1676037725
transform 1 0 496524 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5397
timestamp 1676037725
transform 1 0 497628 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5403
timestamp 1676037725
transform 1 0 498180 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5405
timestamp 1676037725
transform 1 0 498364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5417
timestamp 1676037725
transform 1 0 499468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5429
timestamp 1676037725
transform 1 0 500572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5441
timestamp 1676037725
transform 1 0 501676 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5453
timestamp 1676037725
transform 1 0 502780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5459
timestamp 1676037725
transform 1 0 503332 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5461
timestamp 1676037725
transform 1 0 503516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5473
timestamp 1676037725
transform 1 0 504620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5485
timestamp 1676037725
transform 1 0 505724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5497
timestamp 1676037725
transform 1 0 506828 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5509
timestamp 1676037725
transform 1 0 507932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5515
timestamp 1676037725
transform 1 0 508484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5517
timestamp 1676037725
transform 1 0 508668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5529
timestamp 1676037725
transform 1 0 509772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5541
timestamp 1676037725
transform 1 0 510876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5553
timestamp 1676037725
transform 1 0 511980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5565
timestamp 1676037725
transform 1 0 513084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5571
timestamp 1676037725
transform 1 0 513636 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5573
timestamp 1676037725
transform 1 0 513820 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5585
timestamp 1676037725
transform 1 0 514924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5597
timestamp 1676037725
transform 1 0 516028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5609
timestamp 1676037725
transform 1 0 517132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5621
timestamp 1676037725
transform 1 0 518236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5627
timestamp 1676037725
transform 1 0 518788 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5629
timestamp 1676037725
transform 1 0 518972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5641
timestamp 1676037725
transform 1 0 520076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5653
timestamp 1676037725
transform 1 0 521180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5665
timestamp 1676037725
transform 1 0 522284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_5677
timestamp 1676037725
transform 1 0 523388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_5683
timestamp 1676037725
transform 1 0 523940 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5685
timestamp 1676037725
transform 1 0 524124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5697
timestamp 1676037725
transform 1 0 525228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5709
timestamp 1676037725
transform 1 0 526332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5721
timestamp 1676037725
transform 1 0 527436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1676037725
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1676037725
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1676037725
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1676037725
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1676037725
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1676037725
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1676037725
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1676037725
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1676037725
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1676037725
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1676037725
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1676037725
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1676037725
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1676037725
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1676037725
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1676037725
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1676037725
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1676037725
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1676037725
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1676037725
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1676037725
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1676037725
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1676037725
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1676037725
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1676037725
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1676037725
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_821
timestamp 1676037725
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1676037725
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1676037725
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1676037725
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1676037725
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_865
timestamp 1676037725
transform 1 0 80684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_877
timestamp 1676037725
transform 1 0 81788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_889
timestamp 1676037725
transform 1 0 82892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_895
timestamp 1676037725
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1676037725
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1676037725
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_921
timestamp 1676037725
transform 1 0 85836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_933
timestamp 1676037725
transform 1 0 86940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_945
timestamp 1676037725
transform 1 0 88044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_951
timestamp 1676037725
transform 1 0 88596 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1676037725
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_965
timestamp 1676037725
transform 1 0 89884 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_971
timestamp 1676037725
transform 1 0 90436 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_974
timestamp 1676037725
transform 1 0 90712 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_987
timestamp 1676037725
transform 1 0 91908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_993
timestamp 1676037725
transform 1 0 92460 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1006
timestamp 1676037725
transform 1 0 93656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1009
timestamp 1676037725
transform 1 0 93932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1021
timestamp 1676037725
transform 1 0 95036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1034
timestamp 1676037725
transform 1 0 96232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1047
timestamp 1676037725
transform 1 0 97428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1060
timestamp 1676037725
transform 1 0 98624 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1065
timestamp 1676037725
transform 1 0 99084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1071
timestamp 1676037725
transform 1 0 99636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1084
timestamp 1676037725
transform 1 0 100832 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1097
timestamp 1676037725
transform 1 0 102028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1109
timestamp 1676037725
transform 1 0 103132 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1112
timestamp 1676037725
transform 1 0 103408 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1676037725
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1676037725
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1145
timestamp 1676037725
transform 1 0 106444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1157
timestamp 1676037725
transform 1 0 107548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1169
timestamp 1676037725
transform 1 0 108652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1175
timestamp 1676037725
transform 1 0 109204 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1676037725
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1189
timestamp 1676037725
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1201
timestamp 1676037725
transform 1 0 111596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1213
timestamp 1676037725
transform 1 0 112700 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1219
timestamp 1676037725
transform 1 0 113252 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1222
timestamp 1676037725
transform 1 0 113528 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1230
timestamp 1676037725
transform 1 0 114264 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1676037725
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1676037725
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1257
timestamp 1676037725
transform 1 0 116748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1269
timestamp 1676037725
transform 1 0 117852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1281
timestamp 1676037725
transform 1 0 118956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1287
timestamp 1676037725
transform 1 0 119508 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1289
timestamp 1676037725
transform 1 0 119692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1301
timestamp 1676037725
transform 1 0 120796 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1313
timestamp 1676037725
transform 1 0 121900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1325
timestamp 1676037725
transform 1 0 123004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1337
timestamp 1676037725
transform 1 0 124108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1343
timestamp 1676037725
transform 1 0 124660 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1345
timestamp 1676037725
transform 1 0 124844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1357
timestamp 1676037725
transform 1 0 125948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1369
timestamp 1676037725
transform 1 0 127052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1381
timestamp 1676037725
transform 1 0 128156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1393
timestamp 1676037725
transform 1 0 129260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1399
timestamp 1676037725
transform 1 0 129812 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1401
timestamp 1676037725
transform 1 0 129996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1413
timestamp 1676037725
transform 1 0 131100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1425
timestamp 1676037725
transform 1 0 132204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1437
timestamp 1676037725
transform 1 0 133308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1449
timestamp 1676037725
transform 1 0 134412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1455
timestamp 1676037725
transform 1 0 134964 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1457
timestamp 1676037725
transform 1 0 135148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1469
timestamp 1676037725
transform 1 0 136252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1481
timestamp 1676037725
transform 1 0 137356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1493
timestamp 1676037725
transform 1 0 138460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1505
timestamp 1676037725
transform 1 0 139564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1511
timestamp 1676037725
transform 1 0 140116 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1513
timestamp 1676037725
transform 1 0 140300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1525
timestamp 1676037725
transform 1 0 141404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1537
timestamp 1676037725
transform 1 0 142508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1549
timestamp 1676037725
transform 1 0 143612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1561
timestamp 1676037725
transform 1 0 144716 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1567
timestamp 1676037725
transform 1 0 145268 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1569
timestamp 1676037725
transform 1 0 145452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1581
timestamp 1676037725
transform 1 0 146556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1593
timestamp 1676037725
transform 1 0 147660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1605
timestamp 1676037725
transform 1 0 148764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1617
timestamp 1676037725
transform 1 0 149868 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1623
timestamp 1676037725
transform 1 0 150420 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1625
timestamp 1676037725
transform 1 0 150604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1637
timestamp 1676037725
transform 1 0 151708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1649
timestamp 1676037725
transform 1 0 152812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1661
timestamp 1676037725
transform 1 0 153916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1673
timestamp 1676037725
transform 1 0 155020 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1679
timestamp 1676037725
transform 1 0 155572 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1681
timestamp 1676037725
transform 1 0 155756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1693
timestamp 1676037725
transform 1 0 156860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1705
timestamp 1676037725
transform 1 0 157964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1717
timestamp 1676037725
transform 1 0 159068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1729
timestamp 1676037725
transform 1 0 160172 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1735
timestamp 1676037725
transform 1 0 160724 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1737
timestamp 1676037725
transform 1 0 160908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1749
timestamp 1676037725
transform 1 0 162012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1761
timestamp 1676037725
transform 1 0 163116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1773
timestamp 1676037725
transform 1 0 164220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1785
timestamp 1676037725
transform 1 0 165324 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1791
timestamp 1676037725
transform 1 0 165876 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1793
timestamp 1676037725
transform 1 0 166060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1805
timestamp 1676037725
transform 1 0 167164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1817
timestamp 1676037725
transform 1 0 168268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1829
timestamp 1676037725
transform 1 0 169372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1841
timestamp 1676037725
transform 1 0 170476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1847
timestamp 1676037725
transform 1 0 171028 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1849
timestamp 1676037725
transform 1 0 171212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1861
timestamp 1676037725
transform 1 0 172316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1873
timestamp 1676037725
transform 1 0 173420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1885
timestamp 1676037725
transform 1 0 174524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1897
timestamp 1676037725
transform 1 0 175628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1903
timestamp 1676037725
transform 1 0 176180 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1905
timestamp 1676037725
transform 1 0 176364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1917
timestamp 1676037725
transform 1 0 177468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1929
timestamp 1676037725
transform 1 0 178572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1941
timestamp 1676037725
transform 1 0 179676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1953
timestamp 1676037725
transform 1 0 180780 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1959
timestamp 1676037725
transform 1 0 181332 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1961
timestamp 1676037725
transform 1 0 181516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1973
timestamp 1676037725
transform 1 0 182620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1985
timestamp 1676037725
transform 1 0 183724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1997
timestamp 1676037725
transform 1 0 184828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2009
timestamp 1676037725
transform 1 0 185932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2015
timestamp 1676037725
transform 1 0 186484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2017
timestamp 1676037725
transform 1 0 186668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2029
timestamp 1676037725
transform 1 0 187772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2041
timestamp 1676037725
transform 1 0 188876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2053
timestamp 1676037725
transform 1 0 189980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2065
timestamp 1676037725
transform 1 0 191084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2071
timestamp 1676037725
transform 1 0 191636 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2073
timestamp 1676037725
transform 1 0 191820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2085
timestamp 1676037725
transform 1 0 192924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2097
timestamp 1676037725
transform 1 0 194028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2109
timestamp 1676037725
transform 1 0 195132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2121
timestamp 1676037725
transform 1 0 196236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2127
timestamp 1676037725
transform 1 0 196788 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2129
timestamp 1676037725
transform 1 0 196972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2141
timestamp 1676037725
transform 1 0 198076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2153
timestamp 1676037725
transform 1 0 199180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2165
timestamp 1676037725
transform 1 0 200284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2177
timestamp 1676037725
transform 1 0 201388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2183
timestamp 1676037725
transform 1 0 201940 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2185
timestamp 1676037725
transform 1 0 202124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2197
timestamp 1676037725
transform 1 0 203228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2209
timestamp 1676037725
transform 1 0 204332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2221
timestamp 1676037725
transform 1 0 205436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2233
timestamp 1676037725
transform 1 0 206540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2239
timestamp 1676037725
transform 1 0 207092 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2241
timestamp 1676037725
transform 1 0 207276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2253
timestamp 1676037725
transform 1 0 208380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2265
timestamp 1676037725
transform 1 0 209484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2277
timestamp 1676037725
transform 1 0 210588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2289
timestamp 1676037725
transform 1 0 211692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2295
timestamp 1676037725
transform 1 0 212244 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2297
timestamp 1676037725
transform 1 0 212428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2309
timestamp 1676037725
transform 1 0 213532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2321
timestamp 1676037725
transform 1 0 214636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2333
timestamp 1676037725
transform 1 0 215740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2345
timestamp 1676037725
transform 1 0 216844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2351
timestamp 1676037725
transform 1 0 217396 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2353
timestamp 1676037725
transform 1 0 217580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2365
timestamp 1676037725
transform 1 0 218684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2377
timestamp 1676037725
transform 1 0 219788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2389
timestamp 1676037725
transform 1 0 220892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2401
timestamp 1676037725
transform 1 0 221996 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2407
timestamp 1676037725
transform 1 0 222548 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2409
timestamp 1676037725
transform 1 0 222732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2421
timestamp 1676037725
transform 1 0 223836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2433
timestamp 1676037725
transform 1 0 224940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2445
timestamp 1676037725
transform 1 0 226044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2457
timestamp 1676037725
transform 1 0 227148 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2463
timestamp 1676037725
transform 1 0 227700 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2465
timestamp 1676037725
transform 1 0 227884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2477
timestamp 1676037725
transform 1 0 228988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2489
timestamp 1676037725
transform 1 0 230092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2501
timestamp 1676037725
transform 1 0 231196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2513
timestamp 1676037725
transform 1 0 232300 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2519
timestamp 1676037725
transform 1 0 232852 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2521
timestamp 1676037725
transform 1 0 233036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2533
timestamp 1676037725
transform 1 0 234140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2545
timestamp 1676037725
transform 1 0 235244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2557
timestamp 1676037725
transform 1 0 236348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2569
timestamp 1676037725
transform 1 0 237452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2575
timestamp 1676037725
transform 1 0 238004 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2577
timestamp 1676037725
transform 1 0 238188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2589
timestamp 1676037725
transform 1 0 239292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2601
timestamp 1676037725
transform 1 0 240396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2613
timestamp 1676037725
transform 1 0 241500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2625
timestamp 1676037725
transform 1 0 242604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2631
timestamp 1676037725
transform 1 0 243156 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2633
timestamp 1676037725
transform 1 0 243340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2645
timestamp 1676037725
transform 1 0 244444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2657
timestamp 1676037725
transform 1 0 245548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2669
timestamp 1676037725
transform 1 0 246652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2681
timestamp 1676037725
transform 1 0 247756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2687
timestamp 1676037725
transform 1 0 248308 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2689
timestamp 1676037725
transform 1 0 248492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2703
timestamp 1676037725
transform 1 0 249780 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2716
timestamp 1676037725
transform 1 0 250976 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2729
timestamp 1676037725
transform 1 0 252172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_2742
timestamp 1676037725
transform 1 0 253368 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2745
timestamp 1676037725
transform 1 0 253644 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2749
timestamp 1676037725
transform 1 0 254012 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2759
timestamp 1676037725
transform 1 0 254932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2776
timestamp 1676037725
transform 1 0 256496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2782
timestamp 1676037725
transform 1 0 257048 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2794
timestamp 1676037725
transform 1 0 258152 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2801
timestamp 1676037725
transform 1 0 258796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2813
timestamp 1676037725
transform 1 0 259900 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2821
timestamp 1676037725
transform 1 0 260636 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2831
timestamp 1676037725
transform 1 0 261556 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2837
timestamp 1676037725
transform 1 0 262108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2849
timestamp 1676037725
transform 1 0 263212 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2855
timestamp 1676037725
transform 1 0 263764 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2857
timestamp 1676037725
transform 1 0 263948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2869
timestamp 1676037725
transform 1 0 265052 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2886
timestamp 1676037725
transform 1 0 266616 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2892
timestamp 1676037725
transform 1 0 267168 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2904
timestamp 1676037725
transform 1 0 268272 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2913
timestamp 1676037725
transform 1 0 269100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_2925
timestamp 1676037725
transform 1 0 270204 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2931
timestamp 1676037725
transform 1 0 270756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_2941
timestamp 1676037725
transform 1 0 271676 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2947
timestamp 1676037725
transform 1 0 272228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_2959
timestamp 1676037725
transform 1 0 273332 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_2967
timestamp 1676037725
transform 1 0 274068 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2969
timestamp 1676037725
transform 1 0 274252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2981
timestamp 1676037725
transform 1 0 275356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_2993
timestamp 1676037725
transform 1 0 276460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3005
timestamp 1676037725
transform 1 0 277564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3017
timestamp 1676037725
transform 1 0 278668 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3023
timestamp 1676037725
transform 1 0 279220 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3025
timestamp 1676037725
transform 1 0 279404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3037
timestamp 1676037725
transform 1 0 280508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3049
timestamp 1676037725
transform 1 0 281612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3061
timestamp 1676037725
transform 1 0 282716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3073
timestamp 1676037725
transform 1 0 283820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3079
timestamp 1676037725
transform 1 0 284372 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3081
timestamp 1676037725
transform 1 0 284556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3093
timestamp 1676037725
transform 1 0 285660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3105
timestamp 1676037725
transform 1 0 286764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3117
timestamp 1676037725
transform 1 0 287868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3129
timestamp 1676037725
transform 1 0 288972 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3135
timestamp 1676037725
transform 1 0 289524 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3137
timestamp 1676037725
transform 1 0 289708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3149
timestamp 1676037725
transform 1 0 290812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3161
timestamp 1676037725
transform 1 0 291916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3173
timestamp 1676037725
transform 1 0 293020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3185
timestamp 1676037725
transform 1 0 294124 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3191
timestamp 1676037725
transform 1 0 294676 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3193
timestamp 1676037725
transform 1 0 294860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3205
timestamp 1676037725
transform 1 0 295964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3217
timestamp 1676037725
transform 1 0 297068 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3229
timestamp 1676037725
transform 1 0 298172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3241
timestamp 1676037725
transform 1 0 299276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3247
timestamp 1676037725
transform 1 0 299828 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3249
timestamp 1676037725
transform 1 0 300012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3261
timestamp 1676037725
transform 1 0 301116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3273
timestamp 1676037725
transform 1 0 302220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3285
timestamp 1676037725
transform 1 0 303324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3297
timestamp 1676037725
transform 1 0 304428 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3303
timestamp 1676037725
transform 1 0 304980 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3305
timestamp 1676037725
transform 1 0 305164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3317
timestamp 1676037725
transform 1 0 306268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3329
timestamp 1676037725
transform 1 0 307372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3341
timestamp 1676037725
transform 1 0 308476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3353
timestamp 1676037725
transform 1 0 309580 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3359
timestamp 1676037725
transform 1 0 310132 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3361
timestamp 1676037725
transform 1 0 310316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3373
timestamp 1676037725
transform 1 0 311420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3385
timestamp 1676037725
transform 1 0 312524 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3397
timestamp 1676037725
transform 1 0 313628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3409
timestamp 1676037725
transform 1 0 314732 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3415
timestamp 1676037725
transform 1 0 315284 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3417
timestamp 1676037725
transform 1 0 315468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3429
timestamp 1676037725
transform 1 0 316572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3441
timestamp 1676037725
transform 1 0 317676 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3453
timestamp 1676037725
transform 1 0 318780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3465
timestamp 1676037725
transform 1 0 319884 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3471
timestamp 1676037725
transform 1 0 320436 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3473
timestamp 1676037725
transform 1 0 320620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3485
timestamp 1676037725
transform 1 0 321724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3497
timestamp 1676037725
transform 1 0 322828 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3509
timestamp 1676037725
transform 1 0 323932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3521
timestamp 1676037725
transform 1 0 325036 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3527
timestamp 1676037725
transform 1 0 325588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3529
timestamp 1676037725
transform 1 0 325772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3541
timestamp 1676037725
transform 1 0 326876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3553
timestamp 1676037725
transform 1 0 327980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3565
timestamp 1676037725
transform 1 0 329084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3577
timestamp 1676037725
transform 1 0 330188 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3583
timestamp 1676037725
transform 1 0 330740 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3585
timestamp 1676037725
transform 1 0 330924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3597
timestamp 1676037725
transform 1 0 332028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3609
timestamp 1676037725
transform 1 0 333132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3621
timestamp 1676037725
transform 1 0 334236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3633
timestamp 1676037725
transform 1 0 335340 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3639
timestamp 1676037725
transform 1 0 335892 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3641
timestamp 1676037725
transform 1 0 336076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3653
timestamp 1676037725
transform 1 0 337180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3665
timestamp 1676037725
transform 1 0 338284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3677
timestamp 1676037725
transform 1 0 339388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3689
timestamp 1676037725
transform 1 0 340492 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3695
timestamp 1676037725
transform 1 0 341044 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3697
timestamp 1676037725
transform 1 0 341228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3709
timestamp 1676037725
transform 1 0 342332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3721
timestamp 1676037725
transform 1 0 343436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3733
timestamp 1676037725
transform 1 0 344540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3745
timestamp 1676037725
transform 1 0 345644 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3751
timestamp 1676037725
transform 1 0 346196 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3753
timestamp 1676037725
transform 1 0 346380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3765
timestamp 1676037725
transform 1 0 347484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3777
timestamp 1676037725
transform 1 0 348588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3789
timestamp 1676037725
transform 1 0 349692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3801
timestamp 1676037725
transform 1 0 350796 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3807
timestamp 1676037725
transform 1 0 351348 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3809
timestamp 1676037725
transform 1 0 351532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3821
timestamp 1676037725
transform 1 0 352636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3833
timestamp 1676037725
transform 1 0 353740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3845
timestamp 1676037725
transform 1 0 354844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3857
timestamp 1676037725
transform 1 0 355948 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3863
timestamp 1676037725
transform 1 0 356500 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3865
timestamp 1676037725
transform 1 0 356684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3877
timestamp 1676037725
transform 1 0 357788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3889
timestamp 1676037725
transform 1 0 358892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3901
timestamp 1676037725
transform 1 0 359996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3913
timestamp 1676037725
transform 1 0 361100 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3919
timestamp 1676037725
transform 1 0 361652 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3921
timestamp 1676037725
transform 1 0 361836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3933
timestamp 1676037725
transform 1 0 362940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3945
timestamp 1676037725
transform 1 0 364044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3957
timestamp 1676037725
transform 1 0 365148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3969
timestamp 1676037725
transform 1 0 366252 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3975
timestamp 1676037725
transform 1 0 366804 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3977
timestamp 1676037725
transform 1 0 366988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3989
timestamp 1676037725
transform 1 0 368092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4001
timestamp 1676037725
transform 1 0 369196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4013
timestamp 1676037725
transform 1 0 370300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4025
timestamp 1676037725
transform 1 0 371404 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4031
timestamp 1676037725
transform 1 0 371956 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4033
timestamp 1676037725
transform 1 0 372140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4045
timestamp 1676037725
transform 1 0 373244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4057
timestamp 1676037725
transform 1 0 374348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4069
timestamp 1676037725
transform 1 0 375452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4081
timestamp 1676037725
transform 1 0 376556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4087
timestamp 1676037725
transform 1 0 377108 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4089
timestamp 1676037725
transform 1 0 377292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4101
timestamp 1676037725
transform 1 0 378396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4113
timestamp 1676037725
transform 1 0 379500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4125
timestamp 1676037725
transform 1 0 380604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4137
timestamp 1676037725
transform 1 0 381708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4143
timestamp 1676037725
transform 1 0 382260 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4145
timestamp 1676037725
transform 1 0 382444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4157
timestamp 1676037725
transform 1 0 383548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4169
timestamp 1676037725
transform 1 0 384652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4181
timestamp 1676037725
transform 1 0 385756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4193
timestamp 1676037725
transform 1 0 386860 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4199
timestamp 1676037725
transform 1 0 387412 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4201
timestamp 1676037725
transform 1 0 387596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4213
timestamp 1676037725
transform 1 0 388700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4225
timestamp 1676037725
transform 1 0 389804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4237
timestamp 1676037725
transform 1 0 390908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4249
timestamp 1676037725
transform 1 0 392012 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4255
timestamp 1676037725
transform 1 0 392564 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4257
timestamp 1676037725
transform 1 0 392748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4269
timestamp 1676037725
transform 1 0 393852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4281
timestamp 1676037725
transform 1 0 394956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4293
timestamp 1676037725
transform 1 0 396060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4305
timestamp 1676037725
transform 1 0 397164 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4311
timestamp 1676037725
transform 1 0 397716 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4313
timestamp 1676037725
transform 1 0 397900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4325
timestamp 1676037725
transform 1 0 399004 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4337
timestamp 1676037725
transform 1 0 400108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4349
timestamp 1676037725
transform 1 0 401212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4361
timestamp 1676037725
transform 1 0 402316 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4367
timestamp 1676037725
transform 1 0 402868 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4369
timestamp 1676037725
transform 1 0 403052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4381
timestamp 1676037725
transform 1 0 404156 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4393
timestamp 1676037725
transform 1 0 405260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4405
timestamp 1676037725
transform 1 0 406364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4417
timestamp 1676037725
transform 1 0 407468 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4423
timestamp 1676037725
transform 1 0 408020 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4425
timestamp 1676037725
transform 1 0 408204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4437
timestamp 1676037725
transform 1 0 409308 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4449
timestamp 1676037725
transform 1 0 410412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4461
timestamp 1676037725
transform 1 0 411516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4473
timestamp 1676037725
transform 1 0 412620 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4479
timestamp 1676037725
transform 1 0 413172 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4481
timestamp 1676037725
transform 1 0 413356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4493
timestamp 1676037725
transform 1 0 414460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4505
timestamp 1676037725
transform 1 0 415564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4517
timestamp 1676037725
transform 1 0 416668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4529
timestamp 1676037725
transform 1 0 417772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4535
timestamp 1676037725
transform 1 0 418324 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4537
timestamp 1676037725
transform 1 0 418508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4549
timestamp 1676037725
transform 1 0 419612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4561
timestamp 1676037725
transform 1 0 420716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4573
timestamp 1676037725
transform 1 0 421820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4585
timestamp 1676037725
transform 1 0 422924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4591
timestamp 1676037725
transform 1 0 423476 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4593
timestamp 1676037725
transform 1 0 423660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4605
timestamp 1676037725
transform 1 0 424764 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4617
timestamp 1676037725
transform 1 0 425868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4629
timestamp 1676037725
transform 1 0 426972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4641
timestamp 1676037725
transform 1 0 428076 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4647
timestamp 1676037725
transform 1 0 428628 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4649
timestamp 1676037725
transform 1 0 428812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4661
timestamp 1676037725
transform 1 0 429916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4673
timestamp 1676037725
transform 1 0 431020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4685
timestamp 1676037725
transform 1 0 432124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4697
timestamp 1676037725
transform 1 0 433228 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4703
timestamp 1676037725
transform 1 0 433780 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4705
timestamp 1676037725
transform 1 0 433964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4717
timestamp 1676037725
transform 1 0 435068 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4729
timestamp 1676037725
transform 1 0 436172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4741
timestamp 1676037725
transform 1 0 437276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4753
timestamp 1676037725
transform 1 0 438380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4759
timestamp 1676037725
transform 1 0 438932 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4761
timestamp 1676037725
transform 1 0 439116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4773
timestamp 1676037725
transform 1 0 440220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4785
timestamp 1676037725
transform 1 0 441324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4797
timestamp 1676037725
transform 1 0 442428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4809
timestamp 1676037725
transform 1 0 443532 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4815
timestamp 1676037725
transform 1 0 444084 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4817
timestamp 1676037725
transform 1 0 444268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4829
timestamp 1676037725
transform 1 0 445372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4841
timestamp 1676037725
transform 1 0 446476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4853
timestamp 1676037725
transform 1 0 447580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4865
timestamp 1676037725
transform 1 0 448684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4871
timestamp 1676037725
transform 1 0 449236 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4873
timestamp 1676037725
transform 1 0 449420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4885
timestamp 1676037725
transform 1 0 450524 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4897
timestamp 1676037725
transform 1 0 451628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4909
timestamp 1676037725
transform 1 0 452732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4921
timestamp 1676037725
transform 1 0 453836 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4927
timestamp 1676037725
transform 1 0 454388 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4929
timestamp 1676037725
transform 1 0 454572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4941
timestamp 1676037725
transform 1 0 455676 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4953
timestamp 1676037725
transform 1 0 456780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4965
timestamp 1676037725
transform 1 0 457884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_4977
timestamp 1676037725
transform 1 0 458988 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_4983
timestamp 1676037725
transform 1 0 459540 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4985
timestamp 1676037725
transform 1 0 459724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_4997
timestamp 1676037725
transform 1 0 460828 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5009
timestamp 1676037725
transform 1 0 461932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5021
timestamp 1676037725
transform 1 0 463036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5033
timestamp 1676037725
transform 1 0 464140 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5039
timestamp 1676037725
transform 1 0 464692 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5041
timestamp 1676037725
transform 1 0 464876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5053
timestamp 1676037725
transform 1 0 465980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5065
timestamp 1676037725
transform 1 0 467084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5077
timestamp 1676037725
transform 1 0 468188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5089
timestamp 1676037725
transform 1 0 469292 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5095
timestamp 1676037725
transform 1 0 469844 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5097
timestamp 1676037725
transform 1 0 470028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5109
timestamp 1676037725
transform 1 0 471132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5121
timestamp 1676037725
transform 1 0 472236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5133
timestamp 1676037725
transform 1 0 473340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5145
timestamp 1676037725
transform 1 0 474444 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5151
timestamp 1676037725
transform 1 0 474996 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5153
timestamp 1676037725
transform 1 0 475180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5165
timestamp 1676037725
transform 1 0 476284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5177
timestamp 1676037725
transform 1 0 477388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5189
timestamp 1676037725
transform 1 0 478492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5201
timestamp 1676037725
transform 1 0 479596 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5207
timestamp 1676037725
transform 1 0 480148 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5209
timestamp 1676037725
transform 1 0 480332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5221
timestamp 1676037725
transform 1 0 481436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5233
timestamp 1676037725
transform 1 0 482540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5245
timestamp 1676037725
transform 1 0 483644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5257
timestamp 1676037725
transform 1 0 484748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5263
timestamp 1676037725
transform 1 0 485300 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5265
timestamp 1676037725
transform 1 0 485484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5277
timestamp 1676037725
transform 1 0 486588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5289
timestamp 1676037725
transform 1 0 487692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5301
timestamp 1676037725
transform 1 0 488796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5313
timestamp 1676037725
transform 1 0 489900 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5319
timestamp 1676037725
transform 1 0 490452 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5321
timestamp 1676037725
transform 1 0 490636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5333
timestamp 1676037725
transform 1 0 491740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5345
timestamp 1676037725
transform 1 0 492844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5357
timestamp 1676037725
transform 1 0 493948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5369
timestamp 1676037725
transform 1 0 495052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5375
timestamp 1676037725
transform 1 0 495604 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5377
timestamp 1676037725
transform 1 0 495788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5389
timestamp 1676037725
transform 1 0 496892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5401
timestamp 1676037725
transform 1 0 497996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5413
timestamp 1676037725
transform 1 0 499100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5425
timestamp 1676037725
transform 1 0 500204 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5431
timestamp 1676037725
transform 1 0 500756 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5433
timestamp 1676037725
transform 1 0 500940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5445
timestamp 1676037725
transform 1 0 502044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5457
timestamp 1676037725
transform 1 0 503148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5469
timestamp 1676037725
transform 1 0 504252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5481
timestamp 1676037725
transform 1 0 505356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5487
timestamp 1676037725
transform 1 0 505908 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5489
timestamp 1676037725
transform 1 0 506092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5501
timestamp 1676037725
transform 1 0 507196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5513
timestamp 1676037725
transform 1 0 508300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5525
timestamp 1676037725
transform 1 0 509404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5537
timestamp 1676037725
transform 1 0 510508 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5543
timestamp 1676037725
transform 1 0 511060 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5545
timestamp 1676037725
transform 1 0 511244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5557
timestamp 1676037725
transform 1 0 512348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5569
timestamp 1676037725
transform 1 0 513452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5581
timestamp 1676037725
transform 1 0 514556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5593
timestamp 1676037725
transform 1 0 515660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5599
timestamp 1676037725
transform 1 0 516212 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5601
timestamp 1676037725
transform 1 0 516396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5613
timestamp 1676037725
transform 1 0 517500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5625
timestamp 1676037725
transform 1 0 518604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5637
timestamp 1676037725
transform 1 0 519708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5649
timestamp 1676037725
transform 1 0 520812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5655
timestamp 1676037725
transform 1 0 521364 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5657
timestamp 1676037725
transform 1 0 521548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5669
timestamp 1676037725
transform 1 0 522652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5681
timestamp 1676037725
transform 1 0 523756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5693
timestamp 1676037725
transform 1 0 524860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_5705
timestamp 1676037725
transform 1 0 525964 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_5711
timestamp 1676037725
transform 1 0 526516 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5713
timestamp 1676037725
transform 1 0 526700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_5725
timestamp 1676037725
transform 1 0 527804 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1676037725
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1676037725
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1676037725
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1676037725
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1676037725
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1676037725
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1676037725
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1676037725
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1676037725
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1676037725
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1676037725
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1676037725
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1676037725
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1676037725
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1676037725
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1676037725
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1676037725
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1676037725
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1676037725
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1676037725
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1676037725
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1676037725
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1676037725
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1676037725
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1676037725
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1676037725
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1676037725
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1676037725
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1676037725
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1676037725
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1676037725
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_813
timestamp 1676037725
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_825
timestamp 1676037725
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_837
timestamp 1676037725
transform 1 0 78108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_849
timestamp 1676037725
transform 1 0 79212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_861
timestamp 1676037725
transform 1 0 80316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_867
timestamp 1676037725
transform 1 0 80868 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_869
timestamp 1676037725
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_881
timestamp 1676037725
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_893
timestamp 1676037725
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_905
timestamp 1676037725
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_917
timestamp 1676037725
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_923
timestamp 1676037725
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_925
timestamp 1676037725
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_937
timestamp 1676037725
transform 1 0 87308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_949
timestamp 1676037725
transform 1 0 88412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_961
timestamp 1676037725
transform 1 0 89516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_973
timestamp 1676037725
transform 1 0 90620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_979
timestamp 1676037725
transform 1 0 91172 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_981
timestamp 1676037725
transform 1 0 91356 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_986
timestamp 1676037725
transform 1 0 91816 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_999
timestamp 1676037725
transform 1 0 93012 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1007
timestamp 1676037725
transform 1 0 93748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1012
timestamp 1676037725
transform 1 0 94208 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1020
timestamp 1676037725
transform 1 0 94944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1025
timestamp 1676037725
transform 1 0 95404 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1033
timestamp 1676037725
transform 1 0 96140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1037
timestamp 1676037725
transform 1 0 96508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1041
timestamp 1676037725
transform 1 0 96876 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1051
timestamp 1676037725
transform 1 0 97796 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1063
timestamp 1676037725
transform 1 0 98900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1075
timestamp 1676037725
transform 1 0 100004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1083
timestamp 1676037725
transform 1 0 100740 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1088
timestamp 1676037725
transform 1 0 101200 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1093
timestamp 1676037725
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1105
timestamp 1676037725
transform 1 0 102764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1117
timestamp 1676037725
transform 1 0 103868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1129
timestamp 1676037725
transform 1 0 104972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1141
timestamp 1676037725
transform 1 0 106076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1147
timestamp 1676037725
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1149
timestamp 1676037725
transform 1 0 106812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1161
timestamp 1676037725
transform 1 0 107916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1173
timestamp 1676037725
transform 1 0 109020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1185
timestamp 1676037725
transform 1 0 110124 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1197
timestamp 1676037725
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1203
timestamp 1676037725
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1205
timestamp 1676037725
transform 1 0 111964 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1217
timestamp 1676037725
transform 1 0 113068 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1221
timestamp 1676037725
transform 1 0 113436 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1231
timestamp 1676037725
transform 1 0 114356 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1237
timestamp 1676037725
transform 1 0 114908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1249
timestamp 1676037725
transform 1 0 116012 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1257
timestamp 1676037725
transform 1 0 116748 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1261
timestamp 1676037725
transform 1 0 117116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1273
timestamp 1676037725
transform 1 0 118220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1285
timestamp 1676037725
transform 1 0 119324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1297
timestamp 1676037725
transform 1 0 120428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1314
timestamp 1676037725
transform 1 0 121992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1317
timestamp 1676037725
transform 1 0 122268 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1321
timestamp 1676037725
transform 1 0 122636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1333
timestamp 1676037725
transform 1 0 123740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1345
timestamp 1676037725
transform 1 0 124844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1357
timestamp 1676037725
transform 1 0 125948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1369
timestamp 1676037725
transform 1 0 127052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1373
timestamp 1676037725
transform 1 0 127420 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1377
timestamp 1676037725
transform 1 0 127788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1389
timestamp 1676037725
transform 1 0 128892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1401
timestamp 1676037725
transform 1 0 129996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1413
timestamp 1676037725
transform 1 0 131100 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1424
timestamp 1676037725
transform 1 0 132112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1429
timestamp 1676037725
transform 1 0 132572 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1433
timestamp 1676037725
transform 1 0 132940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1445
timestamp 1676037725
transform 1 0 134044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1457
timestamp 1676037725
transform 1 0 135148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1469
timestamp 1676037725
transform 1 0 136252 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1479
timestamp 1676037725
transform 1 0 137172 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1483
timestamp 1676037725
transform 1 0 137540 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_1485
timestamp 1676037725
transform 1 0 137724 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1489
timestamp 1676037725
transform 1 0 138092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1501
timestamp 1676037725
transform 1 0 139196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1513
timestamp 1676037725
transform 1 0 140300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1525
timestamp 1676037725
transform 1 0 141404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1537
timestamp 1676037725
transform 1 0 142508 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1541
timestamp 1676037725
transform 1 0 142876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1553
timestamp 1676037725
transform 1 0 143980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1565
timestamp 1676037725
transform 1 0 145084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1577
timestamp 1676037725
transform 1 0 146188 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1589
timestamp 1676037725
transform 1 0 147292 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1595
timestamp 1676037725
transform 1 0 147844 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1597
timestamp 1676037725
transform 1 0 148028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1609
timestamp 1676037725
transform 1 0 149132 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1619
timestamp 1676037725
transform 1 0 150052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1631
timestamp 1676037725
transform 1 0 151156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1643
timestamp 1676037725
transform 1 0 152260 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1651
timestamp 1676037725
transform 1 0 152996 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1653
timestamp 1676037725
transform 1 0 153180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1665
timestamp 1676037725
transform 1 0 154284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1677
timestamp 1676037725
transform 1 0 155388 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1689
timestamp 1676037725
transform 1 0 156492 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1701
timestamp 1676037725
transform 1 0 157596 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1707
timestamp 1676037725
transform 1 0 158148 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1709
timestamp 1676037725
transform 1 0 158332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1721
timestamp 1676037725
transform 1 0 159436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1733
timestamp 1676037725
transform 1 0 160540 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1745
timestamp 1676037725
transform 1 0 161644 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1757
timestamp 1676037725
transform 1 0 162748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1763
timestamp 1676037725
transform 1 0 163300 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1765
timestamp 1676037725
transform 1 0 163484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1777
timestamp 1676037725
transform 1 0 164588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1789
timestamp 1676037725
transform 1 0 165692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1801
timestamp 1676037725
transform 1 0 166796 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1813
timestamp 1676037725
transform 1 0 167900 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1819
timestamp 1676037725
transform 1 0 168452 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1821
timestamp 1676037725
transform 1 0 168636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1833
timestamp 1676037725
transform 1 0 169740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1845
timestamp 1676037725
transform 1 0 170844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1857
timestamp 1676037725
transform 1 0 171948 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1869
timestamp 1676037725
transform 1 0 173052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1875
timestamp 1676037725
transform 1 0 173604 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1877
timestamp 1676037725
transform 1 0 173788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1889
timestamp 1676037725
transform 1 0 174892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1901
timestamp 1676037725
transform 1 0 175996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1913
timestamp 1676037725
transform 1 0 177100 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1925
timestamp 1676037725
transform 1 0 178204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1931
timestamp 1676037725
transform 1 0 178756 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1933
timestamp 1676037725
transform 1 0 178940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1945
timestamp 1676037725
transform 1 0 180044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1957
timestamp 1676037725
transform 1 0 181148 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1969
timestamp 1676037725
transform 1 0 182252 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1981
timestamp 1676037725
transform 1 0 183356 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1987
timestamp 1676037725
transform 1 0 183908 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1989
timestamp 1676037725
transform 1 0 184092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2001
timestamp 1676037725
transform 1 0 185196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2013
timestamp 1676037725
transform 1 0 186300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2025
timestamp 1676037725
transform 1 0 187404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2037
timestamp 1676037725
transform 1 0 188508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2043
timestamp 1676037725
transform 1 0 189060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2045
timestamp 1676037725
transform 1 0 189244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2057
timestamp 1676037725
transform 1 0 190348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2069
timestamp 1676037725
transform 1 0 191452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2081
timestamp 1676037725
transform 1 0 192556 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2093
timestamp 1676037725
transform 1 0 193660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2099
timestamp 1676037725
transform 1 0 194212 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2101
timestamp 1676037725
transform 1 0 194396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2113
timestamp 1676037725
transform 1 0 195500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2125
timestamp 1676037725
transform 1 0 196604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2137
timestamp 1676037725
transform 1 0 197708 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2149
timestamp 1676037725
transform 1 0 198812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2155
timestamp 1676037725
transform 1 0 199364 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2157
timestamp 1676037725
transform 1 0 199548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2169
timestamp 1676037725
transform 1 0 200652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2181
timestamp 1676037725
transform 1 0 201756 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2193
timestamp 1676037725
transform 1 0 202860 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2205
timestamp 1676037725
transform 1 0 203964 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2211
timestamp 1676037725
transform 1 0 204516 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2213
timestamp 1676037725
transform 1 0 204700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2225
timestamp 1676037725
transform 1 0 205804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2237
timestamp 1676037725
transform 1 0 206908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2249
timestamp 1676037725
transform 1 0 208012 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2261
timestamp 1676037725
transform 1 0 209116 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2267
timestamp 1676037725
transform 1 0 209668 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2269
timestamp 1676037725
transform 1 0 209852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2281
timestamp 1676037725
transform 1 0 210956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2293
timestamp 1676037725
transform 1 0 212060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2305
timestamp 1676037725
transform 1 0 213164 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2317
timestamp 1676037725
transform 1 0 214268 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2323
timestamp 1676037725
transform 1 0 214820 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2325
timestamp 1676037725
transform 1 0 215004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2337
timestamp 1676037725
transform 1 0 216108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2349
timestamp 1676037725
transform 1 0 217212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2361
timestamp 1676037725
transform 1 0 218316 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2373
timestamp 1676037725
transform 1 0 219420 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2379
timestamp 1676037725
transform 1 0 219972 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2381
timestamp 1676037725
transform 1 0 220156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2393
timestamp 1676037725
transform 1 0 221260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2405
timestamp 1676037725
transform 1 0 222364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2417
timestamp 1676037725
transform 1 0 223468 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2429
timestamp 1676037725
transform 1 0 224572 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2435
timestamp 1676037725
transform 1 0 225124 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2437
timestamp 1676037725
transform 1 0 225308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2449
timestamp 1676037725
transform 1 0 226412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2461
timestamp 1676037725
transform 1 0 227516 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2473
timestamp 1676037725
transform 1 0 228620 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2485
timestamp 1676037725
transform 1 0 229724 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2491
timestamp 1676037725
transform 1 0 230276 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2493
timestamp 1676037725
transform 1 0 230460 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2505
timestamp 1676037725
transform 1 0 231564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2517
timestamp 1676037725
transform 1 0 232668 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2529
timestamp 1676037725
transform 1 0 233772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2541
timestamp 1676037725
transform 1 0 234876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2547
timestamp 1676037725
transform 1 0 235428 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2549
timestamp 1676037725
transform 1 0 235612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2561
timestamp 1676037725
transform 1 0 236716 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2573
timestamp 1676037725
transform 1 0 237820 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2585
timestamp 1676037725
transform 1 0 238924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2597
timestamp 1676037725
transform 1 0 240028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2603
timestamp 1676037725
transform 1 0 240580 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2605
timestamp 1676037725
transform 1 0 240764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2617
timestamp 1676037725
transform 1 0 241868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2629
timestamp 1676037725
transform 1 0 242972 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2641
timestamp 1676037725
transform 1 0 244076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2653
timestamp 1676037725
transform 1 0 245180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2659
timestamp 1676037725
transform 1 0 245732 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2661
timestamp 1676037725
transform 1 0 245916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2673
timestamp 1676037725
transform 1 0 247020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2685
timestamp 1676037725
transform 1 0 248124 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2697
timestamp 1676037725
transform 1 0 249228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2709
timestamp 1676037725
transform 1 0 250332 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2715
timestamp 1676037725
transform 1 0 250884 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_2717
timestamp 1676037725
transform 1 0 251068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_2721
timestamp 1676037725
transform 1 0 251436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_2729
timestamp 1676037725
transform 1 0 252172 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2733
timestamp 1676037725
transform 1 0 252540 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2745
timestamp 1676037725
transform 1 0 253644 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2757
timestamp 1676037725
transform 1 0 254748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_2769
timestamp 1676037725
transform 1 0 255852 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2773
timestamp 1676037725
transform 1 0 256220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2785
timestamp 1676037725
transform 1 0 257324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2797
timestamp 1676037725
transform 1 0 258428 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2809
timestamp 1676037725
transform 1 0 259532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2821
timestamp 1676037725
transform 1 0 260636 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2827
timestamp 1676037725
transform 1 0 261188 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2829
timestamp 1676037725
transform 1 0 261372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2841
timestamp 1676037725
transform 1 0 262476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2853
timestamp 1676037725
transform 1 0 263580 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2865
timestamp 1676037725
transform 1 0 264684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2877
timestamp 1676037725
transform 1 0 265788 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2883
timestamp 1676037725
transform 1 0 266340 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2885
timestamp 1676037725
transform 1 0 266524 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2897
timestamp 1676037725
transform 1 0 267628 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2909
timestamp 1676037725
transform 1 0 268732 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2921
timestamp 1676037725
transform 1 0 269836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_2933
timestamp 1676037725
transform 1 0 270940 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_2939
timestamp 1676037725
transform 1 0 271492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2941
timestamp 1676037725
transform 1 0 271676 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2953
timestamp 1676037725
transform 1 0 272780 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_2965
timestamp 1676037725
transform 1 0 273884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_2977
timestamp 1676037725
transform 1 0 274988 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_2994
timestamp 1676037725
transform 1 0 276552 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_2997
timestamp 1676037725
transform 1 0 276828 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3001
timestamp 1676037725
transform 1 0 277196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3013
timestamp 1676037725
transform 1 0 278300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3025
timestamp 1676037725
transform 1 0 279404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3037
timestamp 1676037725
transform 1 0 280508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3050
timestamp 1676037725
transform 1 0 281704 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3053
timestamp 1676037725
transform 1 0 281980 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3057
timestamp 1676037725
transform 1 0 282348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3069
timestamp 1676037725
transform 1 0 283452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3081
timestamp 1676037725
transform 1 0 284556 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3093
timestamp 1676037725
transform 1 0 285660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3106
timestamp 1676037725
transform 1 0 286856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3109
timestamp 1676037725
transform 1 0 287132 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3113
timestamp 1676037725
transform 1 0 287500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3125
timestamp 1676037725
transform 1 0 288604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3137
timestamp 1676037725
transform 1 0 289708 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3149
timestamp 1676037725
transform 1 0 290812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3161
timestamp 1676037725
transform 1 0 291916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3165
timestamp 1676037725
transform 1 0 292284 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3169
timestamp 1676037725
transform 1 0 292652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3181
timestamp 1676037725
transform 1 0 293756 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3193
timestamp 1676037725
transform 1 0 294860 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3205
timestamp 1676037725
transform 1 0 295964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3215
timestamp 1676037725
transform 1 0 296884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3219
timestamp 1676037725
transform 1 0 297252 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3221
timestamp 1676037725
transform 1 0 297436 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3225
timestamp 1676037725
transform 1 0 297804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3237
timestamp 1676037725
transform 1 0 298908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3249
timestamp 1676037725
transform 1 0 300012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3261
timestamp 1676037725
transform 1 0 301116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3273
timestamp 1676037725
transform 1 0 302220 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3277
timestamp 1676037725
transform 1 0 302588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3289
timestamp 1676037725
transform 1 0 303692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3301
timestamp 1676037725
transform 1 0 304796 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3313
timestamp 1676037725
transform 1 0 305900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3325
timestamp 1676037725
transform 1 0 307004 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3331
timestamp 1676037725
transform 1 0 307556 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3333
timestamp 1676037725
transform 1 0 307740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3345
timestamp 1676037725
transform 1 0 308844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3357
timestamp 1676037725
transform 1 0 309948 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3369
timestamp 1676037725
transform 1 0 311052 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3381
timestamp 1676037725
transform 1 0 312156 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3387
timestamp 1676037725
transform 1 0 312708 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3389
timestamp 1676037725
transform 1 0 312892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3401
timestamp 1676037725
transform 1 0 313996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3413
timestamp 1676037725
transform 1 0 315100 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3425
timestamp 1676037725
transform 1 0 316204 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3437
timestamp 1676037725
transform 1 0 317308 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3443
timestamp 1676037725
transform 1 0 317860 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3445
timestamp 1676037725
transform 1 0 318044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3457
timestamp 1676037725
transform 1 0 319148 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3469
timestamp 1676037725
transform 1 0 320252 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3481
timestamp 1676037725
transform 1 0 321356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3493
timestamp 1676037725
transform 1 0 322460 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3499
timestamp 1676037725
transform 1 0 323012 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3501
timestamp 1676037725
transform 1 0 323196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3513
timestamp 1676037725
transform 1 0 324300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3525
timestamp 1676037725
transform 1 0 325404 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3537
timestamp 1676037725
transform 1 0 326508 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3549
timestamp 1676037725
transform 1 0 327612 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3555
timestamp 1676037725
transform 1 0 328164 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3557
timestamp 1676037725
transform 1 0 328348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3569
timestamp 1676037725
transform 1 0 329452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3581
timestamp 1676037725
transform 1 0 330556 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3593
timestamp 1676037725
transform 1 0 331660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3605
timestamp 1676037725
transform 1 0 332764 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3611
timestamp 1676037725
transform 1 0 333316 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3613
timestamp 1676037725
transform 1 0 333500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3625
timestamp 1676037725
transform 1 0 334604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3637
timestamp 1676037725
transform 1 0 335708 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3649
timestamp 1676037725
transform 1 0 336812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3661
timestamp 1676037725
transform 1 0 337916 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3667
timestamp 1676037725
transform 1 0 338468 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3669
timestamp 1676037725
transform 1 0 338652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3681
timestamp 1676037725
transform 1 0 339756 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3693
timestamp 1676037725
transform 1 0 340860 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3705
timestamp 1676037725
transform 1 0 341964 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3717
timestamp 1676037725
transform 1 0 343068 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3723
timestamp 1676037725
transform 1 0 343620 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3725
timestamp 1676037725
transform 1 0 343804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3737
timestamp 1676037725
transform 1 0 344908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3749
timestamp 1676037725
transform 1 0 346012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3761
timestamp 1676037725
transform 1 0 347116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3773
timestamp 1676037725
transform 1 0 348220 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3779
timestamp 1676037725
transform 1 0 348772 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3781
timestamp 1676037725
transform 1 0 348956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3793
timestamp 1676037725
transform 1 0 350060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3805
timestamp 1676037725
transform 1 0 351164 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3817
timestamp 1676037725
transform 1 0 352268 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3829
timestamp 1676037725
transform 1 0 353372 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3835
timestamp 1676037725
transform 1 0 353924 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3837
timestamp 1676037725
transform 1 0 354108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3849
timestamp 1676037725
transform 1 0 355212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3861
timestamp 1676037725
transform 1 0 356316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3873
timestamp 1676037725
transform 1 0 357420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3885
timestamp 1676037725
transform 1 0 358524 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3891
timestamp 1676037725
transform 1 0 359076 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3893
timestamp 1676037725
transform 1 0 359260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3905
timestamp 1676037725
transform 1 0 360364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3917
timestamp 1676037725
transform 1 0 361468 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3929
timestamp 1676037725
transform 1 0 362572 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3941
timestamp 1676037725
transform 1 0 363676 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3947
timestamp 1676037725
transform 1 0 364228 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3949
timestamp 1676037725
transform 1 0 364412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3961
timestamp 1676037725
transform 1 0 365516 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3973
timestamp 1676037725
transform 1 0 366620 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3985
timestamp 1676037725
transform 1 0 367724 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3997
timestamp 1676037725
transform 1 0 368828 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4003
timestamp 1676037725
transform 1 0 369380 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4005
timestamp 1676037725
transform 1 0 369564 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4017
timestamp 1676037725
transform 1 0 370668 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4029
timestamp 1676037725
transform 1 0 371772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4041
timestamp 1676037725
transform 1 0 372876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4053
timestamp 1676037725
transform 1 0 373980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4059
timestamp 1676037725
transform 1 0 374532 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4061
timestamp 1676037725
transform 1 0 374716 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4073
timestamp 1676037725
transform 1 0 375820 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4085
timestamp 1676037725
transform 1 0 376924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4097
timestamp 1676037725
transform 1 0 378028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4109
timestamp 1676037725
transform 1 0 379132 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4115
timestamp 1676037725
transform 1 0 379684 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4117
timestamp 1676037725
transform 1 0 379868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4129
timestamp 1676037725
transform 1 0 380972 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4141
timestamp 1676037725
transform 1 0 382076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4153
timestamp 1676037725
transform 1 0 383180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4165
timestamp 1676037725
transform 1 0 384284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4171
timestamp 1676037725
transform 1 0 384836 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4173
timestamp 1676037725
transform 1 0 385020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4185
timestamp 1676037725
transform 1 0 386124 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4197
timestamp 1676037725
transform 1 0 387228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4209
timestamp 1676037725
transform 1 0 388332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4221
timestamp 1676037725
transform 1 0 389436 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4227
timestamp 1676037725
transform 1 0 389988 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4229
timestamp 1676037725
transform 1 0 390172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4241
timestamp 1676037725
transform 1 0 391276 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4253
timestamp 1676037725
transform 1 0 392380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4265
timestamp 1676037725
transform 1 0 393484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4277
timestamp 1676037725
transform 1 0 394588 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4283
timestamp 1676037725
transform 1 0 395140 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4285
timestamp 1676037725
transform 1 0 395324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4297
timestamp 1676037725
transform 1 0 396428 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4309
timestamp 1676037725
transform 1 0 397532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4321
timestamp 1676037725
transform 1 0 398636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4333
timestamp 1676037725
transform 1 0 399740 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4339
timestamp 1676037725
transform 1 0 400292 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4341
timestamp 1676037725
transform 1 0 400476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4353
timestamp 1676037725
transform 1 0 401580 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4365
timestamp 1676037725
transform 1 0 402684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4377
timestamp 1676037725
transform 1 0 403788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4389
timestamp 1676037725
transform 1 0 404892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4395
timestamp 1676037725
transform 1 0 405444 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4397
timestamp 1676037725
transform 1 0 405628 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4409
timestamp 1676037725
transform 1 0 406732 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4421
timestamp 1676037725
transform 1 0 407836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4433
timestamp 1676037725
transform 1 0 408940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4445
timestamp 1676037725
transform 1 0 410044 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4451
timestamp 1676037725
transform 1 0 410596 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4453
timestamp 1676037725
transform 1 0 410780 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4465
timestamp 1676037725
transform 1 0 411884 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4477
timestamp 1676037725
transform 1 0 412988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4489
timestamp 1676037725
transform 1 0 414092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4501
timestamp 1676037725
transform 1 0 415196 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4507
timestamp 1676037725
transform 1 0 415748 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4509
timestamp 1676037725
transform 1 0 415932 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4521
timestamp 1676037725
transform 1 0 417036 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4533
timestamp 1676037725
transform 1 0 418140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4545
timestamp 1676037725
transform 1 0 419244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4557
timestamp 1676037725
transform 1 0 420348 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4563
timestamp 1676037725
transform 1 0 420900 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4565
timestamp 1676037725
transform 1 0 421084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4577
timestamp 1676037725
transform 1 0 422188 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4589
timestamp 1676037725
transform 1 0 423292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4601
timestamp 1676037725
transform 1 0 424396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4613
timestamp 1676037725
transform 1 0 425500 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4619
timestamp 1676037725
transform 1 0 426052 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4621
timestamp 1676037725
transform 1 0 426236 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4633
timestamp 1676037725
transform 1 0 427340 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4645
timestamp 1676037725
transform 1 0 428444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4657
timestamp 1676037725
transform 1 0 429548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4669
timestamp 1676037725
transform 1 0 430652 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4675
timestamp 1676037725
transform 1 0 431204 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4677
timestamp 1676037725
transform 1 0 431388 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4689
timestamp 1676037725
transform 1 0 432492 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4701
timestamp 1676037725
transform 1 0 433596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4713
timestamp 1676037725
transform 1 0 434700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4725
timestamp 1676037725
transform 1 0 435804 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4731
timestamp 1676037725
transform 1 0 436356 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4733
timestamp 1676037725
transform 1 0 436540 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4745
timestamp 1676037725
transform 1 0 437644 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4757
timestamp 1676037725
transform 1 0 438748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4769
timestamp 1676037725
transform 1 0 439852 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4781
timestamp 1676037725
transform 1 0 440956 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4787
timestamp 1676037725
transform 1 0 441508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4789
timestamp 1676037725
transform 1 0 441692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4801
timestamp 1676037725
transform 1 0 442796 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4813
timestamp 1676037725
transform 1 0 443900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4825
timestamp 1676037725
transform 1 0 445004 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4837
timestamp 1676037725
transform 1 0 446108 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4843
timestamp 1676037725
transform 1 0 446660 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4845
timestamp 1676037725
transform 1 0 446844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4857
timestamp 1676037725
transform 1 0 447948 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4869
timestamp 1676037725
transform 1 0 449052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4881
timestamp 1676037725
transform 1 0 450156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4893
timestamp 1676037725
transform 1 0 451260 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4899
timestamp 1676037725
transform 1 0 451812 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4901
timestamp 1676037725
transform 1 0 451996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4913
timestamp 1676037725
transform 1 0 453100 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4925
timestamp 1676037725
transform 1 0 454204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4937
timestamp 1676037725
transform 1 0 455308 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_4949
timestamp 1676037725
transform 1 0 456412 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_4955
timestamp 1676037725
transform 1 0 456964 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4957
timestamp 1676037725
transform 1 0 457148 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4969
timestamp 1676037725
transform 1 0 458252 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4981
timestamp 1676037725
transform 1 0 459356 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_4993
timestamp 1676037725
transform 1 0 460460 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5005
timestamp 1676037725
transform 1 0 461564 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5011
timestamp 1676037725
transform 1 0 462116 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5013
timestamp 1676037725
transform 1 0 462300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5025
timestamp 1676037725
transform 1 0 463404 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5037
timestamp 1676037725
transform 1 0 464508 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5049
timestamp 1676037725
transform 1 0 465612 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5061
timestamp 1676037725
transform 1 0 466716 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5067
timestamp 1676037725
transform 1 0 467268 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5069
timestamp 1676037725
transform 1 0 467452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5081
timestamp 1676037725
transform 1 0 468556 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5093
timestamp 1676037725
transform 1 0 469660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5105
timestamp 1676037725
transform 1 0 470764 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5117
timestamp 1676037725
transform 1 0 471868 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5123
timestamp 1676037725
transform 1 0 472420 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5125
timestamp 1676037725
transform 1 0 472604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5137
timestamp 1676037725
transform 1 0 473708 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5149
timestamp 1676037725
transform 1 0 474812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5161
timestamp 1676037725
transform 1 0 475916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5173
timestamp 1676037725
transform 1 0 477020 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5179
timestamp 1676037725
transform 1 0 477572 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5181
timestamp 1676037725
transform 1 0 477756 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5193
timestamp 1676037725
transform 1 0 478860 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5205
timestamp 1676037725
transform 1 0 479964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5217
timestamp 1676037725
transform 1 0 481068 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5229
timestamp 1676037725
transform 1 0 482172 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5235
timestamp 1676037725
transform 1 0 482724 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5237
timestamp 1676037725
transform 1 0 482908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5249
timestamp 1676037725
transform 1 0 484012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5261
timestamp 1676037725
transform 1 0 485116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5273
timestamp 1676037725
transform 1 0 486220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5285
timestamp 1676037725
transform 1 0 487324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5291
timestamp 1676037725
transform 1 0 487876 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5293
timestamp 1676037725
transform 1 0 488060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5305
timestamp 1676037725
transform 1 0 489164 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5317
timestamp 1676037725
transform 1 0 490268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5329
timestamp 1676037725
transform 1 0 491372 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5341
timestamp 1676037725
transform 1 0 492476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5347
timestamp 1676037725
transform 1 0 493028 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5349
timestamp 1676037725
transform 1 0 493212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5361
timestamp 1676037725
transform 1 0 494316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5373
timestamp 1676037725
transform 1 0 495420 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5385
timestamp 1676037725
transform 1 0 496524 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5397
timestamp 1676037725
transform 1 0 497628 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5403
timestamp 1676037725
transform 1 0 498180 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5405
timestamp 1676037725
transform 1 0 498364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5417
timestamp 1676037725
transform 1 0 499468 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5429
timestamp 1676037725
transform 1 0 500572 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5441
timestamp 1676037725
transform 1 0 501676 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5453
timestamp 1676037725
transform 1 0 502780 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5459
timestamp 1676037725
transform 1 0 503332 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5461
timestamp 1676037725
transform 1 0 503516 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5473
timestamp 1676037725
transform 1 0 504620 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5485
timestamp 1676037725
transform 1 0 505724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5497
timestamp 1676037725
transform 1 0 506828 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5509
timestamp 1676037725
transform 1 0 507932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5515
timestamp 1676037725
transform 1 0 508484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5517
timestamp 1676037725
transform 1 0 508668 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5529
timestamp 1676037725
transform 1 0 509772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5541
timestamp 1676037725
transform 1 0 510876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5553
timestamp 1676037725
transform 1 0 511980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5565
timestamp 1676037725
transform 1 0 513084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5571
timestamp 1676037725
transform 1 0 513636 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5573
timestamp 1676037725
transform 1 0 513820 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5585
timestamp 1676037725
transform 1 0 514924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5597
timestamp 1676037725
transform 1 0 516028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5609
timestamp 1676037725
transform 1 0 517132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5621
timestamp 1676037725
transform 1 0 518236 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5627
timestamp 1676037725
transform 1 0 518788 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5629
timestamp 1676037725
transform 1 0 518972 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5641
timestamp 1676037725
transform 1 0 520076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5653
timestamp 1676037725
transform 1 0 521180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5665
timestamp 1676037725
transform 1 0 522284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_5677
timestamp 1676037725
transform 1 0 523388 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5683
timestamp 1676037725
transform 1 0 523940 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5685
timestamp 1676037725
transform 1 0 524124 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5697
timestamp 1676037725
transform 1 0 525228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5709
timestamp 1676037725
transform 1 0 526332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_5721
timestamp 1676037725
transform 1 0 527436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1676037725
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1676037725
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1676037725
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1676037725
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1676037725
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1676037725
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1676037725
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1676037725
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1676037725
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1676037725
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1676037725
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1676037725
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1676037725
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1676037725
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1676037725
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1676037725
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1676037725
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1676037725
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1676037725
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1676037725
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1676037725
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1676037725
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1676037725
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1676037725
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1676037725
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1676037725
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1676037725
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1676037725
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1676037725
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1676037725
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1676037725
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_821
timestamp 1676037725
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1676037725
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1676037725
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_841
timestamp 1676037725
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_853
timestamp 1676037725
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_865
timestamp 1676037725
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_877
timestamp 1676037725
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1676037725
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1676037725
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_897
timestamp 1676037725
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_909
timestamp 1676037725
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_921
timestamp 1676037725
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_933
timestamp 1676037725
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_945
timestamp 1676037725
transform 1 0 88044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1676037725
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_953
timestamp 1676037725
transform 1 0 88780 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_965
timestamp 1676037725
transform 1 0 89884 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_977
timestamp 1676037725
transform 1 0 90988 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_989
timestamp 1676037725
transform 1 0 92092 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1001
timestamp 1676037725
transform 1 0 93196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1007
timestamp 1676037725
transform 1 0 93748 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1009
timestamp 1676037725
transform 1 0 93932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1021
timestamp 1676037725
transform 1 0 95036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1033
timestamp 1676037725
transform 1 0 96140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1045
timestamp 1676037725
transform 1 0 97244 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1057
timestamp 1676037725
transform 1 0 98348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1063
timestamp 1676037725
transform 1 0 98900 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1065
timestamp 1676037725
transform 1 0 99084 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1077
timestamp 1676037725
transform 1 0 100188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1089
timestamp 1676037725
transform 1 0 101292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1101
timestamp 1676037725
transform 1 0 102396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1113
timestamp 1676037725
transform 1 0 103500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1119
timestamp 1676037725
transform 1 0 104052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1121
timestamp 1676037725
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1133
timestamp 1676037725
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1145
timestamp 1676037725
transform 1 0 106444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1157
timestamp 1676037725
transform 1 0 107548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1169
timestamp 1676037725
transform 1 0 108652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1175
timestamp 1676037725
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1177
timestamp 1676037725
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1189
timestamp 1676037725
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1201
timestamp 1676037725
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1213
timestamp 1676037725
transform 1 0 112700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1225
timestamp 1676037725
transform 1 0 113804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1231
timestamp 1676037725
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1233
timestamp 1676037725
transform 1 0 114540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1245
timestamp 1676037725
transform 1 0 115644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1257
timestamp 1676037725
transform 1 0 116748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1269
timestamp 1676037725
transform 1 0 117852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1281
timestamp 1676037725
transform 1 0 118956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1287
timestamp 1676037725
transform 1 0 119508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1289
timestamp 1676037725
transform 1 0 119692 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1301
timestamp 1676037725
transform 1 0 120796 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1313
timestamp 1676037725
transform 1 0 121900 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1325
timestamp 1676037725
transform 1 0 123004 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1337
timestamp 1676037725
transform 1 0 124108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1343
timestamp 1676037725
transform 1 0 124660 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1345
timestamp 1676037725
transform 1 0 124844 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1357
timestamp 1676037725
transform 1 0 125948 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1369
timestamp 1676037725
transform 1 0 127052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1381
timestamp 1676037725
transform 1 0 128156 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1393
timestamp 1676037725
transform 1 0 129260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1399
timestamp 1676037725
transform 1 0 129812 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1401
timestamp 1676037725
transform 1 0 129996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1413
timestamp 1676037725
transform 1 0 131100 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1425
timestamp 1676037725
transform 1 0 132204 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1437
timestamp 1676037725
transform 1 0 133308 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1449
timestamp 1676037725
transform 1 0 134412 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1455
timestamp 1676037725
transform 1 0 134964 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1457
timestamp 1676037725
transform 1 0 135148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1469
timestamp 1676037725
transform 1 0 136252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1481
timestamp 1676037725
transform 1 0 137356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1493
timestamp 1676037725
transform 1 0 138460 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1505
timestamp 1676037725
transform 1 0 139564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1511
timestamp 1676037725
transform 1 0 140116 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1513
timestamp 1676037725
transform 1 0 140300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1534
timestamp 1676037725
transform 1 0 142232 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1540
timestamp 1676037725
transform 1 0 142784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1552
timestamp 1676037725
transform 1 0 143888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1556
timestamp 1676037725
transform 1 0 144256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1566
timestamp 1676037725
transform 1 0 145176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1569
timestamp 1676037725
transform 1 0 145452 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1573
timestamp 1676037725
transform 1 0 145820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1585
timestamp 1676037725
transform 1 0 146924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1597
timestamp 1676037725
transform 1 0 148028 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_1605
timestamp 1676037725
transform 1 0 148764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1617
timestamp 1676037725
transform 1 0 149868 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1623
timestamp 1676037725
transform 1 0 150420 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1625
timestamp 1676037725
transform 1 0 150604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1637
timestamp 1676037725
transform 1 0 151708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1649
timestamp 1676037725
transform 1 0 152812 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1661
timestamp 1676037725
transform 1 0 153916 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1673
timestamp 1676037725
transform 1 0 155020 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1679
timestamp 1676037725
transform 1 0 155572 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1681
timestamp 1676037725
transform 1 0 155756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1689
timestamp 1676037725
transform 1 0 156492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1699
timestamp 1676037725
transform 1 0 157412 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1705
timestamp 1676037725
transform 1 0 157964 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1717
timestamp 1676037725
transform 1 0 159068 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1729
timestamp 1676037725
transform 1 0 160172 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1735
timestamp 1676037725
transform 1 0 160724 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1737
timestamp 1676037725
transform 1 0 160908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1749
timestamp 1676037725
transform 1 0 162012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1761
timestamp 1676037725
transform 1 0 163116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1782
timestamp 1676037725
transform 1 0 165048 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1788
timestamp 1676037725
transform 1 0 165600 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1793
timestamp 1676037725
transform 1 0 166060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1805
timestamp 1676037725
transform 1 0 167164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1817
timestamp 1676037725
transform 1 0 168268 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1829
timestamp 1676037725
transform 1 0 169372 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1841
timestamp 1676037725
transform 1 0 170476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1847
timestamp 1676037725
transform 1 0 171028 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1849
timestamp 1676037725
transform 1 0 171212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1861
timestamp 1676037725
transform 1 0 172316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1873
timestamp 1676037725
transform 1 0 173420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1885
timestamp 1676037725
transform 1 0 174524 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1897
timestamp 1676037725
transform 1 0 175628 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1903
timestamp 1676037725
transform 1 0 176180 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1905
timestamp 1676037725
transform 1 0 176364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1917
timestamp 1676037725
transform 1 0 177468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1929
timestamp 1676037725
transform 1 0 178572 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1941
timestamp 1676037725
transform 1 0 179676 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1953
timestamp 1676037725
transform 1 0 180780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1959
timestamp 1676037725
transform 1 0 181332 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1961
timestamp 1676037725
transform 1 0 181516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1973
timestamp 1676037725
transform 1 0 182620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1985
timestamp 1676037725
transform 1 0 183724 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1997
timestamp 1676037725
transform 1 0 184828 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2009
timestamp 1676037725
transform 1 0 185932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2015
timestamp 1676037725
transform 1 0 186484 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2017
timestamp 1676037725
transform 1 0 186668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2029
timestamp 1676037725
transform 1 0 187772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2041
timestamp 1676037725
transform 1 0 188876 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2053
timestamp 1676037725
transform 1 0 189980 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2065
timestamp 1676037725
transform 1 0 191084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2071
timestamp 1676037725
transform 1 0 191636 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2073
timestamp 1676037725
transform 1 0 191820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2085
timestamp 1676037725
transform 1 0 192924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2097
timestamp 1676037725
transform 1 0 194028 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2109
timestamp 1676037725
transform 1 0 195132 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2121
timestamp 1676037725
transform 1 0 196236 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2127
timestamp 1676037725
transform 1 0 196788 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2129
timestamp 1676037725
transform 1 0 196972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2141
timestamp 1676037725
transform 1 0 198076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2153
timestamp 1676037725
transform 1 0 199180 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2165
timestamp 1676037725
transform 1 0 200284 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2177
timestamp 1676037725
transform 1 0 201388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2183
timestamp 1676037725
transform 1 0 201940 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2185
timestamp 1676037725
transform 1 0 202124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2197
timestamp 1676037725
transform 1 0 203228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2209
timestamp 1676037725
transform 1 0 204332 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2221
timestamp 1676037725
transform 1 0 205436 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2233
timestamp 1676037725
transform 1 0 206540 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2239
timestamp 1676037725
transform 1 0 207092 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2241
timestamp 1676037725
transform 1 0 207276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2253
timestamp 1676037725
transform 1 0 208380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2265
timestamp 1676037725
transform 1 0 209484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2277
timestamp 1676037725
transform 1 0 210588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2289
timestamp 1676037725
transform 1 0 211692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2295
timestamp 1676037725
transform 1 0 212244 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2297
timestamp 1676037725
transform 1 0 212428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2309
timestamp 1676037725
transform 1 0 213532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2321
timestamp 1676037725
transform 1 0 214636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2333
timestamp 1676037725
transform 1 0 215740 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2345
timestamp 1676037725
transform 1 0 216844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2351
timestamp 1676037725
transform 1 0 217396 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2353
timestamp 1676037725
transform 1 0 217580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2365
timestamp 1676037725
transform 1 0 218684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2377
timestamp 1676037725
transform 1 0 219788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2389
timestamp 1676037725
transform 1 0 220892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2401
timestamp 1676037725
transform 1 0 221996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2407
timestamp 1676037725
transform 1 0 222548 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2409
timestamp 1676037725
transform 1 0 222732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2421
timestamp 1676037725
transform 1 0 223836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2433
timestamp 1676037725
transform 1 0 224940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2445
timestamp 1676037725
transform 1 0 226044 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2457
timestamp 1676037725
transform 1 0 227148 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2463
timestamp 1676037725
transform 1 0 227700 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2465
timestamp 1676037725
transform 1 0 227884 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2477
timestamp 1676037725
transform 1 0 228988 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2489
timestamp 1676037725
transform 1 0 230092 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2501
timestamp 1676037725
transform 1 0 231196 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2513
timestamp 1676037725
transform 1 0 232300 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2519
timestamp 1676037725
transform 1 0 232852 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2521
timestamp 1676037725
transform 1 0 233036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2533
timestamp 1676037725
transform 1 0 234140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2545
timestamp 1676037725
transform 1 0 235244 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2557
timestamp 1676037725
transform 1 0 236348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2569
timestamp 1676037725
transform 1 0 237452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2575
timestamp 1676037725
transform 1 0 238004 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2577
timestamp 1676037725
transform 1 0 238188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2589
timestamp 1676037725
transform 1 0 239292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2601
timestamp 1676037725
transform 1 0 240396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2613
timestamp 1676037725
transform 1 0 241500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2625
timestamp 1676037725
transform 1 0 242604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2631
timestamp 1676037725
transform 1 0 243156 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2633
timestamp 1676037725
transform 1 0 243340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2645
timestamp 1676037725
transform 1 0 244444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2657
timestamp 1676037725
transform 1 0 245548 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2669
timestamp 1676037725
transform 1 0 246652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2681
timestamp 1676037725
transform 1 0 247756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2687
timestamp 1676037725
transform 1 0 248308 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2689
timestamp 1676037725
transform 1 0 248492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2701
timestamp 1676037725
transform 1 0 249596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2713
timestamp 1676037725
transform 1 0 250700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2725
timestamp 1676037725
transform 1 0 251804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2737
timestamp 1676037725
transform 1 0 252908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2743
timestamp 1676037725
transform 1 0 253460 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2745
timestamp 1676037725
transform 1 0 253644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2757
timestamp 1676037725
transform 1 0 254748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2769
timestamp 1676037725
transform 1 0 255852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2781
timestamp 1676037725
transform 1 0 256956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2793
timestamp 1676037725
transform 1 0 258060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2799
timestamp 1676037725
transform 1 0 258612 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2801
timestamp 1676037725
transform 1 0 258796 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2813
timestamp 1676037725
transform 1 0 259900 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2825
timestamp 1676037725
transform 1 0 261004 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2837
timestamp 1676037725
transform 1 0 262108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2849
timestamp 1676037725
transform 1 0 263212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2855
timestamp 1676037725
transform 1 0 263764 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2857
timestamp 1676037725
transform 1 0 263948 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2869
timestamp 1676037725
transform 1 0 265052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2881
timestamp 1676037725
transform 1 0 266156 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2893
timestamp 1676037725
transform 1 0 267260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2905
timestamp 1676037725
transform 1 0 268364 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2911
timestamp 1676037725
transform 1 0 268916 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2913
timestamp 1676037725
transform 1 0 269100 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2925
timestamp 1676037725
transform 1 0 270204 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2937
timestamp 1676037725
transform 1 0 271308 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2949
timestamp 1676037725
transform 1 0 272412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_2961
timestamp 1676037725
transform 1 0 273516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_2967
timestamp 1676037725
transform 1 0 274068 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2969
timestamp 1676037725
transform 1 0 274252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2981
timestamp 1676037725
transform 1 0 275356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_2993
timestamp 1676037725
transform 1 0 276460 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3005
timestamp 1676037725
transform 1 0 277564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3017
timestamp 1676037725
transform 1 0 278668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3023
timestamp 1676037725
transform 1 0 279220 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3025
timestamp 1676037725
transform 1 0 279404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3037
timestamp 1676037725
transform 1 0 280508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3049
timestamp 1676037725
transform 1 0 281612 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3061
timestamp 1676037725
transform 1 0 282716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3073
timestamp 1676037725
transform 1 0 283820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3079
timestamp 1676037725
transform 1 0 284372 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3081
timestamp 1676037725
transform 1 0 284556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3093
timestamp 1676037725
transform 1 0 285660 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3105
timestamp 1676037725
transform 1 0 286764 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3117
timestamp 1676037725
transform 1 0 287868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3129
timestamp 1676037725
transform 1 0 288972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3135
timestamp 1676037725
transform 1 0 289524 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3137
timestamp 1676037725
transform 1 0 289708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3149
timestamp 1676037725
transform 1 0 290812 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3161
timestamp 1676037725
transform 1 0 291916 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3173
timestamp 1676037725
transform 1 0 293020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3185
timestamp 1676037725
transform 1 0 294124 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3191
timestamp 1676037725
transform 1 0 294676 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3193
timestamp 1676037725
transform 1 0 294860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3205
timestamp 1676037725
transform 1 0 295964 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3217
timestamp 1676037725
transform 1 0 297068 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3229
timestamp 1676037725
transform 1 0 298172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3241
timestamp 1676037725
transform 1 0 299276 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3247
timestamp 1676037725
transform 1 0 299828 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3249
timestamp 1676037725
transform 1 0 300012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3270
timestamp 1676037725
transform 1 0 301944 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3276
timestamp 1676037725
transform 1 0 302496 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3288
timestamp 1676037725
transform 1 0 303600 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3300
timestamp 1676037725
transform 1 0 304704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3305
timestamp 1676037725
transform 1 0 305164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3313
timestamp 1676037725
transform 1 0 305900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3325
timestamp 1676037725
transform 1 0 307004 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3331
timestamp 1676037725
transform 1 0 307556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3343
timestamp 1676037725
transform 1 0 308660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3355
timestamp 1676037725
transform 1 0 309764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3359
timestamp 1676037725
transform 1 0 310132 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3361
timestamp 1676037725
transform 1 0 310316 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3369
timestamp 1676037725
transform 1 0 311052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3379
timestamp 1676037725
transform 1 0 311972 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3385
timestamp 1676037725
transform 1 0 312524 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3397
timestamp 1676037725
transform 1 0 313628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3409
timestamp 1676037725
transform 1 0 314732 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3415
timestamp 1676037725
transform 1 0 315284 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3417
timestamp 1676037725
transform 1 0 315468 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3434
timestamp 1676037725
transform 1 0 317032 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3440
timestamp 1676037725
transform 1 0 317584 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3452
timestamp 1676037725
transform 1 0 318688 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3464
timestamp 1676037725
transform 1 0 319792 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3473
timestamp 1676037725
transform 1 0 320620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3485
timestamp 1676037725
transform 1 0 321724 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3497
timestamp 1676037725
transform 1 0 322828 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3509
timestamp 1676037725
transform 1 0 323932 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3521
timestamp 1676037725
transform 1 0 325036 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3527
timestamp 1676037725
transform 1 0 325588 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3529
timestamp 1676037725
transform 1 0 325772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3541
timestamp 1676037725
transform 1 0 326876 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3553
timestamp 1676037725
transform 1 0 327980 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3565
timestamp 1676037725
transform 1 0 329084 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3577
timestamp 1676037725
transform 1 0 330188 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3583
timestamp 1676037725
transform 1 0 330740 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3585
timestamp 1676037725
transform 1 0 330924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3597
timestamp 1676037725
transform 1 0 332028 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3609
timestamp 1676037725
transform 1 0 333132 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3621
timestamp 1676037725
transform 1 0 334236 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3633
timestamp 1676037725
transform 1 0 335340 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3639
timestamp 1676037725
transform 1 0 335892 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3641
timestamp 1676037725
transform 1 0 336076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3653
timestamp 1676037725
transform 1 0 337180 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3665
timestamp 1676037725
transform 1 0 338284 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3677
timestamp 1676037725
transform 1 0 339388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3689
timestamp 1676037725
transform 1 0 340492 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3695
timestamp 1676037725
transform 1 0 341044 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3697
timestamp 1676037725
transform 1 0 341228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3709
timestamp 1676037725
transform 1 0 342332 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3721
timestamp 1676037725
transform 1 0 343436 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3733
timestamp 1676037725
transform 1 0 344540 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3745
timestamp 1676037725
transform 1 0 345644 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3751
timestamp 1676037725
transform 1 0 346196 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3753
timestamp 1676037725
transform 1 0 346380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3765
timestamp 1676037725
transform 1 0 347484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3777
timestamp 1676037725
transform 1 0 348588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3789
timestamp 1676037725
transform 1 0 349692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3801
timestamp 1676037725
transform 1 0 350796 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3807
timestamp 1676037725
transform 1 0 351348 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3809
timestamp 1676037725
transform 1 0 351532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3821
timestamp 1676037725
transform 1 0 352636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3833
timestamp 1676037725
transform 1 0 353740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3845
timestamp 1676037725
transform 1 0 354844 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3857
timestamp 1676037725
transform 1 0 355948 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3863
timestamp 1676037725
transform 1 0 356500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3865
timestamp 1676037725
transform 1 0 356684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3877
timestamp 1676037725
transform 1 0 357788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3889
timestamp 1676037725
transform 1 0 358892 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3901
timestamp 1676037725
transform 1 0 359996 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3913
timestamp 1676037725
transform 1 0 361100 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3919
timestamp 1676037725
transform 1 0 361652 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3921
timestamp 1676037725
transform 1 0 361836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3933
timestamp 1676037725
transform 1 0 362940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3945
timestamp 1676037725
transform 1 0 364044 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3957
timestamp 1676037725
transform 1 0 365148 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3969
timestamp 1676037725
transform 1 0 366252 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3975
timestamp 1676037725
transform 1 0 366804 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3977
timestamp 1676037725
transform 1 0 366988 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3989
timestamp 1676037725
transform 1 0 368092 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4001
timestamp 1676037725
transform 1 0 369196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4013
timestamp 1676037725
transform 1 0 370300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4025
timestamp 1676037725
transform 1 0 371404 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4031
timestamp 1676037725
transform 1 0 371956 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4033
timestamp 1676037725
transform 1 0 372140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4045
timestamp 1676037725
transform 1 0 373244 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4057
timestamp 1676037725
transform 1 0 374348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4069
timestamp 1676037725
transform 1 0 375452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4081
timestamp 1676037725
transform 1 0 376556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4087
timestamp 1676037725
transform 1 0 377108 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4089
timestamp 1676037725
transform 1 0 377292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4101
timestamp 1676037725
transform 1 0 378396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4113
timestamp 1676037725
transform 1 0 379500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4125
timestamp 1676037725
transform 1 0 380604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4137
timestamp 1676037725
transform 1 0 381708 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4143
timestamp 1676037725
transform 1 0 382260 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4145
timestamp 1676037725
transform 1 0 382444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4157
timestamp 1676037725
transform 1 0 383548 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4169
timestamp 1676037725
transform 1 0 384652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4181
timestamp 1676037725
transform 1 0 385756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4193
timestamp 1676037725
transform 1 0 386860 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4199
timestamp 1676037725
transform 1 0 387412 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4201
timestamp 1676037725
transform 1 0 387596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4213
timestamp 1676037725
transform 1 0 388700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4225
timestamp 1676037725
transform 1 0 389804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4237
timestamp 1676037725
transform 1 0 390908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4249
timestamp 1676037725
transform 1 0 392012 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4255
timestamp 1676037725
transform 1 0 392564 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4257
timestamp 1676037725
transform 1 0 392748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4269
timestamp 1676037725
transform 1 0 393852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4281
timestamp 1676037725
transform 1 0 394956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4293
timestamp 1676037725
transform 1 0 396060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4305
timestamp 1676037725
transform 1 0 397164 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4311
timestamp 1676037725
transform 1 0 397716 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4313
timestamp 1676037725
transform 1 0 397900 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4325
timestamp 1676037725
transform 1 0 399004 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4337
timestamp 1676037725
transform 1 0 400108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4349
timestamp 1676037725
transform 1 0 401212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4361
timestamp 1676037725
transform 1 0 402316 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4367
timestamp 1676037725
transform 1 0 402868 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4369
timestamp 1676037725
transform 1 0 403052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4381
timestamp 1676037725
transform 1 0 404156 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4393
timestamp 1676037725
transform 1 0 405260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4405
timestamp 1676037725
transform 1 0 406364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4417
timestamp 1676037725
transform 1 0 407468 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4423
timestamp 1676037725
transform 1 0 408020 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4425
timestamp 1676037725
transform 1 0 408204 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4437
timestamp 1676037725
transform 1 0 409308 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4449
timestamp 1676037725
transform 1 0 410412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4461
timestamp 1676037725
transform 1 0 411516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4473
timestamp 1676037725
transform 1 0 412620 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4479
timestamp 1676037725
transform 1 0 413172 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4481
timestamp 1676037725
transform 1 0 413356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4493
timestamp 1676037725
transform 1 0 414460 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4505
timestamp 1676037725
transform 1 0 415564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4517
timestamp 1676037725
transform 1 0 416668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4529
timestamp 1676037725
transform 1 0 417772 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4535
timestamp 1676037725
transform 1 0 418324 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4537
timestamp 1676037725
transform 1 0 418508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4549
timestamp 1676037725
transform 1 0 419612 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4561
timestamp 1676037725
transform 1 0 420716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4573
timestamp 1676037725
transform 1 0 421820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4585
timestamp 1676037725
transform 1 0 422924 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4591
timestamp 1676037725
transform 1 0 423476 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4593
timestamp 1676037725
transform 1 0 423660 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4605
timestamp 1676037725
transform 1 0 424764 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4617
timestamp 1676037725
transform 1 0 425868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4629
timestamp 1676037725
transform 1 0 426972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4641
timestamp 1676037725
transform 1 0 428076 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4647
timestamp 1676037725
transform 1 0 428628 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4649
timestamp 1676037725
transform 1 0 428812 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4661
timestamp 1676037725
transform 1 0 429916 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4673
timestamp 1676037725
transform 1 0 431020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4685
timestamp 1676037725
transform 1 0 432124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4697
timestamp 1676037725
transform 1 0 433228 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4703
timestamp 1676037725
transform 1 0 433780 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4705
timestamp 1676037725
transform 1 0 433964 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4717
timestamp 1676037725
transform 1 0 435068 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4729
timestamp 1676037725
transform 1 0 436172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4741
timestamp 1676037725
transform 1 0 437276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4753
timestamp 1676037725
transform 1 0 438380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4759
timestamp 1676037725
transform 1 0 438932 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4761
timestamp 1676037725
transform 1 0 439116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4773
timestamp 1676037725
transform 1 0 440220 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4785
timestamp 1676037725
transform 1 0 441324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4797
timestamp 1676037725
transform 1 0 442428 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4809
timestamp 1676037725
transform 1 0 443532 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4815
timestamp 1676037725
transform 1 0 444084 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4817
timestamp 1676037725
transform 1 0 444268 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4829
timestamp 1676037725
transform 1 0 445372 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4841
timestamp 1676037725
transform 1 0 446476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4853
timestamp 1676037725
transform 1 0 447580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4865
timestamp 1676037725
transform 1 0 448684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4871
timestamp 1676037725
transform 1 0 449236 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4873
timestamp 1676037725
transform 1 0 449420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4885
timestamp 1676037725
transform 1 0 450524 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4897
timestamp 1676037725
transform 1 0 451628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4909
timestamp 1676037725
transform 1 0 452732 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4921
timestamp 1676037725
transform 1 0 453836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4927
timestamp 1676037725
transform 1 0 454388 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4929
timestamp 1676037725
transform 1 0 454572 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4941
timestamp 1676037725
transform 1 0 455676 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4953
timestamp 1676037725
transform 1 0 456780 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4965
timestamp 1676037725
transform 1 0 457884 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_4977
timestamp 1676037725
transform 1 0 458988 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_4983
timestamp 1676037725
transform 1 0 459540 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4985
timestamp 1676037725
transform 1 0 459724 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_4997
timestamp 1676037725
transform 1 0 460828 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5009
timestamp 1676037725
transform 1 0 461932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5021
timestamp 1676037725
transform 1 0 463036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5033
timestamp 1676037725
transform 1 0 464140 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5039
timestamp 1676037725
transform 1 0 464692 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5041
timestamp 1676037725
transform 1 0 464876 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5053
timestamp 1676037725
transform 1 0 465980 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5065
timestamp 1676037725
transform 1 0 467084 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5077
timestamp 1676037725
transform 1 0 468188 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5089
timestamp 1676037725
transform 1 0 469292 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5095
timestamp 1676037725
transform 1 0 469844 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5097
timestamp 1676037725
transform 1 0 470028 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5109
timestamp 1676037725
transform 1 0 471132 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5121
timestamp 1676037725
transform 1 0 472236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5133
timestamp 1676037725
transform 1 0 473340 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5145
timestamp 1676037725
transform 1 0 474444 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5151
timestamp 1676037725
transform 1 0 474996 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5153
timestamp 1676037725
transform 1 0 475180 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5165
timestamp 1676037725
transform 1 0 476284 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5177
timestamp 1676037725
transform 1 0 477388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5189
timestamp 1676037725
transform 1 0 478492 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5201
timestamp 1676037725
transform 1 0 479596 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5207
timestamp 1676037725
transform 1 0 480148 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5209
timestamp 1676037725
transform 1 0 480332 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5221
timestamp 1676037725
transform 1 0 481436 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5233
timestamp 1676037725
transform 1 0 482540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5245
timestamp 1676037725
transform 1 0 483644 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5257
timestamp 1676037725
transform 1 0 484748 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5263
timestamp 1676037725
transform 1 0 485300 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5265
timestamp 1676037725
transform 1 0 485484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5277
timestamp 1676037725
transform 1 0 486588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5289
timestamp 1676037725
transform 1 0 487692 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5301
timestamp 1676037725
transform 1 0 488796 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5313
timestamp 1676037725
transform 1 0 489900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5319
timestamp 1676037725
transform 1 0 490452 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5321
timestamp 1676037725
transform 1 0 490636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5333
timestamp 1676037725
transform 1 0 491740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5345
timestamp 1676037725
transform 1 0 492844 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5357
timestamp 1676037725
transform 1 0 493948 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5369
timestamp 1676037725
transform 1 0 495052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5375
timestamp 1676037725
transform 1 0 495604 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5377
timestamp 1676037725
transform 1 0 495788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5389
timestamp 1676037725
transform 1 0 496892 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5401
timestamp 1676037725
transform 1 0 497996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5413
timestamp 1676037725
transform 1 0 499100 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5425
timestamp 1676037725
transform 1 0 500204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5431
timestamp 1676037725
transform 1 0 500756 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5433
timestamp 1676037725
transform 1 0 500940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5445
timestamp 1676037725
transform 1 0 502044 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5457
timestamp 1676037725
transform 1 0 503148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5469
timestamp 1676037725
transform 1 0 504252 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5481
timestamp 1676037725
transform 1 0 505356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5487
timestamp 1676037725
transform 1 0 505908 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5489
timestamp 1676037725
transform 1 0 506092 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5501
timestamp 1676037725
transform 1 0 507196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5513
timestamp 1676037725
transform 1 0 508300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5525
timestamp 1676037725
transform 1 0 509404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5537
timestamp 1676037725
transform 1 0 510508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5543
timestamp 1676037725
transform 1 0 511060 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5545
timestamp 1676037725
transform 1 0 511244 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5557
timestamp 1676037725
transform 1 0 512348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5569
timestamp 1676037725
transform 1 0 513452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5581
timestamp 1676037725
transform 1 0 514556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5593
timestamp 1676037725
transform 1 0 515660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5599
timestamp 1676037725
transform 1 0 516212 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5601
timestamp 1676037725
transform 1 0 516396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5613
timestamp 1676037725
transform 1 0 517500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5625
timestamp 1676037725
transform 1 0 518604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5637
timestamp 1676037725
transform 1 0 519708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5649
timestamp 1676037725
transform 1 0 520812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5655
timestamp 1676037725
transform 1 0 521364 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5657
timestamp 1676037725
transform 1 0 521548 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5669
timestamp 1676037725
transform 1 0 522652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5681
timestamp 1676037725
transform 1 0 523756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5693
timestamp 1676037725
transform 1 0 524860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_5705
timestamp 1676037725
transform 1 0 525964 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5711
timestamp 1676037725
transform 1 0 526516 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_5713
timestamp 1676037725
transform 1 0 526700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_5725
timestamp 1676037725
transform 1 0 527804 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1676037725
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1676037725
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1676037725
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1676037725
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1676037725
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1676037725
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1676037725
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1676037725
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1676037725
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1676037725
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1676037725
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1676037725
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1676037725
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1676037725
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1676037725
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1676037725
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1676037725
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1676037725
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1676037725
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1676037725
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1676037725
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1676037725
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1676037725
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1676037725
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1676037725
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1676037725
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1676037725
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1676037725
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1676037725
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1676037725
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1676037725
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1676037725
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_813
timestamp 1676037725
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_825
timestamp 1676037725
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_837
timestamp 1676037725
transform 1 0 78108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_849
timestamp 1676037725
transform 1 0 79212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_861
timestamp 1676037725
transform 1 0 80316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_867
timestamp 1676037725
transform 1 0 80868 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_869
timestamp 1676037725
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_881
timestamp 1676037725
transform 1 0 82156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_893
timestamp 1676037725
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_905
timestamp 1676037725
transform 1 0 84364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1676037725
transform 1 0 85468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1676037725
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_925
timestamp 1676037725
transform 1 0 86204 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_937
timestamp 1676037725
transform 1 0 87308 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_949
timestamp 1676037725
transform 1 0 88412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_961
timestamp 1676037725
transform 1 0 89516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_973
timestamp 1676037725
transform 1 0 90620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_979
timestamp 1676037725
transform 1 0 91172 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_981
timestamp 1676037725
transform 1 0 91356 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_993
timestamp 1676037725
transform 1 0 92460 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1005
timestamp 1676037725
transform 1 0 93564 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1017
timestamp 1676037725
transform 1 0 94668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1029
timestamp 1676037725
transform 1 0 95772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1035
timestamp 1676037725
transform 1 0 96324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1037
timestamp 1676037725
transform 1 0 96508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1049
timestamp 1676037725
transform 1 0 97612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1061
timestamp 1676037725
transform 1 0 98716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1073
timestamp 1676037725
transform 1 0 99820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1085
timestamp 1676037725
transform 1 0 100924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1091
timestamp 1676037725
transform 1 0 101476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1093
timestamp 1676037725
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1105
timestamp 1676037725
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1117
timestamp 1676037725
transform 1 0 103868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1129
timestamp 1676037725
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1141
timestamp 1676037725
transform 1 0 106076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1147
timestamp 1676037725
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1149
timestamp 1676037725
transform 1 0 106812 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1161
timestamp 1676037725
transform 1 0 107916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1173
timestamp 1676037725
transform 1 0 109020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1185
timestamp 1676037725
transform 1 0 110124 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1197
timestamp 1676037725
transform 1 0 111228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1203
timestamp 1676037725
transform 1 0 111780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1205
timestamp 1676037725
transform 1 0 111964 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1217
timestamp 1676037725
transform 1 0 113068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1229
timestamp 1676037725
transform 1 0 114172 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1241
timestamp 1676037725
transform 1 0 115276 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1253
timestamp 1676037725
transform 1 0 116380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1259
timestamp 1676037725
transform 1 0 116932 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1261
timestamp 1676037725
transform 1 0 117116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1273
timestamp 1676037725
transform 1 0 118220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1285
timestamp 1676037725
transform 1 0 119324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1297
timestamp 1676037725
transform 1 0 120428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1309
timestamp 1676037725
transform 1 0 121532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1315
timestamp 1676037725
transform 1 0 122084 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1317
timestamp 1676037725
transform 1 0 122268 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1329
timestamp 1676037725
transform 1 0 123372 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1341
timestamp 1676037725
transform 1 0 124476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1353
timestamp 1676037725
transform 1 0 125580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1365
timestamp 1676037725
transform 1 0 126684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1371
timestamp 1676037725
transform 1 0 127236 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1373
timestamp 1676037725
transform 1 0 127420 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1385
timestamp 1676037725
transform 1 0 128524 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1397
timestamp 1676037725
transform 1 0 129628 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1409
timestamp 1676037725
transform 1 0 130732 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1421
timestamp 1676037725
transform 1 0 131836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1427
timestamp 1676037725
transform 1 0 132388 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1429
timestamp 1676037725
transform 1 0 132572 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1441
timestamp 1676037725
transform 1 0 133676 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1453
timestamp 1676037725
transform 1 0 134780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1465
timestamp 1676037725
transform 1 0 135884 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1477
timestamp 1676037725
transform 1 0 136988 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1483
timestamp 1676037725
transform 1 0 137540 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1485
timestamp 1676037725
transform 1 0 137724 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1497
timestamp 1676037725
transform 1 0 138828 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1509
timestamp 1676037725
transform 1 0 139932 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1521
timestamp 1676037725
transform 1 0 141036 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1533
timestamp 1676037725
transform 1 0 142140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1539
timestamp 1676037725
transform 1 0 142692 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1541
timestamp 1676037725
transform 1 0 142876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1553
timestamp 1676037725
transform 1 0 143980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1565
timestamp 1676037725
transform 1 0 145084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1577
timestamp 1676037725
transform 1 0 146188 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1589
timestamp 1676037725
transform 1 0 147292 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1595
timestamp 1676037725
transform 1 0 147844 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1597
timestamp 1676037725
transform 1 0 148028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1609
timestamp 1676037725
transform 1 0 149132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1621
timestamp 1676037725
transform 1 0 150236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1633
timestamp 1676037725
transform 1 0 151340 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1650
timestamp 1676037725
transform 1 0 152904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1653
timestamp 1676037725
transform 1 0 153180 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1657
timestamp 1676037725
transform 1 0 153548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1669
timestamp 1676037725
transform 1 0 154652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1681
timestamp 1676037725
transform 1 0 155756 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1693
timestamp 1676037725
transform 1 0 156860 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1705
timestamp 1676037725
transform 1 0 157964 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1709
timestamp 1676037725
transform 1 0 158332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1721
timestamp 1676037725
transform 1 0 159436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1734
timestamp 1676037725
transform 1 0 160632 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1740
timestamp 1676037725
transform 1 0 161184 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1752
timestamp 1676037725
transform 1 0 162288 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1765
timestamp 1676037725
transform 1 0 163484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1777
timestamp 1676037725
transform 1 0 164588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1789
timestamp 1676037725
transform 1 0 165692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1801
timestamp 1676037725
transform 1 0 166796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1807
timestamp 1676037725
transform 1 0 167348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1817
timestamp 1676037725
transform 1 0 168268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1821
timestamp 1676037725
transform 1 0 168636 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1825
timestamp 1676037725
transform 1 0 169004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1837
timestamp 1676037725
transform 1 0 170108 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1849
timestamp 1676037725
transform 1 0 171212 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1864
timestamp 1676037725
transform 1 0 172592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1870
timestamp 1676037725
transform 1 0 173144 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1877
timestamp 1676037725
transform 1 0 173788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1889
timestamp 1676037725
transform 1 0 174892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1899
timestamp 1676037725
transform 1 0 175812 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1905
timestamp 1676037725
transform 1 0 176364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1917
timestamp 1676037725
transform 1 0 177468 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1929
timestamp 1676037725
transform 1 0 178572 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1933
timestamp 1676037725
transform 1 0 178940 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1946
timestamp 1676037725
transform 1 0 180136 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1952
timestamp 1676037725
transform 1 0 180688 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1964
timestamp 1676037725
transform 1 0 181792 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1976
timestamp 1676037725
transform 1 0 182896 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1989
timestamp 1676037725
transform 1 0 184092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2001
timestamp 1676037725
transform 1 0 185196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2013
timestamp 1676037725
transform 1 0 186300 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2019
timestamp 1676037725
transform 1 0 186852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_2029
timestamp 1676037725
transform 1 0 187772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_2035
timestamp 1676037725
transform 1 0 188324 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2043
timestamp 1676037725
transform 1 0 189060 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2045
timestamp 1676037725
transform 1 0 189244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2057
timestamp 1676037725
transform 1 0 190348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2069
timestamp 1676037725
transform 1 0 191452 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2081
timestamp 1676037725
transform 1 0 192556 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2093
timestamp 1676037725
transform 1 0 193660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2099
timestamp 1676037725
transform 1 0 194212 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2101
timestamp 1676037725
transform 1 0 194396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2113
timestamp 1676037725
transform 1 0 195500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2125
timestamp 1676037725
transform 1 0 196604 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2137
timestamp 1676037725
transform 1 0 197708 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2149
timestamp 1676037725
transform 1 0 198812 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2155
timestamp 1676037725
transform 1 0 199364 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2157
timestamp 1676037725
transform 1 0 199548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2169
timestamp 1676037725
transform 1 0 200652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2181
timestamp 1676037725
transform 1 0 201756 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2193
timestamp 1676037725
transform 1 0 202860 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2205
timestamp 1676037725
transform 1 0 203964 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2211
timestamp 1676037725
transform 1 0 204516 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2213
timestamp 1676037725
transform 1 0 204700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2225
timestamp 1676037725
transform 1 0 205804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2237
timestamp 1676037725
transform 1 0 206908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2249
timestamp 1676037725
transform 1 0 208012 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2261
timestamp 1676037725
transform 1 0 209116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2267
timestamp 1676037725
transform 1 0 209668 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2269
timestamp 1676037725
transform 1 0 209852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2281
timestamp 1676037725
transform 1 0 210956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2293
timestamp 1676037725
transform 1 0 212060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2305
timestamp 1676037725
transform 1 0 213164 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2317
timestamp 1676037725
transform 1 0 214268 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2323
timestamp 1676037725
transform 1 0 214820 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2325
timestamp 1676037725
transform 1 0 215004 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2337
timestamp 1676037725
transform 1 0 216108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2349
timestamp 1676037725
transform 1 0 217212 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2361
timestamp 1676037725
transform 1 0 218316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2373
timestamp 1676037725
transform 1 0 219420 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2379
timestamp 1676037725
transform 1 0 219972 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2381
timestamp 1676037725
transform 1 0 220156 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2393
timestamp 1676037725
transform 1 0 221260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2405
timestamp 1676037725
transform 1 0 222364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2417
timestamp 1676037725
transform 1 0 223468 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2429
timestamp 1676037725
transform 1 0 224572 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2435
timestamp 1676037725
transform 1 0 225124 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2437
timestamp 1676037725
transform 1 0 225308 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2449
timestamp 1676037725
transform 1 0 226412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2461
timestamp 1676037725
transform 1 0 227516 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2473
timestamp 1676037725
transform 1 0 228620 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2485
timestamp 1676037725
transform 1 0 229724 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2491
timestamp 1676037725
transform 1 0 230276 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2493
timestamp 1676037725
transform 1 0 230460 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2505
timestamp 1676037725
transform 1 0 231564 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2517
timestamp 1676037725
transform 1 0 232668 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2529
timestamp 1676037725
transform 1 0 233772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2541
timestamp 1676037725
transform 1 0 234876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2547
timestamp 1676037725
transform 1 0 235428 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2549
timestamp 1676037725
transform 1 0 235612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2561
timestamp 1676037725
transform 1 0 236716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2573
timestamp 1676037725
transform 1 0 237820 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2585
timestamp 1676037725
transform 1 0 238924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_2599
timestamp 1676037725
transform 1 0 240212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2603
timestamp 1676037725
transform 1 0 240580 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2605
timestamp 1676037725
transform 1 0 240764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2617
timestamp 1676037725
transform 1 0 241868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2629
timestamp 1676037725
transform 1 0 242972 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2641
timestamp 1676037725
transform 1 0 244076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2653
timestamp 1676037725
transform 1 0 245180 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2659
timestamp 1676037725
transform 1 0 245732 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2661
timestamp 1676037725
transform 1 0 245916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2673
timestamp 1676037725
transform 1 0 247020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2685
timestamp 1676037725
transform 1 0 248124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2697
timestamp 1676037725
transform 1 0 249228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2709
timestamp 1676037725
transform 1 0 250332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2715
timestamp 1676037725
transform 1 0 250884 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2717
timestamp 1676037725
transform 1 0 251068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2729
timestamp 1676037725
transform 1 0 252172 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2741
timestamp 1676037725
transform 1 0 253276 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2753
timestamp 1676037725
transform 1 0 254380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2765
timestamp 1676037725
transform 1 0 255484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2771
timestamp 1676037725
transform 1 0 256036 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2773
timestamp 1676037725
transform 1 0 256220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2785
timestamp 1676037725
transform 1 0 257324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2797
timestamp 1676037725
transform 1 0 258428 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2809
timestamp 1676037725
transform 1 0 259532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2821
timestamp 1676037725
transform 1 0 260636 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2827
timestamp 1676037725
transform 1 0 261188 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2829
timestamp 1676037725
transform 1 0 261372 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2841
timestamp 1676037725
transform 1 0 262476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2853
timestamp 1676037725
transform 1 0 263580 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2865
timestamp 1676037725
transform 1 0 264684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2877
timestamp 1676037725
transform 1 0 265788 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2883
timestamp 1676037725
transform 1 0 266340 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2885
timestamp 1676037725
transform 1 0 266524 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2897
timestamp 1676037725
transform 1 0 267628 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2909
timestamp 1676037725
transform 1 0 268732 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2921
timestamp 1676037725
transform 1 0 269836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2933
timestamp 1676037725
transform 1 0 270940 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2939
timestamp 1676037725
transform 1 0 271492 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2941
timestamp 1676037725
transform 1 0 271676 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2953
timestamp 1676037725
transform 1 0 272780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2965
timestamp 1676037725
transform 1 0 273884 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2977
timestamp 1676037725
transform 1 0 274988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_2989
timestamp 1676037725
transform 1 0 276092 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_2995
timestamp 1676037725
transform 1 0 276644 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_2997
timestamp 1676037725
transform 1 0 276828 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3009
timestamp 1676037725
transform 1 0 277932 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3021
timestamp 1676037725
transform 1 0 279036 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3033
timestamp 1676037725
transform 1 0 280140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3045
timestamp 1676037725
transform 1 0 281244 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3051
timestamp 1676037725
transform 1 0 281796 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3053
timestamp 1676037725
transform 1 0 281980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3065
timestamp 1676037725
transform 1 0 283084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3077
timestamp 1676037725
transform 1 0 284188 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3089
timestamp 1676037725
transform 1 0 285292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3101
timestamp 1676037725
transform 1 0 286396 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3107
timestamp 1676037725
transform 1 0 286948 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3109
timestamp 1676037725
transform 1 0 287132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3121
timestamp 1676037725
transform 1 0 288236 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3133
timestamp 1676037725
transform 1 0 289340 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3145
timestamp 1676037725
transform 1 0 290444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3157
timestamp 1676037725
transform 1 0 291548 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3163
timestamp 1676037725
transform 1 0 292100 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3165
timestamp 1676037725
transform 1 0 292284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3177
timestamp 1676037725
transform 1 0 293388 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3189
timestamp 1676037725
transform 1 0 294492 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3201
timestamp 1676037725
transform 1 0 295596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3213
timestamp 1676037725
transform 1 0 296700 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3219
timestamp 1676037725
transform 1 0 297252 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3221
timestamp 1676037725
transform 1 0 297436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3233
timestamp 1676037725
transform 1 0 298540 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3245
timestamp 1676037725
transform 1 0 299644 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3257
timestamp 1676037725
transform 1 0 300748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3269
timestamp 1676037725
transform 1 0 301852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3275
timestamp 1676037725
transform 1 0 302404 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3277
timestamp 1676037725
transform 1 0 302588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3289
timestamp 1676037725
transform 1 0 303692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3301
timestamp 1676037725
transform 1 0 304796 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3313
timestamp 1676037725
transform 1 0 305900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3325
timestamp 1676037725
transform 1 0 307004 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3331
timestamp 1676037725
transform 1 0 307556 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3333
timestamp 1676037725
transform 1 0 307740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3345
timestamp 1676037725
transform 1 0 308844 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3357
timestamp 1676037725
transform 1 0 309948 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3369
timestamp 1676037725
transform 1 0 311052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3381
timestamp 1676037725
transform 1 0 312156 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3387
timestamp 1676037725
transform 1 0 312708 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3389
timestamp 1676037725
transform 1 0 312892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3401
timestamp 1676037725
transform 1 0 313996 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3413
timestamp 1676037725
transform 1 0 315100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3425
timestamp 1676037725
transform 1 0 316204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3437
timestamp 1676037725
transform 1 0 317308 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3443
timestamp 1676037725
transform 1 0 317860 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3445
timestamp 1676037725
transform 1 0 318044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3457
timestamp 1676037725
transform 1 0 319148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3469
timestamp 1676037725
transform 1 0 320252 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3477
timestamp 1676037725
transform 1 0 320988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3488
timestamp 1676037725
transform 1 0 322000 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3494
timestamp 1676037725
transform 1 0 322552 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3501
timestamp 1676037725
transform 1 0 323196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3513
timestamp 1676037725
transform 1 0 324300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3525
timestamp 1676037725
transform 1 0 325404 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3533
timestamp 1676037725
transform 1 0 326140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3543
timestamp 1676037725
transform 1 0 327060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3549
timestamp 1676037725
transform 1 0 327612 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3555
timestamp 1676037725
transform 1 0 328164 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3557
timestamp 1676037725
transform 1 0 328348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3569
timestamp 1676037725
transform 1 0 329452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3581
timestamp 1676037725
transform 1 0 330556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3587
timestamp 1676037725
transform 1 0 331108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3597
timestamp 1676037725
transform 1 0 332028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3603
timestamp 1676037725
transform 1 0 332580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3611
timestamp 1676037725
transform 1 0 333316 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3613
timestamp 1676037725
transform 1 0 333500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3625
timestamp 1676037725
transform 1 0 334604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3637
timestamp 1676037725
transform 1 0 335708 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3641
timestamp 1676037725
transform 1 0 336076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3651
timestamp 1676037725
transform 1 0 336996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3657
timestamp 1676037725
transform 1 0 337548 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3665
timestamp 1676037725
transform 1 0 338284 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3669
timestamp 1676037725
transform 1 0 338652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3681
timestamp 1676037725
transform 1 0 339756 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3693
timestamp 1676037725
transform 1 0 340860 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3705
timestamp 1676037725
transform 1 0 341964 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3717
timestamp 1676037725
transform 1 0 343068 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3723
timestamp 1676037725
transform 1 0 343620 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3725
timestamp 1676037725
transform 1 0 343804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3737
timestamp 1676037725
transform 1 0 344908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3749
timestamp 1676037725
transform 1 0 346012 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3761
timestamp 1676037725
transform 1 0 347116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3773
timestamp 1676037725
transform 1 0 348220 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3779
timestamp 1676037725
transform 1 0 348772 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3781
timestamp 1676037725
transform 1 0 348956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3793
timestamp 1676037725
transform 1 0 350060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3805
timestamp 1676037725
transform 1 0 351164 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3817
timestamp 1676037725
transform 1 0 352268 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3829
timestamp 1676037725
transform 1 0 353372 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3835
timestamp 1676037725
transform 1 0 353924 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3837
timestamp 1676037725
transform 1 0 354108 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3849
timestamp 1676037725
transform 1 0 355212 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3861
timestamp 1676037725
transform 1 0 356316 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3873
timestamp 1676037725
transform 1 0 357420 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3885
timestamp 1676037725
transform 1 0 358524 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3891
timestamp 1676037725
transform 1 0 359076 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3893
timestamp 1676037725
transform 1 0 359260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3905
timestamp 1676037725
transform 1 0 360364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3917
timestamp 1676037725
transform 1 0 361468 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3929
timestamp 1676037725
transform 1 0 362572 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3941
timestamp 1676037725
transform 1 0 363676 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3947
timestamp 1676037725
transform 1 0 364228 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3949
timestamp 1676037725
transform 1 0 364412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3961
timestamp 1676037725
transform 1 0 365516 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3973
timestamp 1676037725
transform 1 0 366620 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3985
timestamp 1676037725
transform 1 0 367724 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3997
timestamp 1676037725
transform 1 0 368828 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4003
timestamp 1676037725
transform 1 0 369380 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4005
timestamp 1676037725
transform 1 0 369564 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_4017
timestamp 1676037725
transform 1 0 370668 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4027
timestamp 1676037725
transform 1 0 371588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4039
timestamp 1676037725
transform 1 0 372692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_4051
timestamp 1676037725
transform 1 0 373796 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4059
timestamp 1676037725
transform 1 0 374532 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4061
timestamp 1676037725
transform 1 0 374716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4073
timestamp 1676037725
transform 1 0 375820 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4085
timestamp 1676037725
transform 1 0 376924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4097
timestamp 1676037725
transform 1 0 378028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4109
timestamp 1676037725
transform 1 0 379132 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4115
timestamp 1676037725
transform 1 0 379684 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4117
timestamp 1676037725
transform 1 0 379868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4129
timestamp 1676037725
transform 1 0 380972 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4141
timestamp 1676037725
transform 1 0 382076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4153
timestamp 1676037725
transform 1 0 383180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4165
timestamp 1676037725
transform 1 0 384284 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4171
timestamp 1676037725
transform 1 0 384836 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4173
timestamp 1676037725
transform 1 0 385020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4185
timestamp 1676037725
transform 1 0 386124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4197
timestamp 1676037725
transform 1 0 387228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4209
timestamp 1676037725
transform 1 0 388332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4221
timestamp 1676037725
transform 1 0 389436 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4227
timestamp 1676037725
transform 1 0 389988 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4229
timestamp 1676037725
transform 1 0 390172 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4241
timestamp 1676037725
transform 1 0 391276 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4253
timestamp 1676037725
transform 1 0 392380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4265
timestamp 1676037725
transform 1 0 393484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4277
timestamp 1676037725
transform 1 0 394588 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4283
timestamp 1676037725
transform 1 0 395140 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4285
timestamp 1676037725
transform 1 0 395324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4297
timestamp 1676037725
transform 1 0 396428 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4309
timestamp 1676037725
transform 1 0 397532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4321
timestamp 1676037725
transform 1 0 398636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4333
timestamp 1676037725
transform 1 0 399740 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4339
timestamp 1676037725
transform 1 0 400292 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4341
timestamp 1676037725
transform 1 0 400476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4353
timestamp 1676037725
transform 1 0 401580 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4365
timestamp 1676037725
transform 1 0 402684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4377
timestamp 1676037725
transform 1 0 403788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4389
timestamp 1676037725
transform 1 0 404892 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4395
timestamp 1676037725
transform 1 0 405444 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4397
timestamp 1676037725
transform 1 0 405628 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4409
timestamp 1676037725
transform 1 0 406732 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4421
timestamp 1676037725
transform 1 0 407836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4433
timestamp 1676037725
transform 1 0 408940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4445
timestamp 1676037725
transform 1 0 410044 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4451
timestamp 1676037725
transform 1 0 410596 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4453
timestamp 1676037725
transform 1 0 410780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4465
timestamp 1676037725
transform 1 0 411884 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4477
timestamp 1676037725
transform 1 0 412988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4489
timestamp 1676037725
transform 1 0 414092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4501
timestamp 1676037725
transform 1 0 415196 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4507
timestamp 1676037725
transform 1 0 415748 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4509
timestamp 1676037725
transform 1 0 415932 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4521
timestamp 1676037725
transform 1 0 417036 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4533
timestamp 1676037725
transform 1 0 418140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4545
timestamp 1676037725
transform 1 0 419244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4557
timestamp 1676037725
transform 1 0 420348 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4563
timestamp 1676037725
transform 1 0 420900 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4565
timestamp 1676037725
transform 1 0 421084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4577
timestamp 1676037725
transform 1 0 422188 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4589
timestamp 1676037725
transform 1 0 423292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4601
timestamp 1676037725
transform 1 0 424396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4613
timestamp 1676037725
transform 1 0 425500 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4619
timestamp 1676037725
transform 1 0 426052 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4621
timestamp 1676037725
transform 1 0 426236 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4633
timestamp 1676037725
transform 1 0 427340 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4645
timestamp 1676037725
transform 1 0 428444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4657
timestamp 1676037725
transform 1 0 429548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4669
timestamp 1676037725
transform 1 0 430652 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4675
timestamp 1676037725
transform 1 0 431204 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4677
timestamp 1676037725
transform 1 0 431388 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4689
timestamp 1676037725
transform 1 0 432492 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4701
timestamp 1676037725
transform 1 0 433596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4713
timestamp 1676037725
transform 1 0 434700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4725
timestamp 1676037725
transform 1 0 435804 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4731
timestamp 1676037725
transform 1 0 436356 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4733
timestamp 1676037725
transform 1 0 436540 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4745
timestamp 1676037725
transform 1 0 437644 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4757
timestamp 1676037725
transform 1 0 438748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4769
timestamp 1676037725
transform 1 0 439852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4781
timestamp 1676037725
transform 1 0 440956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4787
timestamp 1676037725
transform 1 0 441508 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4789
timestamp 1676037725
transform 1 0 441692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4801
timestamp 1676037725
transform 1 0 442796 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4813
timestamp 1676037725
transform 1 0 443900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4825
timestamp 1676037725
transform 1 0 445004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4837
timestamp 1676037725
transform 1 0 446108 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4843
timestamp 1676037725
transform 1 0 446660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4845
timestamp 1676037725
transform 1 0 446844 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4857
timestamp 1676037725
transform 1 0 447948 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4869
timestamp 1676037725
transform 1 0 449052 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4881
timestamp 1676037725
transform 1 0 450156 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4893
timestamp 1676037725
transform 1 0 451260 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4899
timestamp 1676037725
transform 1 0 451812 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4901
timestamp 1676037725
transform 1 0 451996 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4913
timestamp 1676037725
transform 1 0 453100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4925
timestamp 1676037725
transform 1 0 454204 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4937
timestamp 1676037725
transform 1 0 455308 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_4949
timestamp 1676037725
transform 1 0 456412 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_4955
timestamp 1676037725
transform 1 0 456964 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4957
timestamp 1676037725
transform 1 0 457148 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4969
timestamp 1676037725
transform 1 0 458252 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4981
timestamp 1676037725
transform 1 0 459356 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_4993
timestamp 1676037725
transform 1 0 460460 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5005
timestamp 1676037725
transform 1 0 461564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5011
timestamp 1676037725
transform 1 0 462116 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5013
timestamp 1676037725
transform 1 0 462300 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5025
timestamp 1676037725
transform 1 0 463404 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5037
timestamp 1676037725
transform 1 0 464508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5049
timestamp 1676037725
transform 1 0 465612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5061
timestamp 1676037725
transform 1 0 466716 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5067
timestamp 1676037725
transform 1 0 467268 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5069
timestamp 1676037725
transform 1 0 467452 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5081
timestamp 1676037725
transform 1 0 468556 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5093
timestamp 1676037725
transform 1 0 469660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5105
timestamp 1676037725
transform 1 0 470764 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5117
timestamp 1676037725
transform 1 0 471868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5123
timestamp 1676037725
transform 1 0 472420 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5125
timestamp 1676037725
transform 1 0 472604 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5137
timestamp 1676037725
transform 1 0 473708 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5149
timestamp 1676037725
transform 1 0 474812 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5161
timestamp 1676037725
transform 1 0 475916 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5173
timestamp 1676037725
transform 1 0 477020 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5179
timestamp 1676037725
transform 1 0 477572 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5181
timestamp 1676037725
transform 1 0 477756 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5193
timestamp 1676037725
transform 1 0 478860 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5205
timestamp 1676037725
transform 1 0 479964 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5217
timestamp 1676037725
transform 1 0 481068 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5229
timestamp 1676037725
transform 1 0 482172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5235
timestamp 1676037725
transform 1 0 482724 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5237
timestamp 1676037725
transform 1 0 482908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5249
timestamp 1676037725
transform 1 0 484012 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5261
timestamp 1676037725
transform 1 0 485116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5273
timestamp 1676037725
transform 1 0 486220 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5285
timestamp 1676037725
transform 1 0 487324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5291
timestamp 1676037725
transform 1 0 487876 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5293
timestamp 1676037725
transform 1 0 488060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5305
timestamp 1676037725
transform 1 0 489164 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5317
timestamp 1676037725
transform 1 0 490268 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5329
timestamp 1676037725
transform 1 0 491372 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5341
timestamp 1676037725
transform 1 0 492476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5347
timestamp 1676037725
transform 1 0 493028 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5349
timestamp 1676037725
transform 1 0 493212 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5361
timestamp 1676037725
transform 1 0 494316 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5373
timestamp 1676037725
transform 1 0 495420 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5385
timestamp 1676037725
transform 1 0 496524 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5397
timestamp 1676037725
transform 1 0 497628 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5403
timestamp 1676037725
transform 1 0 498180 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5405
timestamp 1676037725
transform 1 0 498364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5417
timestamp 1676037725
transform 1 0 499468 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5429
timestamp 1676037725
transform 1 0 500572 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5441
timestamp 1676037725
transform 1 0 501676 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5453
timestamp 1676037725
transform 1 0 502780 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5459
timestamp 1676037725
transform 1 0 503332 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5461
timestamp 1676037725
transform 1 0 503516 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5473
timestamp 1676037725
transform 1 0 504620 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5485
timestamp 1676037725
transform 1 0 505724 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5497
timestamp 1676037725
transform 1 0 506828 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5509
timestamp 1676037725
transform 1 0 507932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5515
timestamp 1676037725
transform 1 0 508484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5517
timestamp 1676037725
transform 1 0 508668 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5529
timestamp 1676037725
transform 1 0 509772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5541
timestamp 1676037725
transform 1 0 510876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5553
timestamp 1676037725
transform 1 0 511980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5565
timestamp 1676037725
transform 1 0 513084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5571
timestamp 1676037725
transform 1 0 513636 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5573
timestamp 1676037725
transform 1 0 513820 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5585
timestamp 1676037725
transform 1 0 514924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5597
timestamp 1676037725
transform 1 0 516028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5609
timestamp 1676037725
transform 1 0 517132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5621
timestamp 1676037725
transform 1 0 518236 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5627
timestamp 1676037725
transform 1 0 518788 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5629
timestamp 1676037725
transform 1 0 518972 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5641
timestamp 1676037725
transform 1 0 520076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5653
timestamp 1676037725
transform 1 0 521180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5665
timestamp 1676037725
transform 1 0 522284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_5677
timestamp 1676037725
transform 1 0 523388 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_5683
timestamp 1676037725
transform 1 0 523940 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5685
timestamp 1676037725
transform 1 0 524124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5697
timestamp 1676037725
transform 1 0 525228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5709
timestamp 1676037725
transform 1 0 526332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5721
timestamp 1676037725
transform 1 0 527436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_29
timestamp 1676037725
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_41
timestamp 1676037725
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1676037725
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_85
timestamp 1676037725
transform 1 0 8924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_97
timestamp 1676037725
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_141
timestamp 1676037725
transform 1 0 14076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_153
timestamp 1676037725
transform 1 0 15180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_197
timestamp 1676037725
transform 1 0 19228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_209
timestamp 1676037725
transform 1 0 20332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1676037725
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_253
timestamp 1676037725
transform 1 0 24380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_265
timestamp 1676037725
transform 1 0 25484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1676037725
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_305
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_309
timestamp 1676037725
transform 1 0 29532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_321
timestamp 1676037725
transform 1 0 30636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_333
timestamp 1676037725
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_365
timestamp 1676037725
transform 1 0 34684 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_377
timestamp 1676037725
transform 1 0 35788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_389
timestamp 1676037725
transform 1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_421
timestamp 1676037725
transform 1 0 39836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_433
timestamp 1676037725
transform 1 0 40940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 1676037725
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_477
timestamp 1676037725
transform 1 0 44988 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_489
timestamp 1676037725
transform 1 0 46092 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_501
timestamp 1676037725
transform 1 0 47196 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_529
timestamp 1676037725
transform 1 0 49772 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_533
timestamp 1676037725
transform 1 0 50140 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_545
timestamp 1676037725
transform 1 0 51244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_557
timestamp 1676037725
transform 1 0 52348 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1676037725
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1676037725
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_585
timestamp 1676037725
transform 1 0 54924 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_589
timestamp 1676037725
transform 1 0 55292 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_601
timestamp 1676037725
transform 1 0 56396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_613
timestamp 1676037725
transform 1 0 57500 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1676037725
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1676037725
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_641
timestamp 1676037725
transform 1 0 60076 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_645
timestamp 1676037725
transform 1 0 60444 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_657
timestamp 1676037725
transform 1 0 61548 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_669
timestamp 1676037725
transform 1 0 62652 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1676037725
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1676037725
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_697
timestamp 1676037725
transform 1 0 65228 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_701
timestamp 1676037725
transform 1 0 65596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_713
timestamp 1676037725
transform 1 0 66700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_725
timestamp 1676037725
transform 1 0 67804 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1676037725
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1676037725
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_753
timestamp 1676037725
transform 1 0 70380 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_757
timestamp 1676037725
transform 1 0 70748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_769
timestamp 1676037725
transform 1 0 71852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_781
timestamp 1676037725
transform 1 0 72956 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1676037725
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1676037725
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_809
timestamp 1676037725
transform 1 0 75532 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_813
timestamp 1676037725
transform 1 0 75900 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_825
timestamp 1676037725
transform 1 0 77004 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_837
timestamp 1676037725
transform 1 0 78108 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_841
timestamp 1676037725
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_853
timestamp 1676037725
transform 1 0 79580 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_865
timestamp 1676037725
transform 1 0 80684 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_869
timestamp 1676037725
transform 1 0 81052 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_881
timestamp 1676037725
transform 1 0 82156 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_893
timestamp 1676037725
transform 1 0 83260 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_897
timestamp 1676037725
transform 1 0 83628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_909
timestamp 1676037725
transform 1 0 84732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_921
timestamp 1676037725
transform 1 0 85836 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_925
timestamp 1676037725
transform 1 0 86204 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_937
timestamp 1676037725
transform 1 0 87308 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_949
timestamp 1676037725
transform 1 0 88412 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_953
timestamp 1676037725
transform 1 0 88780 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_965
timestamp 1676037725
transform 1 0 89884 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_977
timestamp 1676037725
transform 1 0 90988 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_981
timestamp 1676037725
transform 1 0 91356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_993
timestamp 1676037725
transform 1 0 92460 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1005
timestamp 1676037725
transform 1 0 93564 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1009
timestamp 1676037725
transform 1 0 93932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1021
timestamp 1676037725
transform 1 0 95036 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1033
timestamp 1676037725
transform 1 0 96140 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1037
timestamp 1676037725
transform 1 0 96508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1049
timestamp 1676037725
transform 1 0 97612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1061
timestamp 1676037725
transform 1 0 98716 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1065
timestamp 1676037725
transform 1 0 99084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1077
timestamp 1676037725
transform 1 0 100188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1089
timestamp 1676037725
transform 1 0 101292 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1093
timestamp 1676037725
transform 1 0 101660 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1105
timestamp 1676037725
transform 1 0 102764 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1117
timestamp 1676037725
transform 1 0 103868 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1121
timestamp 1676037725
transform 1 0 104236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1133
timestamp 1676037725
transform 1 0 105340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1145
timestamp 1676037725
transform 1 0 106444 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1149
timestamp 1676037725
transform 1 0 106812 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1161
timestamp 1676037725
transform 1 0 107916 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1173
timestamp 1676037725
transform 1 0 109020 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1177
timestamp 1676037725
transform 1 0 109388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1189
timestamp 1676037725
transform 1 0 110492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1201
timestamp 1676037725
transform 1 0 111596 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1205
timestamp 1676037725
transform 1 0 111964 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1217
timestamp 1676037725
transform 1 0 113068 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1229
timestamp 1676037725
transform 1 0 114172 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1233
timestamp 1676037725
transform 1 0 114540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1245
timestamp 1676037725
transform 1 0 115644 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1257
timestamp 1676037725
transform 1 0 116748 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1261
timestamp 1676037725
transform 1 0 117116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1273
timestamp 1676037725
transform 1 0 118220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1285
timestamp 1676037725
transform 1 0 119324 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1289
timestamp 1676037725
transform 1 0 119692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1301
timestamp 1676037725
transform 1 0 120796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1313
timestamp 1676037725
transform 1 0 121900 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1317
timestamp 1676037725
transform 1 0 122268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1329
timestamp 1676037725
transform 1 0 123372 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1341
timestamp 1676037725
transform 1 0 124476 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1345
timestamp 1676037725
transform 1 0 124844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1357
timestamp 1676037725
transform 1 0 125948 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1369
timestamp 1676037725
transform 1 0 127052 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1373
timestamp 1676037725
transform 1 0 127420 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1385
timestamp 1676037725
transform 1 0 128524 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1397
timestamp 1676037725
transform 1 0 129628 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1401
timestamp 1676037725
transform 1 0 129996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1413
timestamp 1676037725
transform 1 0 131100 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1425
timestamp 1676037725
transform 1 0 132204 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1429
timestamp 1676037725
transform 1 0 132572 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1441
timestamp 1676037725
transform 1 0 133676 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1453
timestamp 1676037725
transform 1 0 134780 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1457
timestamp 1676037725
transform 1 0 135148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1469
timestamp 1676037725
transform 1 0 136252 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1481
timestamp 1676037725
transform 1 0 137356 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1485
timestamp 1676037725
transform 1 0 137724 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1497
timestamp 1676037725
transform 1 0 138828 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1509
timestamp 1676037725
transform 1 0 139932 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1513
timestamp 1676037725
transform 1 0 140300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1525
timestamp 1676037725
transform 1 0 141404 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1537
timestamp 1676037725
transform 1 0 142508 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1541
timestamp 1676037725
transform 1 0 142876 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1553
timestamp 1676037725
transform 1 0 143980 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1565
timestamp 1676037725
transform 1 0 145084 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1569
timestamp 1676037725
transform 1 0 145452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1581
timestamp 1676037725
transform 1 0 146556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1593
timestamp 1676037725
transform 1 0 147660 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1597
timestamp 1676037725
transform 1 0 148028 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1609
timestamp 1676037725
transform 1 0 149132 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1621
timestamp 1676037725
transform 1 0 150236 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1625
timestamp 1676037725
transform 1 0 150604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1637
timestamp 1676037725
transform 1 0 151708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1649
timestamp 1676037725
transform 1 0 152812 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1653
timestamp 1676037725
transform 1 0 153180 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1665
timestamp 1676037725
transform 1 0 154284 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1677
timestamp 1676037725
transform 1 0 155388 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1681
timestamp 1676037725
transform 1 0 155756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1693
timestamp 1676037725
transform 1 0 156860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1705
timestamp 1676037725
transform 1 0 157964 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1709
timestamp 1676037725
transform 1 0 158332 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1721
timestamp 1676037725
transform 1 0 159436 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1733
timestamp 1676037725
transform 1 0 160540 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1737
timestamp 1676037725
transform 1 0 160908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1749
timestamp 1676037725
transform 1 0 162012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1761
timestamp 1676037725
transform 1 0 163116 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1765
timestamp 1676037725
transform 1 0 163484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1777
timestamp 1676037725
transform 1 0 164588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1789
timestamp 1676037725
transform 1 0 165692 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1793
timestamp 1676037725
transform 1 0 166060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1805
timestamp 1676037725
transform 1 0 167164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1817
timestamp 1676037725
transform 1 0 168268 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1821
timestamp 1676037725
transform 1 0 168636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1833
timestamp 1676037725
transform 1 0 169740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1845
timestamp 1676037725
transform 1 0 170844 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1849
timestamp 1676037725
transform 1 0 171212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1861
timestamp 1676037725
transform 1 0 172316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1873
timestamp 1676037725
transform 1 0 173420 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1877
timestamp 1676037725
transform 1 0 173788 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1889
timestamp 1676037725
transform 1 0 174892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1901
timestamp 1676037725
transform 1 0 175996 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1905
timestamp 1676037725
transform 1 0 176364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1917
timestamp 1676037725
transform 1 0 177468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1929
timestamp 1676037725
transform 1 0 178572 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1933
timestamp 1676037725
transform 1 0 178940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1945
timestamp 1676037725
transform 1 0 180044 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_1957
timestamp 1676037725
transform 1 0 181148 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1961
timestamp 1676037725
transform 1 0 181516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1982
timestamp 1676037725
transform 1 0 183448 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1989
timestamp 1676037725
transform 1 0 184092 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1993
timestamp 1676037725
transform 1 0 184460 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2005
timestamp 1676037725
transform 1 0 185564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2013
timestamp 1676037725
transform 1 0 186300 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2017
timestamp 1676037725
transform 1 0 186668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2029
timestamp 1676037725
transform 1 0 187772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2041
timestamp 1676037725
transform 1 0 188876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2045
timestamp 1676037725
transform 1 0 189244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2053
timestamp 1676037725
transform 1 0 189980 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2064
timestamp 1676037725
transform 1 0 190992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2070
timestamp 1676037725
transform 1 0 191544 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2073
timestamp 1676037725
transform 1 0 191820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2085
timestamp 1676037725
transform 1 0 192924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2097
timestamp 1676037725
transform 1 0 194028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2101
timestamp 1676037725
transform 1 0 194396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2112
timestamp 1676037725
transform 1 0 195408 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2118
timestamp 1676037725
transform 1 0 195960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2126
timestamp 1676037725
transform 1 0 196696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2129
timestamp 1676037725
transform 1 0 196972 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2146
timestamp 1676037725
transform 1 0 198536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2152
timestamp 1676037725
transform 1 0 199088 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2157
timestamp 1676037725
transform 1 0 199548 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2169
timestamp 1676037725
transform 1 0 200652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2181
timestamp 1676037725
transform 1 0 201756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2185
timestamp 1676037725
transform 1 0 202124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2196
timestamp 1676037725
transform 1 0 203136 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2202
timestamp 1676037725
transform 1 0 203688 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2210
timestamp 1676037725
transform 1 0 204424 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2213
timestamp 1676037725
transform 1 0 204700 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2225
timestamp 1676037725
transform 1 0 205804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2231
timestamp 1676037725
transform 1 0 206356 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2239
timestamp 1676037725
transform 1 0 207092 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2241
timestamp 1676037725
transform 1 0 207276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2253
timestamp 1676037725
transform 1 0 208380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2265
timestamp 1676037725
transform 1 0 209484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2269
timestamp 1676037725
transform 1 0 209852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2277
timestamp 1676037725
transform 1 0 210588 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2283
timestamp 1676037725
transform 1 0 211140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2295
timestamp 1676037725
transform 1 0 212244 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2297
timestamp 1676037725
transform 1 0 212428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2307
timestamp 1676037725
transform 1 0 213348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2313
timestamp 1676037725
transform 1 0 213900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2321
timestamp 1676037725
transform 1 0 214636 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2325
timestamp 1676037725
transform 1 0 215004 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2337
timestamp 1676037725
transform 1 0 216108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2349
timestamp 1676037725
transform 1 0 217212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2353
timestamp 1676037725
transform 1 0 217580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2361
timestamp 1676037725
transform 1 0 218316 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2367
timestamp 1676037725
transform 1 0 218868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2379
timestamp 1676037725
transform 1 0 219972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2381
timestamp 1676037725
transform 1 0 220156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2389
timestamp 1676037725
transform 1 0 220892 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2395
timestamp 1676037725
transform 1 0 221444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2407
timestamp 1676037725
transform 1 0 222548 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2409
timestamp 1676037725
transform 1 0 222732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2421
timestamp 1676037725
transform 1 0 223836 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2427
timestamp 1676037725
transform 1 0 224388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2434
timestamp 1676037725
transform 1 0 225032 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2437
timestamp 1676037725
transform 1 0 225308 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2441
timestamp 1676037725
transform 1 0 225676 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2453
timestamp 1676037725
transform 1 0 226780 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2461
timestamp 1676037725
transform 1 0 227516 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2465
timestamp 1676037725
transform 1 0 227884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2473
timestamp 1676037725
transform 1 0 228620 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2479
timestamp 1676037725
transform 1 0 229172 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2491
timestamp 1676037725
transform 1 0 230276 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2493
timestamp 1676037725
transform 1 0 230460 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2505
timestamp 1676037725
transform 1 0 231564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2509
timestamp 1676037725
transform 1 0 231932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2516
timestamp 1676037725
transform 1 0 232576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2521
timestamp 1676037725
transform 1 0 233036 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2525
timestamp 1676037725
transform 1 0 233404 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_2537
timestamp 1676037725
transform 1 0 234508 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2545
timestamp 1676037725
transform 1 0 235244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2549
timestamp 1676037725
transform 1 0 235612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2557
timestamp 1676037725
transform 1 0 236348 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2563
timestamp 1676037725
transform 1 0 236900 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2575
timestamp 1676037725
transform 1 0 238004 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2577
timestamp 1676037725
transform 1 0 238188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2589
timestamp 1676037725
transform 1 0 239292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_2597
timestamp 1676037725
transform 1 0 240028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2603
timestamp 1676037725
transform 1 0 240580 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2605
timestamp 1676037725
transform 1 0 240764 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2617
timestamp 1676037725
transform 1 0 241868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2629
timestamp 1676037725
transform 1 0 242972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_2633
timestamp 1676037725
transform 1 0 243340 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_2641
timestamp 1676037725
transform 1 0 244076 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2647
timestamp 1676037725
transform 1 0 244628 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_2659
timestamp 1676037725
transform 1 0 245732 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2661
timestamp 1676037725
transform 1 0 245916 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2673
timestamp 1676037725
transform 1 0 247020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2685
timestamp 1676037725
transform 1 0 248124 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2689
timestamp 1676037725
transform 1 0 248492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2701
timestamp 1676037725
transform 1 0 249596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2713
timestamp 1676037725
transform 1 0 250700 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2717
timestamp 1676037725
transform 1 0 251068 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2729
timestamp 1676037725
transform 1 0 252172 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2741
timestamp 1676037725
transform 1 0 253276 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2745
timestamp 1676037725
transform 1 0 253644 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2757
timestamp 1676037725
transform 1 0 254748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2769
timestamp 1676037725
transform 1 0 255852 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2773
timestamp 1676037725
transform 1 0 256220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2785
timestamp 1676037725
transform 1 0 257324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2797
timestamp 1676037725
transform 1 0 258428 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2801
timestamp 1676037725
transform 1 0 258796 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2813
timestamp 1676037725
transform 1 0 259900 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2825
timestamp 1676037725
transform 1 0 261004 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2829
timestamp 1676037725
transform 1 0 261372 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2841
timestamp 1676037725
transform 1 0 262476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2853
timestamp 1676037725
transform 1 0 263580 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2857
timestamp 1676037725
transform 1 0 263948 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2869
timestamp 1676037725
transform 1 0 265052 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2881
timestamp 1676037725
transform 1 0 266156 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2885
timestamp 1676037725
transform 1 0 266524 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2897
timestamp 1676037725
transform 1 0 267628 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2909
timestamp 1676037725
transform 1 0 268732 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2913
timestamp 1676037725
transform 1 0 269100 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2925
timestamp 1676037725
transform 1 0 270204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2937
timestamp 1676037725
transform 1 0 271308 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2941
timestamp 1676037725
transform 1 0 271676 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2953
timestamp 1676037725
transform 1 0 272780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2965
timestamp 1676037725
transform 1 0 273884 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2969
timestamp 1676037725
transform 1 0 274252 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2981
timestamp 1676037725
transform 1 0 275356 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_2993
timestamp 1676037725
transform 1 0 276460 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_2997
timestamp 1676037725
transform 1 0 276828 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3009
timestamp 1676037725
transform 1 0 277932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3021
timestamp 1676037725
transform 1 0 279036 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3025
timestamp 1676037725
transform 1 0 279404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3037
timestamp 1676037725
transform 1 0 280508 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3049
timestamp 1676037725
transform 1 0 281612 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3053
timestamp 1676037725
transform 1 0 281980 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3065
timestamp 1676037725
transform 1 0 283084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3077
timestamp 1676037725
transform 1 0 284188 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3081
timestamp 1676037725
transform 1 0 284556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3093
timestamp 1676037725
transform 1 0 285660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3105
timestamp 1676037725
transform 1 0 286764 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3109
timestamp 1676037725
transform 1 0 287132 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3121
timestamp 1676037725
transform 1 0 288236 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3133
timestamp 1676037725
transform 1 0 289340 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3137
timestamp 1676037725
transform 1 0 289708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3149
timestamp 1676037725
transform 1 0 290812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3161
timestamp 1676037725
transform 1 0 291916 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3165
timestamp 1676037725
transform 1 0 292284 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3177
timestamp 1676037725
transform 1 0 293388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3189
timestamp 1676037725
transform 1 0 294492 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3193
timestamp 1676037725
transform 1 0 294860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3205
timestamp 1676037725
transform 1 0 295964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3217
timestamp 1676037725
transform 1 0 297068 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3221
timestamp 1676037725
transform 1 0 297436 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3233
timestamp 1676037725
transform 1 0 298540 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3245
timestamp 1676037725
transform 1 0 299644 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3249
timestamp 1676037725
transform 1 0 300012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3261
timestamp 1676037725
transform 1 0 301116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3273
timestamp 1676037725
transform 1 0 302220 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3277
timestamp 1676037725
transform 1 0 302588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3289
timestamp 1676037725
transform 1 0 303692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3301
timestamp 1676037725
transform 1 0 304796 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3305
timestamp 1676037725
transform 1 0 305164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3317
timestamp 1676037725
transform 1 0 306268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3329
timestamp 1676037725
transform 1 0 307372 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3333
timestamp 1676037725
transform 1 0 307740 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3345
timestamp 1676037725
transform 1 0 308844 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3357
timestamp 1676037725
transform 1 0 309948 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3361
timestamp 1676037725
transform 1 0 310316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3373
timestamp 1676037725
transform 1 0 311420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3385
timestamp 1676037725
transform 1 0 312524 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3389
timestamp 1676037725
transform 1 0 312892 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3401
timestamp 1676037725
transform 1 0 313996 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3413
timestamp 1676037725
transform 1 0 315100 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3417
timestamp 1676037725
transform 1 0 315468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3429
timestamp 1676037725
transform 1 0 316572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3441
timestamp 1676037725
transform 1 0 317676 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3445
timestamp 1676037725
transform 1 0 318044 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3457
timestamp 1676037725
transform 1 0 319148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3469
timestamp 1676037725
transform 1 0 320252 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3473
timestamp 1676037725
transform 1 0 320620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3485
timestamp 1676037725
transform 1 0 321724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3497
timestamp 1676037725
transform 1 0 322828 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3501
timestamp 1676037725
transform 1 0 323196 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3513
timestamp 1676037725
transform 1 0 324300 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3525
timestamp 1676037725
transform 1 0 325404 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3529
timestamp 1676037725
transform 1 0 325772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3541
timestamp 1676037725
transform 1 0 326876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3553
timestamp 1676037725
transform 1 0 327980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3557
timestamp 1676037725
transform 1 0 328348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3569
timestamp 1676037725
transform 1 0 329452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3581
timestamp 1676037725
transform 1 0 330556 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3585
timestamp 1676037725
transform 1 0 330924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3597
timestamp 1676037725
transform 1 0 332028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3609
timestamp 1676037725
transform 1 0 333132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3613
timestamp 1676037725
transform 1 0 333500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3625
timestamp 1676037725
transform 1 0 334604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3637
timestamp 1676037725
transform 1 0 335708 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3641
timestamp 1676037725
transform 1 0 336076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3653
timestamp 1676037725
transform 1 0 337180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3665
timestamp 1676037725
transform 1 0 338284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3669
timestamp 1676037725
transform 1 0 338652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3680
timestamp 1676037725
transform 1 0 339664 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3686
timestamp 1676037725
transform 1 0 340216 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3694
timestamp 1676037725
transform 1 0 340952 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3697
timestamp 1676037725
transform 1 0 341228 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3708
timestamp 1676037725
transform 1 0 342240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3714
timestamp 1676037725
transform 1 0 342792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3722
timestamp 1676037725
transform 1 0 343528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3725
timestamp 1676037725
transform 1 0 343804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3736
timestamp 1676037725
transform 1 0 344816 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3742
timestamp 1676037725
transform 1 0 345368 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3750
timestamp 1676037725
transform 1 0 346104 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3753
timestamp 1676037725
transform 1 0 346380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3761
timestamp 1676037725
transform 1 0 347116 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3767
timestamp 1676037725
transform 1 0 347668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3779
timestamp 1676037725
transform 1 0 348772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3781
timestamp 1676037725
transform 1 0 348956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3789
timestamp 1676037725
transform 1 0 349692 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3795
timestamp 1676037725
transform 1 0 350244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3807
timestamp 1676037725
transform 1 0 351348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3809
timestamp 1676037725
transform 1 0 351532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3817
timestamp 1676037725
transform 1 0 352268 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3823
timestamp 1676037725
transform 1 0 352820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3835
timestamp 1676037725
transform 1 0 353924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3837
timestamp 1676037725
transform 1 0 354108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3845
timestamp 1676037725
transform 1 0 354844 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3851
timestamp 1676037725
transform 1 0 355396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3863
timestamp 1676037725
transform 1 0 356500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3865
timestamp 1676037725
transform 1 0 356684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3873
timestamp 1676037725
transform 1 0 357420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3879
timestamp 1676037725
transform 1 0 357972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3883
timestamp 1676037725
transform 1 0 358340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3890
timestamp 1676037725
transform 1 0 358984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3893
timestamp 1676037725
transform 1 0 359260 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3897
timestamp 1676037725
transform 1 0 359628 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3909
timestamp 1676037725
transform 1 0 360732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3918
timestamp 1676037725
transform 1 0 361560 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3921
timestamp 1676037725
transform 1 0 361836 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3925
timestamp 1676037725
transform 1 0 362204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3937
timestamp 1676037725
transform 1 0 363308 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3945
timestamp 1676037725
transform 1 0 364044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3949
timestamp 1676037725
transform 1 0 364412 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3953
timestamp 1676037725
transform 1 0 364780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3971
timestamp 1676037725
transform 1 0 366436 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3975
timestamp 1676037725
transform 1 0 366804 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3977
timestamp 1676037725
transform 1 0 366988 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3981
timestamp 1676037725
transform 1 0 367356 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3989
timestamp 1676037725
transform 1 0 368092 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3998
timestamp 1676037725
transform 1 0 368920 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_4005
timestamp 1676037725
transform 1 0 369564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_4009
timestamp 1676037725
transform 1 0 369932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_4017
timestamp 1676037725
transform 1 0 370668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_4025
timestamp 1676037725
transform 1 0 371404 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_4031
timestamp 1676037725
transform 1 0 371956 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4033
timestamp 1676037725
transform 1 0 372140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_4051
timestamp 1676037725
transform 1 0 373796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4057
timestamp 1676037725
transform 1 0 374348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_4061
timestamp 1676037725
transform 1 0 374716 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4069
timestamp 1676037725
transform 1 0 375452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_4078
timestamp 1676037725
transform 1 0 376280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_4084
timestamp 1676037725
transform 1 0 376832 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_4089
timestamp 1676037725
transform 1 0 377292 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_4097
timestamp 1676037725
transform 1 0 378028 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_4104
timestamp 1676037725
transform 1 0 378672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_4110
timestamp 1676037725
transform 1 0 379224 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_4117
timestamp 1676037725
transform 1 0 379868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_4131
timestamp 1676037725
transform 1 0 381156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_4137
timestamp 1676037725
transform 1 0 381708 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_4143
timestamp 1676037725
transform 1 0 382260 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_4145
timestamp 1676037725
transform 1 0 382444 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_4157
timestamp 1676037725
transform 1 0 383548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_4163
timestamp 1676037725
transform 1 0 384100 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_4171
timestamp 1676037725
transform 1 0 384836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4173
timestamp 1676037725
transform 1 0 385020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4185
timestamp 1676037725
transform 1 0 386124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4197
timestamp 1676037725
transform 1 0 387228 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4201
timestamp 1676037725
transform 1 0 387596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4213
timestamp 1676037725
transform 1 0 388700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4225
timestamp 1676037725
transform 1 0 389804 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4229
timestamp 1676037725
transform 1 0 390172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4241
timestamp 1676037725
transform 1 0 391276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4253
timestamp 1676037725
transform 1 0 392380 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4257
timestamp 1676037725
transform 1 0 392748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4269
timestamp 1676037725
transform 1 0 393852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4281
timestamp 1676037725
transform 1 0 394956 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4285
timestamp 1676037725
transform 1 0 395324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4297
timestamp 1676037725
transform 1 0 396428 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4309
timestamp 1676037725
transform 1 0 397532 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4313
timestamp 1676037725
transform 1 0 397900 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4325
timestamp 1676037725
transform 1 0 399004 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4337
timestamp 1676037725
transform 1 0 400108 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4341
timestamp 1676037725
transform 1 0 400476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4353
timestamp 1676037725
transform 1 0 401580 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4365
timestamp 1676037725
transform 1 0 402684 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4369
timestamp 1676037725
transform 1 0 403052 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4381
timestamp 1676037725
transform 1 0 404156 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4393
timestamp 1676037725
transform 1 0 405260 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4397
timestamp 1676037725
transform 1 0 405628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4409
timestamp 1676037725
transform 1 0 406732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4421
timestamp 1676037725
transform 1 0 407836 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4425
timestamp 1676037725
transform 1 0 408204 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4437
timestamp 1676037725
transform 1 0 409308 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4449
timestamp 1676037725
transform 1 0 410412 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4453
timestamp 1676037725
transform 1 0 410780 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4465
timestamp 1676037725
transform 1 0 411884 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4477
timestamp 1676037725
transform 1 0 412988 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4481
timestamp 1676037725
transform 1 0 413356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4493
timestamp 1676037725
transform 1 0 414460 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4505
timestamp 1676037725
transform 1 0 415564 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4509
timestamp 1676037725
transform 1 0 415932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4521
timestamp 1676037725
transform 1 0 417036 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4533
timestamp 1676037725
transform 1 0 418140 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4537
timestamp 1676037725
transform 1 0 418508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4549
timestamp 1676037725
transform 1 0 419612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4561
timestamp 1676037725
transform 1 0 420716 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4565
timestamp 1676037725
transform 1 0 421084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4577
timestamp 1676037725
transform 1 0 422188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4589
timestamp 1676037725
transform 1 0 423292 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4593
timestamp 1676037725
transform 1 0 423660 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4605
timestamp 1676037725
transform 1 0 424764 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4617
timestamp 1676037725
transform 1 0 425868 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4621
timestamp 1676037725
transform 1 0 426236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4633
timestamp 1676037725
transform 1 0 427340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4645
timestamp 1676037725
transform 1 0 428444 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4649
timestamp 1676037725
transform 1 0 428812 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4661
timestamp 1676037725
transform 1 0 429916 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4673
timestamp 1676037725
transform 1 0 431020 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4677
timestamp 1676037725
transform 1 0 431388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4689
timestamp 1676037725
transform 1 0 432492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4701
timestamp 1676037725
transform 1 0 433596 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4705
timestamp 1676037725
transform 1 0 433964 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4717
timestamp 1676037725
transform 1 0 435068 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4729
timestamp 1676037725
transform 1 0 436172 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4733
timestamp 1676037725
transform 1 0 436540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4745
timestamp 1676037725
transform 1 0 437644 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4757
timestamp 1676037725
transform 1 0 438748 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4761
timestamp 1676037725
transform 1 0 439116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4773
timestamp 1676037725
transform 1 0 440220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4785
timestamp 1676037725
transform 1 0 441324 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4789
timestamp 1676037725
transform 1 0 441692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4801
timestamp 1676037725
transform 1 0 442796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4813
timestamp 1676037725
transform 1 0 443900 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4817
timestamp 1676037725
transform 1 0 444268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4829
timestamp 1676037725
transform 1 0 445372 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4841
timestamp 1676037725
transform 1 0 446476 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4845
timestamp 1676037725
transform 1 0 446844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4857
timestamp 1676037725
transform 1 0 447948 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4869
timestamp 1676037725
transform 1 0 449052 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4873
timestamp 1676037725
transform 1 0 449420 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4885
timestamp 1676037725
transform 1 0 450524 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4897
timestamp 1676037725
transform 1 0 451628 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4901
timestamp 1676037725
transform 1 0 451996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4913
timestamp 1676037725
transform 1 0 453100 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4925
timestamp 1676037725
transform 1 0 454204 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4929
timestamp 1676037725
transform 1 0 454572 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4941
timestamp 1676037725
transform 1 0 455676 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4953
timestamp 1676037725
transform 1 0 456780 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4957
timestamp 1676037725
transform 1 0 457148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4969
timestamp 1676037725
transform 1 0 458252 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_4981
timestamp 1676037725
transform 1 0 459356 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4985
timestamp 1676037725
transform 1 0 459724 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_4997
timestamp 1676037725
transform 1 0 460828 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5009
timestamp 1676037725
transform 1 0 461932 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5013
timestamp 1676037725
transform 1 0 462300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5025
timestamp 1676037725
transform 1 0 463404 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5037
timestamp 1676037725
transform 1 0 464508 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5041
timestamp 1676037725
transform 1 0 464876 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5053
timestamp 1676037725
transform 1 0 465980 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5065
timestamp 1676037725
transform 1 0 467084 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5069
timestamp 1676037725
transform 1 0 467452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5081
timestamp 1676037725
transform 1 0 468556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5093
timestamp 1676037725
transform 1 0 469660 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5097
timestamp 1676037725
transform 1 0 470028 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5109
timestamp 1676037725
transform 1 0 471132 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5121
timestamp 1676037725
transform 1 0 472236 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5125
timestamp 1676037725
transform 1 0 472604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5137
timestamp 1676037725
transform 1 0 473708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5149
timestamp 1676037725
transform 1 0 474812 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5153
timestamp 1676037725
transform 1 0 475180 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5165
timestamp 1676037725
transform 1 0 476284 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5177
timestamp 1676037725
transform 1 0 477388 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5181
timestamp 1676037725
transform 1 0 477756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5193
timestamp 1676037725
transform 1 0 478860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5205
timestamp 1676037725
transform 1 0 479964 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5209
timestamp 1676037725
transform 1 0 480332 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5221
timestamp 1676037725
transform 1 0 481436 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5233
timestamp 1676037725
transform 1 0 482540 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5237
timestamp 1676037725
transform 1 0 482908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5249
timestamp 1676037725
transform 1 0 484012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5261
timestamp 1676037725
transform 1 0 485116 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5265
timestamp 1676037725
transform 1 0 485484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5277
timestamp 1676037725
transform 1 0 486588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5289
timestamp 1676037725
transform 1 0 487692 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5293
timestamp 1676037725
transform 1 0 488060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5305
timestamp 1676037725
transform 1 0 489164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5317
timestamp 1676037725
transform 1 0 490268 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5321
timestamp 1676037725
transform 1 0 490636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5333
timestamp 1676037725
transform 1 0 491740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5345
timestamp 1676037725
transform 1 0 492844 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5349
timestamp 1676037725
transform 1 0 493212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5361
timestamp 1676037725
transform 1 0 494316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5373
timestamp 1676037725
transform 1 0 495420 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5377
timestamp 1676037725
transform 1 0 495788 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5389
timestamp 1676037725
transform 1 0 496892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5401
timestamp 1676037725
transform 1 0 497996 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5405
timestamp 1676037725
transform 1 0 498364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5417
timestamp 1676037725
transform 1 0 499468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5429
timestamp 1676037725
transform 1 0 500572 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5433
timestamp 1676037725
transform 1 0 500940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5445
timestamp 1676037725
transform 1 0 502044 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5457
timestamp 1676037725
transform 1 0 503148 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5461
timestamp 1676037725
transform 1 0 503516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5473
timestamp 1676037725
transform 1 0 504620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5485
timestamp 1676037725
transform 1 0 505724 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5489
timestamp 1676037725
transform 1 0 506092 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5501
timestamp 1676037725
transform 1 0 507196 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5513
timestamp 1676037725
transform 1 0 508300 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5517
timestamp 1676037725
transform 1 0 508668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5529
timestamp 1676037725
transform 1 0 509772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5541
timestamp 1676037725
transform 1 0 510876 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5545
timestamp 1676037725
transform 1 0 511244 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5557
timestamp 1676037725
transform 1 0 512348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5569
timestamp 1676037725
transform 1 0 513452 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5573
timestamp 1676037725
transform 1 0 513820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5585
timestamp 1676037725
transform 1 0 514924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5597
timestamp 1676037725
transform 1 0 516028 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5601
timestamp 1676037725
transform 1 0 516396 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5613
timestamp 1676037725
transform 1 0 517500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5625
timestamp 1676037725
transform 1 0 518604 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5629
timestamp 1676037725
transform 1 0 518972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5641
timestamp 1676037725
transform 1 0 520076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5653
timestamp 1676037725
transform 1 0 521180 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5657
timestamp 1676037725
transform 1 0 521548 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5669
timestamp 1676037725
transform 1 0 522652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5681
timestamp 1676037725
transform 1 0 523756 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5685
timestamp 1676037725
transform 1 0 524124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5697
timestamp 1676037725
transform 1 0 525228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_5709
timestamp 1676037725
transform 1 0 526332 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_5713
timestamp 1676037725
transform 1 0 526700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_5725
timestamp 1676037725
transform 1 0 527804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 528816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 528816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 528816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 528816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 528816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 528816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 528816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 528816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 528816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 528816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 528816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 528816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 528816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 528816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1676037725
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1676037725
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1676037725
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1676037725
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1676037725
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1676037725
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1676037725
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1676037725
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 119600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 124752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 129904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 135056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 140208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 145360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 150512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 153088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 155664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 160816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 163392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 165968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 168544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 171120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 173696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 176272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 178848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 181424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 184000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 186576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 189152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 191728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 194304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 196880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 199456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 202032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 204608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 207184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 209760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 212336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 214912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 217488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 220064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 222640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 225216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 227792 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 230368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 232944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 235520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 238096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 240672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 243248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 245824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 248400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 250976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 253552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 256128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 258704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 261280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 263856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 266432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 269008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 271584 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 274160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 276736 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 279312 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 281888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 284464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 287040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 289616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 292192 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 294768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 297344 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 299920 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 302496 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 305072 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 307648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 310224 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 312800 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 315376 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 317952 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 320528 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 323104 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 325680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 328256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 330832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 333408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 335984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 338560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 341136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 343712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 346288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 348864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 351440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 354016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 356592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 359168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 361744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 364320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 366896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 369472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 372048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 374624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 377200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 379776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 382352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 384928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 387504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 390080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 392656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 395232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 397808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 400384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 402960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 405536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 408112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 410688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 413264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 415840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 418416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 420992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 423568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 426144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 428720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 431296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 433872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 436448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 439024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 441600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 444176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 446752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 449328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 451904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 454480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 457056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 459632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 462208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 464784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 467360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 469936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 472512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 475088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 477664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 480240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 482816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 485392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 487968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 490544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 493120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 495696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 498272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 500848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 503424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 506000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 508576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 511152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 513728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 516304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 518880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 521456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 524032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 526608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 150512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 155664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 160816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 165968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 171120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 176272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 181424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 186576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 191728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 196880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 202032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 207184 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 212336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 217488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 222640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 227792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 232944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 238096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 243248 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 248400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 253552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 258704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 263856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 269008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 274160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 279312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 284464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 289616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 294768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 299920 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 305072 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 310224 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 315376 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 320528 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 325680 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 330832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 335984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 341136 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 346288 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 351440 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 356592 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 361744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 366896 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 372048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 377200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 382352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 387504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 392656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 397808 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 402960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 408112 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 413264 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 418416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 423568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 428720 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 433872 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 439024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 444176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 449328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 454480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 459632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 464784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 469936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 475088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 480240 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 485392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 490544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 495696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 500848 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 506000 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 511152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 516304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 521456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 526608 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 153088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 158240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 163392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 168544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 173696 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 178848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 184000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 189152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 194304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 199456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 204608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 209760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 214912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 220064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 225216 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 230368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 235520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 240672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 245824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 250976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 256128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 261280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 266432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 271584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 276736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 281888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 287040 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 292192 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 297344 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 302496 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 307648 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 312800 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 317952 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 323104 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 328256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 333408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 338560 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 343712 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 348864 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 354016 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 359168 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 364320 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 369472 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 374624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 379776 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 384928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 390080 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 395232 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 400384 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 405536 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 410688 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 415840 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 420992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 426144 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 431296 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 436448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 441600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 446752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 451904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 457056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 462208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 467360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 472512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 477664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 482816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 487968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 493120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 498272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 503424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 508576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 513728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 518880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 524032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 150512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 155664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 160816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 165968 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 171120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 176272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 181424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 186576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 191728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 196880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 202032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 207184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 212336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 217488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 222640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 227792 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 232944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 238096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 243248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 248400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 253552 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 258704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 263856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 269008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 274160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 279312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 284464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 289616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 294768 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 299920 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 305072 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 310224 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 315376 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 320528 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 325680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 330832 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 335984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 341136 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 346288 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 351440 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 356592 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 361744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 366896 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 372048 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 377200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 382352 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 387504 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 392656 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 397808 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 402960 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 408112 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 413264 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 418416 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 423568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 428720 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 433872 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 439024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 444176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 449328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 454480 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 459632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 464784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 469936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 475088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 480240 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 485392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 490544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 495696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 500848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 506000 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 511152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 516304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 521456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 526608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 153088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 158240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 163392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 168544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 173696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 178848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 184000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 189152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 194304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 199456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 204608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 209760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 214912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 220064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 225216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 230368 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 235520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 240672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 245824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 250976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 256128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 261280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 266432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 271584 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 276736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 281888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 287040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 292192 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 297344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 302496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 307648 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 312800 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 317952 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 323104 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 328256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 333408 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 338560 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 343712 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 348864 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 354016 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 359168 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 364320 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 369472 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 374624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 379776 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 384928 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 390080 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 395232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 400384 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 405536 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 410688 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 415840 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 420992 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 426144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 431296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 436448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 441600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 446752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 451904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 457056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 462208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 467360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 472512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 477664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 482816 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 487968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 493120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 498272 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 503424 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 508576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 513728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 518880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 524032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 150512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 155664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 160816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 165968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 171120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 176272 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 181424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 186576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 191728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 196880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 202032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 207184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 212336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 217488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 222640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 227792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 232944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 238096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 243248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 248400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 253552 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 258704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 263856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 269008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 274160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 279312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 284464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 289616 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 294768 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 299920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 305072 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 310224 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 315376 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 320528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 325680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 330832 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 335984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 341136 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 346288 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 351440 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 356592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 361744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 366896 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 372048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 377200 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 382352 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 387504 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 392656 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 397808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 402960 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 408112 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 413264 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 418416 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 423568 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 428720 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 433872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 439024 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 444176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 449328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 454480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 459632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 464784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 469936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 475088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 480240 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 485392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 490544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 495696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 500848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 506000 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 511152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 516304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 521456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 526608 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 153088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 158240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 163392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 168544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 173696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 178848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 184000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 189152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 194304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 199456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 204608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 209760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 214912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 220064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 225216 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 230368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 235520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 240672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 245824 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 250976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 256128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 261280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 266432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 271584 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 276736 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 281888 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 287040 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 292192 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 297344 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 302496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 307648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 312800 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 317952 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 323104 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 328256 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 333408 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 338560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 343712 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 348864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 354016 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 359168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 364320 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 369472 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 374624 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 379776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 384928 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 390080 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 395232 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 400384 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 405536 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 410688 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 415840 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 420992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 426144 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 431296 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 436448 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 441600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 446752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 451904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 457056 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 462208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 467360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 472512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 477664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 482816 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 487968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 493120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 498272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 503424 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 508576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 513728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 518880 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 524032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 150512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 155664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 160816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 165968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 171120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 176272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 181424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 186576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 191728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 196880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 202032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 207184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 212336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 217488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 222640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 227792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 232944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 238096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 243248 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 248400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 253552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 258704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 263856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 269008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 274160 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 279312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 284464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 289616 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 294768 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 299920 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 305072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 310224 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 315376 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 320528 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 325680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 330832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 335984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 341136 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 346288 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 351440 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 356592 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 361744 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 366896 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 372048 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 377200 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 382352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 387504 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 392656 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 397808 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 402960 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 408112 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 413264 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 418416 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 423568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 428720 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 433872 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 439024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 444176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 449328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 454480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 459632 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 464784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 469936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 475088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 480240 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 485392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 490544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 495696 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 500848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 506000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 511152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 516304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 521456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 526608 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 153088 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 158240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 163392 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 168544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 173696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 178848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 184000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 189152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 194304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 199456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 204608 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 209760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 214912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 220064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 225216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 230368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 235520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 240672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 245824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 250976 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 256128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 261280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 266432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 271584 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 276736 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 281888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 287040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 292192 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 297344 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 302496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 307648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 312800 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 317952 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 323104 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 328256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 333408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 338560 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 343712 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 348864 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 354016 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 359168 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 364320 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 369472 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 374624 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 379776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 384928 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 390080 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 395232 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 400384 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 405536 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 410688 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 415840 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 420992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 426144 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 431296 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 436448 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 441600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 446752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 451904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 457056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 462208 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 467360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 472512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 477664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 482816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 487968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 493120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 498272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 503424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 508576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 513728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 518880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 524032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1676037725
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1676037725
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1676037725
transform 1 0 150512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1676037725
transform 1 0 155664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1676037725
transform 1 0 160816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1676037725
transform 1 0 165968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1676037725
transform 1 0 171120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1676037725
transform 1 0 176272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1676037725
transform 1 0 181424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1676037725
transform 1 0 186576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1676037725
transform 1 0 191728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1676037725
transform 1 0 196880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1676037725
transform 1 0 202032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1676037725
transform 1 0 207184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1676037725
transform 1 0 212336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1676037725
transform 1 0 217488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1676037725
transform 1 0 222640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1676037725
transform 1 0 227792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1676037725
transform 1 0 232944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1676037725
transform 1 0 238096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1676037725
transform 1 0 243248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1676037725
transform 1 0 248400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1676037725
transform 1 0 253552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1676037725
transform 1 0 258704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1676037725
transform 1 0 263856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1676037725
transform 1 0 269008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1676037725
transform 1 0 274160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1676037725
transform 1 0 279312 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1676037725
transform 1 0 284464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1676037725
transform 1 0 289616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1676037725
transform 1 0 294768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1676037725
transform 1 0 299920 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1676037725
transform 1 0 305072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1676037725
transform 1 0 310224 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1676037725
transform 1 0 315376 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1676037725
transform 1 0 320528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1676037725
transform 1 0 325680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1676037725
transform 1 0 330832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1676037725
transform 1 0 335984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1676037725
transform 1 0 341136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1676037725
transform 1 0 346288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1676037725
transform 1 0 351440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1676037725
transform 1 0 356592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1676037725
transform 1 0 361744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1676037725
transform 1 0 366896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1676037725
transform 1 0 372048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1676037725
transform 1 0 377200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1676037725
transform 1 0 382352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1676037725
transform 1 0 387504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1676037725
transform 1 0 392656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1676037725
transform 1 0 397808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1676037725
transform 1 0 402960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1676037725
transform 1 0 408112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1676037725
transform 1 0 413264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1676037725
transform 1 0 418416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1676037725
transform 1 0 423568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1676037725
transform 1 0 428720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1676037725
transform 1 0 433872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1676037725
transform 1 0 439024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1676037725
transform 1 0 444176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1676037725
transform 1 0 449328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1676037725
transform 1 0 454480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1676037725
transform 1 0 459632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1676037725
transform 1 0 464784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1676037725
transform 1 0 469936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1676037725
transform 1 0 475088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1676037725
transform 1 0 480240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1676037725
transform 1 0 485392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1676037725
transform 1 0 490544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1676037725
transform 1 0 495696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1676037725
transform 1 0 500848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1676037725
transform 1 0 506000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1676037725
transform 1 0 511152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1676037725
transform 1 0 516304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1676037725
transform 1 0 521456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1676037725
transform 1 0 526608 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1676037725
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1676037725
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1676037725
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1676037725
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1676037725
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1676037725
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1676037725
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1676037725
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1676037725
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1676037725
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1676037725
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1676037725
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1676037725
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1676037725
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1676037725
transform 1 0 122176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1676037725
transform 1 0 127328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1676037725
transform 1 0 132480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1676037725
transform 1 0 137632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1676037725
transform 1 0 142784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1676037725
transform 1 0 147936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1676037725
transform 1 0 153088 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1676037725
transform 1 0 158240 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1676037725
transform 1 0 163392 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1676037725
transform 1 0 168544 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1676037725
transform 1 0 173696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1676037725
transform 1 0 178848 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1676037725
transform 1 0 184000 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1676037725
transform 1 0 189152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1676037725
transform 1 0 194304 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1676037725
transform 1 0 199456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1676037725
transform 1 0 204608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1676037725
transform 1 0 209760 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1676037725
transform 1 0 214912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1676037725
transform 1 0 220064 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1676037725
transform 1 0 225216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1676037725
transform 1 0 230368 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1676037725
transform 1 0 235520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1676037725
transform 1 0 240672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1676037725
transform 1 0 245824 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1676037725
transform 1 0 250976 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1676037725
transform 1 0 256128 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1676037725
transform 1 0 261280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1676037725
transform 1 0 266432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1676037725
transform 1 0 271584 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1676037725
transform 1 0 276736 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1676037725
transform 1 0 281888 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1676037725
transform 1 0 287040 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1676037725
transform 1 0 292192 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1676037725
transform 1 0 297344 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1676037725
transform 1 0 302496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1676037725
transform 1 0 307648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1676037725
transform 1 0 312800 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1676037725
transform 1 0 317952 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1676037725
transform 1 0 323104 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1676037725
transform 1 0 328256 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1676037725
transform 1 0 333408 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1676037725
transform 1 0 338560 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1676037725
transform 1 0 343712 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1676037725
transform 1 0 348864 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1676037725
transform 1 0 354016 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1676037725
transform 1 0 359168 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1676037725
transform 1 0 364320 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1676037725
transform 1 0 369472 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1676037725
transform 1 0 374624 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1676037725
transform 1 0 379776 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1676037725
transform 1 0 384928 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1676037725
transform 1 0 390080 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1676037725
transform 1 0 395232 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1676037725
transform 1 0 400384 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1676037725
transform 1 0 405536 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1676037725
transform 1 0 410688 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1676037725
transform 1 0 415840 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1676037725
transform 1 0 420992 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1676037725
transform 1 0 426144 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1676037725
transform 1 0 431296 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1676037725
transform 1 0 436448 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1676037725
transform 1 0 441600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1676037725
transform 1 0 446752 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1676037725
transform 1 0 451904 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1676037725
transform 1 0 457056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1676037725
transform 1 0 462208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1676037725
transform 1 0 467360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1676037725
transform 1 0 472512 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1676037725
transform 1 0 477664 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1676037725
transform 1 0 482816 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1676037725
transform 1 0 487968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1676037725
transform 1 0 493120 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1676037725
transform 1 0 498272 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1676037725
transform 1 0 503424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1676037725
transform 1 0 508576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1676037725
transform 1 0 513728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1676037725
transform 1 0 518880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1676037725
transform 1 0 524032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1676037725
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1676037725
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1676037725
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1676037725
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1676037725
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1676037725
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1676037725
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1676037725
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1676037725
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1676037725
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1676037725
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1676037725
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1676037725
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1676037725
transform 1 0 119600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1676037725
transform 1 0 124752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1676037725
transform 1 0 129904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1676037725
transform 1 0 135056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1676037725
transform 1 0 140208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1676037725
transform 1 0 145360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1676037725
transform 1 0 150512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1676037725
transform 1 0 155664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1676037725
transform 1 0 160816 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1676037725
transform 1 0 165968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1676037725
transform 1 0 171120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1676037725
transform 1 0 176272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1676037725
transform 1 0 181424 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1676037725
transform 1 0 186576 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1676037725
transform 1 0 191728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1676037725
transform 1 0 196880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1676037725
transform 1 0 202032 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1676037725
transform 1 0 207184 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1676037725
transform 1 0 212336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1676037725
transform 1 0 217488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1676037725
transform 1 0 222640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1676037725
transform 1 0 227792 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1676037725
transform 1 0 232944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1676037725
transform 1 0 238096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1676037725
transform 1 0 243248 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1676037725
transform 1 0 248400 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1676037725
transform 1 0 253552 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1676037725
transform 1 0 258704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1676037725
transform 1 0 263856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1676037725
transform 1 0 269008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1676037725
transform 1 0 274160 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1676037725
transform 1 0 279312 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1676037725
transform 1 0 284464 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1676037725
transform 1 0 289616 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1676037725
transform 1 0 294768 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1676037725
transform 1 0 299920 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1676037725
transform 1 0 305072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1676037725
transform 1 0 310224 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1676037725
transform 1 0 315376 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1676037725
transform 1 0 320528 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1676037725
transform 1 0 325680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1676037725
transform 1 0 330832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1676037725
transform 1 0 335984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1676037725
transform 1 0 341136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1676037725
transform 1 0 346288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1676037725
transform 1 0 351440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1676037725
transform 1 0 356592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1676037725
transform 1 0 361744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1676037725
transform 1 0 366896 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1676037725
transform 1 0 372048 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1676037725
transform 1 0 377200 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1676037725
transform 1 0 382352 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1676037725
transform 1 0 387504 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1676037725
transform 1 0 392656 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1676037725
transform 1 0 397808 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1676037725
transform 1 0 402960 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1676037725
transform 1 0 408112 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1676037725
transform 1 0 413264 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1676037725
transform 1 0 418416 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1676037725
transform 1 0 423568 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1676037725
transform 1 0 428720 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1676037725
transform 1 0 433872 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1676037725
transform 1 0 439024 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1676037725
transform 1 0 444176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1676037725
transform 1 0 449328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1676037725
transform 1 0 454480 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1676037725
transform 1 0 459632 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1676037725
transform 1 0 464784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1676037725
transform 1 0 469936 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1676037725
transform 1 0 475088 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1676037725
transform 1 0 480240 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1676037725
transform 1 0 485392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1676037725
transform 1 0 490544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1676037725
transform 1 0 495696 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1676037725
transform 1 0 500848 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1676037725
transform 1 0 506000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1676037725
transform 1 0 511152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1676037725
transform 1 0 516304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1676037725
transform 1 0 521456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1676037725
transform 1 0 526608 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1676037725
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1676037725
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1676037725
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1676037725
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1676037725
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1676037725
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1676037725
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1676037725
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1676037725
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1676037725
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1676037725
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1676037725
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1676037725
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1676037725
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1676037725
transform 1 0 122176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1676037725
transform 1 0 127328 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1676037725
transform 1 0 132480 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1676037725
transform 1 0 137632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1676037725
transform 1 0 142784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1676037725
transform 1 0 147936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1676037725
transform 1 0 153088 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1676037725
transform 1 0 158240 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1676037725
transform 1 0 163392 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1676037725
transform 1 0 168544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1676037725
transform 1 0 173696 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1676037725
transform 1 0 178848 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1676037725
transform 1 0 184000 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1676037725
transform 1 0 189152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1676037725
transform 1 0 194304 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1676037725
transform 1 0 199456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1676037725
transform 1 0 204608 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1676037725
transform 1 0 209760 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1676037725
transform 1 0 214912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1676037725
transform 1 0 220064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1676037725
transform 1 0 225216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1676037725
transform 1 0 230368 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1676037725
transform 1 0 235520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1676037725
transform 1 0 240672 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1676037725
transform 1 0 245824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1676037725
transform 1 0 250976 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1676037725
transform 1 0 256128 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1676037725
transform 1 0 261280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1676037725
transform 1 0 266432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1676037725
transform 1 0 271584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1676037725
transform 1 0 276736 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1676037725
transform 1 0 281888 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1676037725
transform 1 0 287040 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1676037725
transform 1 0 292192 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1676037725
transform 1 0 297344 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1676037725
transform 1 0 302496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1676037725
transform 1 0 307648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1676037725
transform 1 0 312800 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1676037725
transform 1 0 317952 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1676037725
transform 1 0 323104 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1676037725
transform 1 0 328256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1676037725
transform 1 0 333408 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1676037725
transform 1 0 338560 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1676037725
transform 1 0 343712 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1676037725
transform 1 0 348864 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1676037725
transform 1 0 354016 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1676037725
transform 1 0 359168 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1676037725
transform 1 0 364320 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1676037725
transform 1 0 369472 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1676037725
transform 1 0 374624 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1676037725
transform 1 0 379776 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1676037725
transform 1 0 384928 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1676037725
transform 1 0 390080 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1676037725
transform 1 0 395232 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1676037725
transform 1 0 400384 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1676037725
transform 1 0 405536 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1676037725
transform 1 0 410688 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1676037725
transform 1 0 415840 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1676037725
transform 1 0 420992 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1676037725
transform 1 0 426144 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1676037725
transform 1 0 431296 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1676037725
transform 1 0 436448 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1676037725
transform 1 0 441600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1676037725
transform 1 0 446752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1676037725
transform 1 0 451904 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1676037725
transform 1 0 457056 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1676037725
transform 1 0 462208 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1676037725
transform 1 0 467360 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1676037725
transform 1 0 472512 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1676037725
transform 1 0 477664 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1676037725
transform 1 0 482816 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1676037725
transform 1 0 487968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1676037725
transform 1 0 493120 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1676037725
transform 1 0 498272 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1676037725
transform 1 0 503424 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1676037725
transform 1 0 508576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1676037725
transform 1 0 513728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1676037725
transform 1 0 518880 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1676037725
transform 1 0 524032 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1676037725
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1676037725
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1676037725
transform 1 0 13984 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1676037725
transform 1 0 19136 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1676037725
transform 1 0 24288 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1676037725
transform 1 0 29440 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1676037725
transform 1 0 34592 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1676037725
transform 1 0 39744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1676037725
transform 1 0 44896 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1676037725
transform 1 0 50048 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1676037725
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1676037725
transform 1 0 55200 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1676037725
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1676037725
transform 1 0 60352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1676037725
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1676037725
transform 1 0 65504 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1676037725
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1676037725
transform 1 0 70656 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1676037725
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1676037725
transform 1 0 75808 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1676037725
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1676037725
transform 1 0 80960 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1676037725
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1676037725
transform 1 0 86112 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1676037725
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1676037725
transform 1 0 91264 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1676037725
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1676037725
transform 1 0 96416 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1676037725
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1676037725
transform 1 0 101568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1676037725
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1676037725
transform 1 0 106720 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1676037725
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1676037725
transform 1 0 111872 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1676037725
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1676037725
transform 1 0 117024 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1676037725
transform 1 0 119600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1676037725
transform 1 0 122176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1676037725
transform 1 0 124752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1676037725
transform 1 0 127328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1676037725
transform 1 0 129904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1676037725
transform 1 0 132480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1676037725
transform 1 0 135056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1676037725
transform 1 0 137632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1676037725
transform 1 0 140208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1676037725
transform 1 0 142784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1676037725
transform 1 0 145360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1676037725
transform 1 0 147936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1676037725
transform 1 0 150512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1676037725
transform 1 0 153088 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1676037725
transform 1 0 155664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1676037725
transform 1 0 158240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1676037725
transform 1 0 160816 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1676037725
transform 1 0 163392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1676037725
transform 1 0 165968 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1676037725
transform 1 0 168544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1676037725
transform 1 0 171120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1676037725
transform 1 0 173696 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1676037725
transform 1 0 176272 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1676037725
transform 1 0 178848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1676037725
transform 1 0 181424 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1676037725
transform 1 0 184000 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1676037725
transform 1 0 186576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1676037725
transform 1 0 189152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1676037725
transform 1 0 191728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1676037725
transform 1 0 194304 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1676037725
transform 1 0 196880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1676037725
transform 1 0 199456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1676037725
transform 1 0 202032 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1676037725
transform 1 0 204608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1676037725
transform 1 0 207184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1676037725
transform 1 0 209760 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1676037725
transform 1 0 212336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1676037725
transform 1 0 214912 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1676037725
transform 1 0 217488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1676037725
transform 1 0 220064 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1676037725
transform 1 0 222640 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1676037725
transform 1 0 225216 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1676037725
transform 1 0 227792 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1676037725
transform 1 0 230368 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1676037725
transform 1 0 232944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1676037725
transform 1 0 235520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1676037725
transform 1 0 238096 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1676037725
transform 1 0 240672 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1676037725
transform 1 0 243248 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1676037725
transform 1 0 245824 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1676037725
transform 1 0 248400 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1676037725
transform 1 0 250976 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1676037725
transform 1 0 253552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1676037725
transform 1 0 256128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1676037725
transform 1 0 258704 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1676037725
transform 1 0 261280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1676037725
transform 1 0 263856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1676037725
transform 1 0 266432 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1676037725
transform 1 0 269008 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1676037725
transform 1 0 271584 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1676037725
transform 1 0 274160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1676037725
transform 1 0 276736 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1676037725
transform 1 0 279312 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1676037725
transform 1 0 281888 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1676037725
transform 1 0 284464 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1676037725
transform 1 0 287040 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1676037725
transform 1 0 289616 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1676037725
transform 1 0 292192 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1676037725
transform 1 0 294768 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1676037725
transform 1 0 297344 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1676037725
transform 1 0 299920 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1676037725
transform 1 0 302496 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1676037725
transform 1 0 305072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1676037725
transform 1 0 307648 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1676037725
transform 1 0 310224 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1676037725
transform 1 0 312800 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1676037725
transform 1 0 315376 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1676037725
transform 1 0 317952 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1676037725
transform 1 0 320528 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1676037725
transform 1 0 323104 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1676037725
transform 1 0 325680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1676037725
transform 1 0 328256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1676037725
transform 1 0 330832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1676037725
transform 1 0 333408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1676037725
transform 1 0 335984 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1676037725
transform 1 0 338560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1676037725
transform 1 0 341136 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1676037725
transform 1 0 343712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1676037725
transform 1 0 346288 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1676037725
transform 1 0 348864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1676037725
transform 1 0 351440 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1676037725
transform 1 0 354016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1676037725
transform 1 0 356592 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1676037725
transform 1 0 359168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1676037725
transform 1 0 361744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1676037725
transform 1 0 364320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1676037725
transform 1 0 366896 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1676037725
transform 1 0 369472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1676037725
transform 1 0 372048 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1676037725
transform 1 0 374624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1676037725
transform 1 0 377200 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1676037725
transform 1 0 379776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1676037725
transform 1 0 382352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1676037725
transform 1 0 384928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1676037725
transform 1 0 387504 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1676037725
transform 1 0 390080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1676037725
transform 1 0 392656 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1676037725
transform 1 0 395232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1676037725
transform 1 0 397808 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1676037725
transform 1 0 400384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1676037725
transform 1 0 402960 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1676037725
transform 1 0 405536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1676037725
transform 1 0 408112 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1676037725
transform 1 0 410688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1676037725
transform 1 0 413264 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1676037725
transform 1 0 415840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1676037725
transform 1 0 418416 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1676037725
transform 1 0 420992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1676037725
transform 1 0 423568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1676037725
transform 1 0 426144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1676037725
transform 1 0 428720 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1676037725
transform 1 0 431296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1676037725
transform 1 0 433872 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1676037725
transform 1 0 436448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1676037725
transform 1 0 439024 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1676037725
transform 1 0 441600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1676037725
transform 1 0 444176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1676037725
transform 1 0 446752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1676037725
transform 1 0 449328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1676037725
transform 1 0 451904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1676037725
transform 1 0 454480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1676037725
transform 1 0 457056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1676037725
transform 1 0 459632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1676037725
transform 1 0 462208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1676037725
transform 1 0 464784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1676037725
transform 1 0 467360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1676037725
transform 1 0 469936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1676037725
transform 1 0 472512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1676037725
transform 1 0 475088 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1676037725
transform 1 0 477664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1676037725
transform 1 0 480240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1676037725
transform 1 0 482816 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1676037725
transform 1 0 485392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1676037725
transform 1 0 487968 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1676037725
transform 1 0 490544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1676037725
transform 1 0 493120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1676037725
transform 1 0 495696 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1676037725
transform 1 0 498272 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1676037725
transform 1 0 500848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1676037725
transform 1 0 503424 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1676037725
transform 1 0 506000 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1676037725
transform 1 0 508576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1676037725
transform 1 0 511152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1676037725
transform 1 0 513728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1676037725
transform 1 0 516304 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1676037725
transform 1 0 518880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1676037725
transform 1 0 521456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1676037725
transform 1 0 524032 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1676037725
transform 1 0 526608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[0\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[1\].u_buf
timestamp 1676037725
transform -1 0 2116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[2\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[3\].u_buf
timestamp 1676037725
transform -1 0 4692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[4\].u_buf
timestamp 1676037725
transform -1 0 7268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[5\].u_buf
timestamp 1676037725
transform -1 0 7268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[6\].u_buf
timestamp 1676037725
transform -1 0 9844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[7\].u_buf
timestamp 1676037725
transform -1 0 9844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[8\].u_buf
timestamp 1676037725
transform -1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[9\].u_buf
timestamp 1676037725
transform -1 0 12420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[10\].u_buf
timestamp 1676037725
transform -1 0 14996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[11\].u_buf
timestamp 1676037725
transform -1 0 14996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[12\].u_buf
timestamp 1676037725
transform -1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[13\].u_buf
timestamp 1676037725
transform -1 0 17572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[14\].u_buf
timestamp 1676037725
transform -1 0 20148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[15\].u_buf
timestamp 1676037725
transform -1 0 20148 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[16\].u_buf
timestamp 1676037725
transform -1 0 22724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[17\].u_buf
timestamp 1676037725
transform -1 0 22724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[18\].u_buf
timestamp 1676037725
transform -1 0 25300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[19\].u_buf
timestamp 1676037725
transform -1 0 25300 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[20\].u_buf
timestamp 1676037725
transform -1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[21\].u_buf
timestamp 1676037725
transform -1 0 27876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[22\].u_buf
timestamp 1676037725
transform -1 0 30452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[23\].u_buf
timestamp 1676037725
transform -1 0 30452 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[24\].u_buf
timestamp 1676037725
transform -1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[25\].u_buf
timestamp 1676037725
transform -1 0 33028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[26\].u_buf
timestamp 1676037725
transform -1 0 35604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[27\].u_buf
timestamp 1676037725
transform -1 0 35604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[28\].u_buf
timestamp 1676037725
transform -1 0 38180 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[29\].u_buf
timestamp 1676037725
transform -1 0 38180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[30\].u_buf
timestamp 1676037725
transform -1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[31\].u_buf
timestamp 1676037725
transform -1 0 40756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[32\].u_buf
timestamp 1676037725
transform -1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[33\].u_buf
timestamp 1676037725
transform -1 0 43332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[34\].u_buf
timestamp 1676037725
transform -1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[35\].u_buf
timestamp 1676037725
transform -1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[36\].u_buf
timestamp 1676037725
transform -1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[37\].u_buf
timestamp 1676037725
transform -1 0 48484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[38\].u_buf
timestamp 1676037725
transform -1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[39\].u_buf
timestamp 1676037725
transform -1 0 51060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[40\].u_buf
timestamp 1676037725
transform -1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[41\].u_buf
timestamp 1676037725
transform -1 0 53636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[42\].u_buf
timestamp 1676037725
transform -1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[43\].u_buf
timestamp 1676037725
transform -1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[44\].u_buf
timestamp 1676037725
transform -1 0 58788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[45\].u_buf
timestamp 1676037725
transform -1 0 58788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[46\].u_buf
timestamp 1676037725
transform -1 0 61364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[47\].u_buf
timestamp 1676037725
transform -1 0 61364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[48\].u_buf
timestamp 1676037725
transform -1 0 63940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[49\].u_buf
timestamp 1676037725
transform -1 0 63940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[50\].u_buf
timestamp 1676037725
transform -1 0 66516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[51\].u_buf
timestamp 1676037725
transform -1 0 66516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[52\].u_buf
timestamp 1676037725
transform -1 0 69092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[53\].u_buf
timestamp 1676037725
transform -1 0 69092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[54\].u_buf
timestamp 1676037725
transform -1 0 71668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[55\].u_buf
timestamp 1676037725
transform -1 0 71668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[56\].u_buf
timestamp 1676037725
transform -1 0 74244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[57\].u_buf
timestamp 1676037725
transform -1 0 74244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[58\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 76820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[59\].u_buf
timestamp 1676037725
transform -1 0 76820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[60\].u_buf
timestamp 1676037725
transform -1 0 79396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[61\].u_buf
timestamp 1676037725
transform -1 0 79396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[62\].u_buf
timestamp 1676037725
transform -1 0 81972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[63\].u_buf
timestamp 1676037725
transform -1 0 81972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[64\].u_buf
timestamp 1676037725
transform -1 0 84548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[65\].u_buf
timestamp 1676037725
transform -1 0 84548 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[66\].u_buf
timestamp 1676037725
transform -1 0 87124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[67\].u_buf
timestamp 1676037725
transform -1 0 87124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[68\].u_buf
timestamp 1676037725
transform -1 0 89700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[69\].u_buf
timestamp 1676037725
transform -1 0 89700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[70\].u_buf
timestamp 1676037725
transform -1 0 92276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[71\].u_buf
timestamp 1676037725
transform -1 0 92276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[72\].u_buf
timestamp 1676037725
transform -1 0 94852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[73\].u_buf
timestamp 1676037725
transform -1 0 94852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[74\].u_buf
timestamp 1676037725
transform -1 0 97428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[75\].u_buf
timestamp 1676037725
transform -1 0 97428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[76\].u_buf
timestamp 1676037725
transform -1 0 100004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[77\].u_buf
timestamp 1676037725
transform -1 0 100004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[78\].u_buf
timestamp 1676037725
transform -1 0 102580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[79\].u_buf
timestamp 1676037725
transform -1 0 102580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[80\].u_buf
timestamp 1676037725
transform -1 0 105156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[81\].u_buf
timestamp 1676037725
transform -1 0 105156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[82\].u_buf
timestamp 1676037725
transform -1 0 107732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[83\].u_buf
timestamp 1676037725
transform -1 0 107732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[84\].u_buf
timestamp 1676037725
transform -1 0 110308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[85\].u_buf
timestamp 1676037725
transform -1 0 110308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[86\].u_buf
timestamp 1676037725
transform -1 0 112884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[87\].u_buf
timestamp 1676037725
transform -1 0 112884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[88\].u_buf
timestamp 1676037725
transform -1 0 115460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[89\].u_buf
timestamp 1676037725
transform -1 0 115460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[90\].u_buf
timestamp 1676037725
transform -1 0 118036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[91\].u_buf
timestamp 1676037725
transform -1 0 118036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[92\].u_buf
timestamp 1676037725
transform -1 0 120612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[93\].u_buf
timestamp 1676037725
transform -1 0 120612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[94\].u_buf
timestamp 1676037725
transform -1 0 123188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[95\].u_buf
timestamp 1676037725
transform -1 0 123188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[96\].u_buf
timestamp 1676037725
transform -1 0 125764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[97\].u_buf
timestamp 1676037725
transform -1 0 125764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[98\].u_buf
timestamp 1676037725
transform -1 0 128340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[99\].u_buf
timestamp 1676037725
transform -1 0 128340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[100\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 130916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[101\].u_buf
timestamp 1676037725
transform -1 0 130916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[102\].u_buf
timestamp 1676037725
transform -1 0 133492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[103\].u_buf
timestamp 1676037725
transform -1 0 133492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  u_rp\[104\].u_buf
timestamp 1676037725
transform -1 0 136068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  u_rp\[105\].u_buf
timestamp 1676037725
transform -1 0 136068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  u_rp\[106\].u_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 138644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[107\].u_buf
timestamp 1676037725
transform -1 0 141220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  u_rp\[108\].u_buf
timestamp 1676037725
transform -1 0 143796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[109\].u_buf
timestamp 1676037725
transform -1 0 146372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  u_rp\[110\].u_buf
timestamp 1676037725
transform -1 0 148948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[111\].u_buf
timestamp 1676037725
transform -1 0 151524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  u_rp\[112\].u_buf
timestamp 1676037725
transform -1 0 154100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[113\].u_buf
timestamp 1676037725
transform -1 0 156676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  u_rp\[114\].u_buf
timestamp 1676037725
transform -1 0 159252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[115\].u_buf
timestamp 1676037725
transform -1 0 161828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[116\].u_buf
timestamp 1676037725
transform -1 0 164404 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[117\].u_buf
timestamp 1676037725
transform -1 0 166980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[118\].u_buf
timestamp 1676037725
transform -1 0 169556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[119\].u_buf
timestamp 1676037725
transform -1 0 172132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[120\].u_buf
timestamp 1676037725
transform -1 0 174708 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[121\].u_buf
timestamp 1676037725
transform -1 0 177284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[122\].u_buf
timestamp 1676037725
transform -1 0 179860 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[123\].u_buf
timestamp 1676037725
transform -1 0 182436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[124\].u_buf
timestamp 1676037725
transform -1 0 185012 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[125\].u_buf
timestamp 1676037725
transform -1 0 187588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[126\].u_buf
timestamp 1676037725
transform -1 0 190164 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[127\].u_buf
timestamp 1676037725
transform -1 0 192740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  u_rp\[128\].u_buf
timestamp 1676037725
transform -1 0 195316 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  u_rp\[129\].u_buf
timestamp 1676037725
transform -1 0 197892 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[130\].u_buf
timestamp 1676037725
transform -1 0 200468 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[131\].u_buf
timestamp 1676037725
transform -1 0 203044 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[132\].u_buf
timestamp 1676037725
transform -1 0 205620 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[133\].u_buf
timestamp 1676037725
transform -1 0 208196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[134\].u_buf
timestamp 1676037725
transform -1 0 210772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[135\].u_buf
timestamp 1676037725
transform -1 0 213348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[136\].u_buf
timestamp 1676037725
transform -1 0 215924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[137\].u_buf
timestamp 1676037725
transform -1 0 218500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[138\].u_buf
timestamp 1676037725
transform -1 0 221076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[139\].u_buf
timestamp 1676037725
transform -1 0 223652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  u_rp\[140\].u_buf
timestamp 1676037725
transform -1 0 226228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[141\].u_buf
timestamp 1676037725
transform -1 0 228804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[142\].u_buf
timestamp 1676037725
transform -1 0 231380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[143\].u_buf
timestamp 1676037725
transform -1 0 233956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[144\].u_buf
timestamp 1676037725
transform -1 0 236532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[145\].u_buf
timestamp 1676037725
transform -1 0 239108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[146\].u_buf
timestamp 1676037725
transform -1 0 241684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[147\].u_buf
timestamp 1676037725
transform -1 0 244260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[148\].u_buf
timestamp 1676037725
transform -1 0 246836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[149\].u_buf
timestamp 1676037725
transform -1 0 249412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[150\].u_buf
timestamp 1676037725
transform -1 0 251988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[151\].u_buf
timestamp 1676037725
transform -1 0 254564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[152\].u_buf
timestamp 1676037725
transform -1 0 257140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[153\].u_buf
timestamp 1676037725
transform -1 0 259716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[154\].u_buf
timestamp 1676037725
transform -1 0 262292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[155\].u_buf
timestamp 1676037725
transform -1 0 264868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[156\].u_buf
timestamp 1676037725
transform -1 0 267444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[157\].u_buf
timestamp 1676037725
transform -1 0 270020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[158\].u_buf
timestamp 1676037725
transform -1 0 272596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[159\].u_buf
timestamp 1676037725
transform -1 0 275172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[160\].u_buf
timestamp 1676037725
transform -1 0 277748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[161\].u_buf
timestamp 1676037725
transform -1 0 280324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[162\].u_buf
timestamp 1676037725
transform -1 0 282900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[163\].u_buf
timestamp 1676037725
transform -1 0 285476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[164\].u_buf
timestamp 1676037725
transform -1 0 288052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[165\].u_buf
timestamp 1676037725
transform -1 0 290628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[166\].u_buf
timestamp 1676037725
transform -1 0 293204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[167\].u_buf
timestamp 1676037725
transform -1 0 295780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[168\].u_buf
timestamp 1676037725
transform -1 0 298356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[169\].u_buf
timestamp 1676037725
transform -1 0 300932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[170\].u_buf
timestamp 1676037725
transform -1 0 303508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[171\].u_buf
timestamp 1676037725
transform -1 0 306084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[172\].u_buf
timestamp 1676037725
transform -1 0 308660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[173\].u_buf
timestamp 1676037725
transform -1 0 311236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[174\].u_buf
timestamp 1676037725
transform -1 0 313812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[175\].u_buf
timestamp 1676037725
transform -1 0 316388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[176\].u_buf
timestamp 1676037725
transform -1 0 318964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[177\].u_buf
timestamp 1676037725
transform -1 0 321540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[178\].u_buf
timestamp 1676037725
transform -1 0 324116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[179\].u_buf
timestamp 1676037725
transform -1 0 326692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[180\].u_buf
timestamp 1676037725
transform -1 0 329268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[181\].u_buf
timestamp 1676037725
transform -1 0 331844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[182\].u_buf
timestamp 1676037725
transform -1 0 334420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[183\].u_buf
timestamp 1676037725
transform -1 0 336996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[184\].u_buf
timestamp 1676037725
transform -1 0 339572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[185\].u_buf
timestamp 1676037725
transform -1 0 342148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[186\].u_buf
timestamp 1676037725
transform -1 0 344724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[187\].u_buf
timestamp 1676037725
transform -1 0 347300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[188\].u_buf
timestamp 1676037725
transform -1 0 349876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[189\].u_buf
timestamp 1676037725
transform -1 0 352452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[190\].u_buf
timestamp 1676037725
transform -1 0 355028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[191\].u_buf
timestamp 1676037725
transform -1 0 357604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[192\].u_buf
timestamp 1676037725
transform -1 0 360180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[193\].u_buf
timestamp 1676037725
transform -1 0 362756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[194\].u_buf
timestamp 1676037725
transform -1 0 365332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[195\].u_buf
timestamp 1676037725
transform -1 0 367908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[196\].u_buf
timestamp 1676037725
transform -1 0 370484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[197\].u_buf
timestamp 1676037725
transform -1 0 373060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[198\].u_buf
timestamp 1676037725
transform -1 0 375636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[199\].u_buf
timestamp 1676037725
transform -1 0 378212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[200\].u_buf
timestamp 1676037725
transform -1 0 380788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[201\].u_buf
timestamp 1676037725
transform -1 0 383364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[202\].u_buf
timestamp 1676037725
transform -1 0 385940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[203\].u_buf
timestamp 1676037725
transform -1 0 388516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[204\].u_buf
timestamp 1676037725
transform -1 0 391092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[205\].u_buf
timestamp 1676037725
transform -1 0 393668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[206\].u_buf
timestamp 1676037725
transform -1 0 396244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[207\].u_buf
timestamp 1676037725
transform -1 0 398820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[208\].u_buf
timestamp 1676037725
transform -1 0 401396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[209\].u_buf
timestamp 1676037725
transform -1 0 403972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[210\].u_buf
timestamp 1676037725
transform -1 0 406548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[211\].u_buf
timestamp 1676037725
transform -1 0 409124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[212\].u_buf
timestamp 1676037725
transform -1 0 411700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[213\].u_buf
timestamp 1676037725
transform -1 0 414276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[214\].u_buf
timestamp 1676037725
transform -1 0 416852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[215\].u_buf
timestamp 1676037725
transform -1 0 419428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[216\].u_buf
timestamp 1676037725
transform -1 0 422004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[217\].u_buf
timestamp 1676037725
transform -1 0 424580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[218\].u_buf
timestamp 1676037725
transform -1 0 427156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[219\].u_buf
timestamp 1676037725
transform -1 0 429732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[220\].u_buf
timestamp 1676037725
transform -1 0 432308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[221\].u_buf
timestamp 1676037725
transform -1 0 434884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[222\].u_buf
timestamp 1676037725
transform -1 0 437460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[223\].u_buf
timestamp 1676037725
transform -1 0 440036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[224\].u_buf
timestamp 1676037725
transform -1 0 442612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[225\].u_buf
timestamp 1676037725
transform -1 0 445188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[226\].u_buf
timestamp 1676037725
transform -1 0 447764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[227\].u_buf
timestamp 1676037725
transform -1 0 450340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[228\].u_buf
timestamp 1676037725
transform -1 0 452916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[229\].u_buf
timestamp 1676037725
transform -1 0 455492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[230\].u_buf
timestamp 1676037725
transform -1 0 458068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[231\].u_buf
timestamp 1676037725
transform -1 0 460644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[232\].u_buf
timestamp 1676037725
transform -1 0 463220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[233\].u_buf
timestamp 1676037725
transform -1 0 465796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[234\].u_buf
timestamp 1676037725
transform -1 0 468372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[235\].u_buf
timestamp 1676037725
transform -1 0 470948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[236\].u_buf
timestamp 1676037725
transform -1 0 473524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[237\].u_buf
timestamp 1676037725
transform -1 0 476100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[238\].u_buf
timestamp 1676037725
transform -1 0 478676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[239\].u_buf
timestamp 1676037725
transform -1 0 481252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[240\].u_buf
timestamp 1676037725
transform -1 0 483828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[241\].u_buf
timestamp 1676037725
transform -1 0 486404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[242\].u_buf
timestamp 1676037725
transform -1 0 488980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[243\].u_buf
timestamp 1676037725
transform -1 0 491556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[244\].u_buf
timestamp 1676037725
transform -1 0 494132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[245\].u_buf
timestamp 1676037725
transform -1 0 496708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[246\].u_buf
timestamp 1676037725
transform -1 0 499284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[247\].u_buf
timestamp 1676037725
transform -1 0 501860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[248\].u_buf
timestamp 1676037725
transform -1 0 504436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[249\].u_buf
timestamp 1676037725
transform -1 0 507012 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[250\].u_buf
timestamp 1676037725
transform -1 0 509588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[251\].u_buf
timestamp 1676037725
transform -1 0 512164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  u_rp\[252\].u_buf
timestamp 1676037725
transform -1 0 514740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  wire1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 95404 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire2
timestamp 1676037725
transform 1 0 147200 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire3
timestamp 1676037725
transform 1 0 145636 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire4
timestamp 1676037725
transform 1 0 144532 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire5
timestamp 1676037725
transform 1 0 145636 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire6
timestamp 1676037725
transform 1 0 143704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire7
timestamp 1676037725
transform 1 0 142140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire8
timestamp 1676037725
transform 1 0 141036 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire9
timestamp 1676037725
transform 1 0 141312 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire10
timestamp 1676037725
transform 1 0 140208 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire11
timestamp 1676037725
transform 1 0 138736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire12
timestamp 1676037725
transform 1 0 137540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire13
timestamp 1676037725
transform 1 0 137908 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire14
timestamp 1676037725
transform 1 0 136712 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire15
timestamp 1676037725
transform 1 0 94208 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire16
timestamp 1676037725
transform 1 0 135240 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire17
timestamp 1676037725
transform 1 0 134136 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire18
timestamp 1676037725
transform 1 0 134320 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire19
timestamp 1676037725
transform 1 0 133216 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire20
timestamp 1676037725
transform 1 0 131744 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire21
timestamp 1676037725
transform 1 0 130640 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire22
timestamp 1676037725
transform 1 0 131376 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire23
timestamp 1676037725
transform 1 0 94484 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire24
timestamp 1676037725
transform 1 0 130180 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire25
timestamp 1676037725
transform 1 0 128340 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire26
timestamp 1676037725
transform 1 0 127144 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire27
timestamp 1676037725
transform 1 0 127420 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire28
timestamp 1676037725
transform 1 0 126224 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire29
timestamp 1676037725
transform 1 0 125028 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire30
timestamp 1676037725
transform 1 0 92828 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire31
timestamp 1676037725
transform 1 0 123740 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire32
timestamp 1676037725
transform 1 0 124016 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire33
timestamp 1676037725
transform 1 0 122820 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire34
timestamp 1676037725
transform 1 0 121532 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire35
timestamp 1676037725
transform 1 0 120336 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire36
timestamp 1676037725
transform 1 0 120612 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire37
timestamp 1676037725
transform 1 0 119416 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire38
timestamp 1676037725
transform 1 0 93288 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire39
timestamp 1676037725
transform 1 0 118128 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire40
timestamp 1676037725
transform 1 0 117300 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire41
timestamp 1676037725
transform 1 0 117300 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire42
timestamp 1676037725
transform 1 0 116012 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire43
timestamp 1676037725
transform 1 0 114724 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire44
timestamp 1676037725
transform 1 0 113528 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire45
timestamp 1676037725
transform 1 0 113436 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire46
timestamp 1676037725
transform 1 0 92184 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire47
timestamp 1676037725
transform 1 0 112240 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire48
timestamp 1676037725
transform 1 0 112148 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire49
timestamp 1676037725
transform 1 0 110216 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire50
timestamp 1676037725
transform 1 0 110308 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire51
timestamp 1676037725
transform 1 0 109204 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire52
timestamp 1676037725
transform 1 0 107916 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire53
timestamp 1676037725
transform 1 0 106812 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire54
timestamp 1676037725
transform 1 0 106996 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire55
timestamp 1676037725
transform 1 0 105616 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire56
timestamp 1676037725
transform 1 0 104604 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire57
timestamp 1676037725
transform 1 0 103408 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire58
timestamp 1676037725
transform 1 0 103132 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire59
timestamp 1676037725
transform 1 0 102212 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire60
timestamp 1676037725
transform 1 0 91080 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire61
timestamp 1676037725
transform 1 0 101200 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire62
timestamp 1676037725
transform 1 0 101292 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire63
timestamp 1676037725
transform 1 0 100004 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire64
timestamp 1676037725
transform 1 0 98900 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire65
timestamp 1676037725
transform 1 0 99268 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire66
timestamp 1676037725
transform 1 0 271032 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire67
timestamp 1676037725
transform 1 0 97796 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire68
timestamp 1676037725
transform 1 0 269836 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire69
timestamp 1676037725
transform 1 0 268548 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire70
timestamp 1676037725
transform 1 0 267352 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire71
timestamp 1676037725
transform 1 0 266156 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire72
timestamp 1676037725
transform 1 0 264868 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire73
timestamp 1676037725
transform 1 0 263672 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire74
timestamp 1676037725
transform 1 0 262476 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire75
timestamp 1676037725
transform 1 0 261280 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire76
timestamp 1676037725
transform 1 0 260084 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire77
timestamp 1676037725
transform 1 0 258888 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire78
timestamp 1676037725
transform 1 0 96600 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire79
timestamp 1676037725
transform 1 0 257692 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire80
timestamp 1676037725
transform 1 0 256496 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire81
timestamp 1676037725
transform 1 0 255116 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire82
timestamp 1676037725
transform 1 0 254104 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire83
timestamp 1676037725
transform 1 0 252540 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire84
timestamp 1676037725
transform 1 0 96784 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire85
timestamp 1676037725
transform 1 0 251344 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire86
timestamp 1676037725
transform 1 0 250148 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire87
timestamp 1676037725
transform 1 0 150788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire88
timestamp 1676037725
transform 1 0 149132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire89
timestamp 1676037725
transform 1 0 148028 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire90
timestamp 1676037725
transform 1 0 148396 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire91
timestamp 1676037725
transform 1 0 91540 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire92
timestamp 1676037725
transform -1 0 236348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire93
timestamp 1676037725
transform -1 0 232576 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire94
timestamp 1676037725
transform -1 0 228620 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire95
timestamp 1676037725
transform -1 0 225032 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire96
timestamp 1676037725
transform -1 0 121992 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire97
timestamp 1676037725
transform -1 0 220892 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire98
timestamp 1676037725
transform -1 0 218316 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire99
timestamp 1676037725
transform -1 0 213348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire100
timestamp 1676037725
transform -1 0 210588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire101
timestamp 1676037725
transform -1 0 205804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire102
timestamp 1676037725
transform -1 0 203136 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire103
timestamp 1676037725
transform -1 0 198536 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire104
timestamp 1676037725
transform -1 0 195408 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire105
timestamp 1676037725
transform -1 0 190992 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire106
timestamp 1676037725
transform -1 0 187772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire107
timestamp 1676037725
transform -1 0 183448 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire108
timestamp 1676037725
transform -1 0 180136 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire109
timestamp 1676037725
transform -1 0 175812 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire110
timestamp 1676037725
transform -1 0 172592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire111
timestamp 1676037725
transform -1 0 168268 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire112
timestamp 1676037725
transform -1 0 165048 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire113
timestamp 1676037725
transform -1 0 160632 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire114
timestamp 1676037725
transform -1 0 157412 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire115
timestamp 1676037725
transform -1 0 152904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire116
timestamp 1676037725
transform -1 0 149868 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire117
timestamp 1676037725
transform -1 0 114356 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire118
timestamp 1676037725
transform -1 0 145176 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire119
timestamp 1676037725
transform -1 0 142232 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire120
timestamp 1676037725
transform -1 0 137172 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire121
timestamp 1676037725
transform -1 0 132112 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire122
timestamp 1676037725
transform -1 0 383548 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire123
timestamp 1676037725
transform -1 0 381156 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire124
timestamp 1676037725
transform -1 0 378672 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire125
timestamp 1676037725
transform -1 0 376280 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire126
timestamp 1676037725
transform -1 0 373796 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire127
timestamp 1676037725
transform -1 0 371404 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire128
timestamp 1676037725
transform -1 0 368920 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire129
timestamp 1676037725
transform -1 0 366436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire130
timestamp 1676037725
transform -1 0 364044 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire131
timestamp 1676037725
transform -1 0 361560 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire132
timestamp 1676037725
transform -1 0 358984 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire133
timestamp 1676037725
transform -1 0 357420 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire134
timestamp 1676037725
transform -1 0 354844 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire135
timestamp 1676037725
transform -1 0 352268 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire136
timestamp 1676037725
transform -1 0 349692 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire137
timestamp 1676037725
transform -1 0 347116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  wire138
timestamp 1676037725
transform -1 0 344816 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire139
timestamp 1676037725
transform -1 0 342240 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire140
timestamp 1676037725
transform -1 0 339664 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire141
timestamp 1676037725
transform -1 0 336996 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire142
timestamp 1676037725
transform -1 0 332028 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire143
timestamp 1676037725
transform -1 0 327060 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire144
timestamp 1676037725
transform -1 0 322000 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire145
timestamp 1676037725
transform -1 0 317032 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire146
timestamp 1676037725
transform -1 0 311972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire147
timestamp 1676037725
transform -1 0 127052 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire148
timestamp 1676037725
transform -1 0 307004 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire149
timestamp 1676037725
transform -1 0 301944 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire150
timestamp 1676037725
transform -1 0 296884 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire151
timestamp 1676037725
transform -1 0 291916 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire152
timestamp 1676037725
transform -1 0 286856 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire153
timestamp 1676037725
transform -1 0 281704 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire154
timestamp 1676037725
transform -1 0 276552 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire155
timestamp 1676037725
transform -1 0 271676 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire156
timestamp 1676037725
transform -1 0 266616 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire157
timestamp 1676037725
transform -1 0 261556 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire158
timestamp 1676037725
transform -1 0 256496 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  wire159
timestamp 1676037725
transform -1 0 252080 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  wire160
timestamp 1676037725
transform -1 0 244076 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  wire161
timestamp 1676037725
transform -1 0 240028 0 -1 9792
box -38 -48 590 592
<< labels >>
flabel metal1 s 74 0 130 800 0 FreeSans 224 90 0 0 ch_in[0]
port 0 nsew signal input
flabel metal1 s 108874 0 108930 800 0 FreeSans 224 90 0 0 ch_in[100]
port 1 nsew signal input
flabel metal1 s 109962 0 110018 800 0 FreeSans 224 90 0 0 ch_in[101]
port 2 nsew signal input
flabel metal1 s 255550 11200 255606 12000 0 FreeSans 224 90 0 0 ch_in[102]
port 3 nsew signal input
flabel metal1 s 112138 0 112194 800 0 FreeSans 224 90 0 0 ch_in[103]
port 4 nsew signal input
flabel metal1 s 113226 0 113282 800 0 FreeSans 224 90 0 0 ch_in[104]
port 5 nsew signal input
flabel metal1 s 257182 11200 257238 12000 0 FreeSans 224 90 0 0 ch_in[105]
port 6 nsew signal input
flabel metal1 s 120026 0 120082 800 0 FreeSans 224 90 0 0 ch_in[106]
port 7 nsew signal input
flabel metal1 s 360610 11200 360666 12000 0 FreeSans 224 90 0 0 ch_in[107]
port 8 nsew signal input
flabel metal1 s 124378 0 124434 800 0 FreeSans 224 90 0 0 ch_in[108]
port 9 nsew signal input
flabel metal1 s 361698 11200 361754 12000 0 FreeSans 224 90 0 0 ch_in[109]
port 10 nsew signal input
flabel metal1 s 10954 0 11010 800 0 FreeSans 224 90 0 0 ch_in[10]
port 11 nsew signal input
flabel metal1 s 128730 0 128786 800 0 FreeSans 224 90 0 0 ch_in[110]
port 12 nsew signal input
flabel metal1 s 362786 11200 362842 12000 0 FreeSans 224 90 0 0 ch_in[111]
port 13 nsew signal input
flabel metal1 s 133082 0 133138 800 0 FreeSans 224 90 0 0 ch_in[112]
port 14 nsew signal input
flabel metal1 s 363874 11200 363930 12000 0 FreeSans 224 90 0 0 ch_in[113]
port 15 nsew signal input
flabel metal1 s 137434 0 137490 800 0 FreeSans 224 90 0 0 ch_in[114]
port 16 nsew signal input
flabel metal1 s 364962 11200 365018 12000 0 FreeSans 224 90 0 0 ch_in[115]
port 17 nsew signal input
flabel metal1 s 141786 0 141842 800 0 FreeSans 224 90 0 0 ch_in[116]
port 18 nsew signal input
flabel metal1 s 366050 11200 366106 12000 0 FreeSans 224 90 0 0 ch_in[117]
port 19 nsew signal input
flabel metal1 s 146138 0 146194 800 0 FreeSans 224 90 0 0 ch_in[118]
port 20 nsew signal input
flabel metal1 s 367138 11200 367194 12000 0 FreeSans 224 90 0 0 ch_in[119]
port 21 nsew signal input
flabel metal1 s 12042 0 12098 800 0 FreeSans 224 90 0 0 ch_in[11]
port 22 nsew signal input
flabel metal1 s 150490 0 150546 800 0 FreeSans 224 90 0 0 ch_in[120]
port 23 nsew signal input
flabel metal1 s 368226 11200 368282 12000 0 FreeSans 224 90 0 0 ch_in[121]
port 24 nsew signal input
flabel metal1 s 154842 0 154898 800 0 FreeSans 224 90 0 0 ch_in[122]
port 25 nsew signal input
flabel metal1 s 369314 11200 369370 12000 0 FreeSans 224 90 0 0 ch_in[123]
port 26 nsew signal input
flabel metal1 s 159194 0 159250 800 0 FreeSans 224 90 0 0 ch_in[124]
port 27 nsew signal input
flabel metal1 s 370402 11200 370458 12000 0 FreeSans 224 90 0 0 ch_in[125]
port 28 nsew signal input
flabel metal1 s 162050 0 162106 800 0 FreeSans 224 90 0 0 ch_in[126]
port 29 nsew signal input
flabel metal1 s 371490 11200 371546 12000 0 FreeSans 224 90 0 0 ch_in[127]
port 30 nsew signal input
flabel metal1 s 166402 0 166458 800 0 FreeSans 224 90 0 0 ch_in[128]
port 31 nsew signal input
flabel metal1 s 372578 11200 372634 12000 0 FreeSans 224 90 0 0 ch_in[129]
port 32 nsew signal input
flabel metal1 s 206590 11200 206646 12000 0 FreeSans 224 90 0 0 ch_in[12]
port 33 nsew signal input
flabel metal1 s 170754 0 170810 800 0 FreeSans 224 90 0 0 ch_in[130]
port 34 nsew signal input
flabel metal1 s 373666 11200 373722 12000 0 FreeSans 224 90 0 0 ch_in[131]
port 35 nsew signal input
flabel metal1 s 175106 0 175162 800 0 FreeSans 224 90 0 0 ch_in[132]
port 36 nsew signal input
flabel metal1 s 374754 11200 374810 12000 0 FreeSans 224 90 0 0 ch_in[133]
port 37 nsew signal input
flabel metal1 s 179458 0 179514 800 0 FreeSans 224 90 0 0 ch_in[134]
port 38 nsew signal input
flabel metal1 s 375842 11200 375898 12000 0 FreeSans 224 90 0 0 ch_in[135]
port 39 nsew signal input
flabel metal1 s 183810 0 183866 800 0 FreeSans 224 90 0 0 ch_in[136]
port 40 nsew signal input
flabel metal1 s 376930 11200 376986 12000 0 FreeSans 224 90 0 0 ch_in[137]
port 41 nsew signal input
flabel metal1 s 188162 0 188218 800 0 FreeSans 224 90 0 0 ch_in[138]
port 42 nsew signal input
flabel metal1 s 378018 11200 378074 12000 0 FreeSans 224 90 0 0 ch_in[139]
port 43 nsew signal input
flabel metal1 s 14218 0 14274 800 0 FreeSans 224 90 0 0 ch_in[13]
port 44 nsew signal input
flabel metal1 s 192514 0 192570 800 0 FreeSans 224 90 0 0 ch_in[140]
port 45 nsew signal input
flabel metal1 s 379106 11200 379162 12000 0 FreeSans 224 90 0 0 ch_in[141]
port 46 nsew signal input
flabel metal1 s 379650 11200 379706 12000 0 FreeSans 224 90 0 0 ch_in[142]
port 47 nsew signal input
flabel metal1 s 380194 11200 380250 12000 0 FreeSans 224 90 0 0 ch_in[143]
port 48 nsew signal input
flabel metal1 s 380738 11200 380794 12000 0 FreeSans 224 90 0 0 ch_in[144]
port 49 nsew signal input
flabel metal1 s 381282 11200 381338 12000 0 FreeSans 224 90 0 0 ch_in[145]
port 50 nsew signal input
flabel metal1 s 381826 11200 381882 12000 0 FreeSans 224 90 0 0 ch_in[146]
port 51 nsew signal input
flabel metal1 s 382370 11200 382426 12000 0 FreeSans 224 90 0 0 ch_in[147]
port 52 nsew signal input
flabel metal1 s 382914 11200 382970 12000 0 FreeSans 224 90 0 0 ch_in[148]
port 53 nsew signal input
flabel metal1 s 383458 11200 383514 12000 0 FreeSans 224 90 0 0 ch_in[149]
port 54 nsew signal input
flabel metal1 s 15306 0 15362 800 0 FreeSans 224 90 0 0 ch_in[14]
port 55 nsew signal input
flabel metal1 s 384002 11200 384058 12000 0 FreeSans 224 90 0 0 ch_in[150]
port 56 nsew signal input
flabel metal1 s 384546 11200 384602 12000 0 FreeSans 224 90 0 0 ch_in[151]
port 57 nsew signal input
flabel metal1 s 385090 11200 385146 12000 0 FreeSans 224 90 0 0 ch_in[152]
port 58 nsew signal input
flabel metal1 s 385634 11200 385690 12000 0 FreeSans 224 90 0 0 ch_in[153]
port 59 nsew signal input
flabel metal1 s 386178 11200 386234 12000 0 FreeSans 224 90 0 0 ch_in[154]
port 60 nsew signal input
flabel metal1 s 386722 11200 386778 12000 0 FreeSans 224 90 0 0 ch_in[155]
port 61 nsew signal input
flabel metal1 s 387266 11200 387322 12000 0 FreeSans 224 90 0 0 ch_in[156]
port 62 nsew signal input
flabel metal1 s 387810 11200 387866 12000 0 FreeSans 224 90 0 0 ch_in[157]
port 63 nsew signal input
flabel metal1 s 388354 11200 388410 12000 0 FreeSans 224 90 0 0 ch_in[158]
port 64 nsew signal input
flabel metal1 s 388898 11200 388954 12000 0 FreeSans 224 90 0 0 ch_in[159]
port 65 nsew signal input
flabel metal1 s 16394 0 16450 800 0 FreeSans 224 90 0 0 ch_in[15]
port 66 nsew signal input
flabel metal1 s 389442 11200 389498 12000 0 FreeSans 224 90 0 0 ch_in[160]
port 67 nsew signal input
flabel metal1 s 389986 11200 390042 12000 0 FreeSans 224 90 0 0 ch_in[161]
port 68 nsew signal input
flabel metal1 s 390530 11200 390586 12000 0 FreeSans 224 90 0 0 ch_in[162]
port 69 nsew signal input
flabel metal1 s 391074 11200 391130 12000 0 FreeSans 224 90 0 0 ch_in[163]
port 70 nsew signal input
flabel metal1 s 391618 11200 391674 12000 0 FreeSans 224 90 0 0 ch_in[164]
port 71 nsew signal input
flabel metal1 s 392162 11200 392218 12000 0 FreeSans 224 90 0 0 ch_in[165]
port 72 nsew signal input
flabel metal1 s 392706 11200 392762 12000 0 FreeSans 224 90 0 0 ch_in[166]
port 73 nsew signal input
flabel metal1 s 393250 11200 393306 12000 0 FreeSans 224 90 0 0 ch_in[167]
port 74 nsew signal input
flabel metal1 s 393794 11200 393850 12000 0 FreeSans 224 90 0 0 ch_in[168]
port 75 nsew signal input
flabel metal1 s 394338 11200 394394 12000 0 FreeSans 224 90 0 0 ch_in[169]
port 76 nsew signal input
flabel metal1 s 208766 11200 208822 12000 0 FreeSans 224 90 0 0 ch_in[16]
port 77 nsew signal input
flabel metal1 s 394882 11200 394938 12000 0 FreeSans 224 90 0 0 ch_in[170]
port 78 nsew signal input
flabel metal1 s 395426 11200 395482 12000 0 FreeSans 224 90 0 0 ch_in[171]
port 79 nsew signal input
flabel metal1 s 395970 11200 396026 12000 0 FreeSans 224 90 0 0 ch_in[172]
port 80 nsew signal input
flabel metal1 s 396514 11200 396570 12000 0 FreeSans 224 90 0 0 ch_in[173]
port 81 nsew signal input
flabel metal1 s 397058 11200 397114 12000 0 FreeSans 224 90 0 0 ch_in[174]
port 82 nsew signal input
flabel metal1 s 397602 11200 397658 12000 0 FreeSans 224 90 0 0 ch_in[175]
port 83 nsew signal input
flabel metal1 s 398146 11200 398202 12000 0 FreeSans 224 90 0 0 ch_in[176]
port 84 nsew signal input
flabel metal1 s 398690 11200 398746 12000 0 FreeSans 224 90 0 0 ch_in[177]
port 85 nsew signal input
flabel metal1 s 399234 11200 399290 12000 0 FreeSans 224 90 0 0 ch_in[178]
port 86 nsew signal input
flabel metal1 s 399778 11200 399834 12000 0 FreeSans 224 90 0 0 ch_in[179]
port 87 nsew signal input
flabel metal1 s 18570 0 18626 800 0 FreeSans 224 90 0 0 ch_in[17]
port 88 nsew signal input
flabel metal1 s 400322 11200 400378 12000 0 FreeSans 224 90 0 0 ch_in[180]
port 89 nsew signal input
flabel metal1 s 400866 11200 400922 12000 0 FreeSans 224 90 0 0 ch_in[181]
port 90 nsew signal input
flabel metal1 s 401410 11200 401466 12000 0 FreeSans 224 90 0 0 ch_in[182]
port 91 nsew signal input
flabel metal1 s 401954 11200 402010 12000 0 FreeSans 224 90 0 0 ch_in[183]
port 92 nsew signal input
flabel metal1 s 402498 11200 402554 12000 0 FreeSans 224 90 0 0 ch_in[184]
port 93 nsew signal input
flabel metal1 s 403042 11200 403098 12000 0 FreeSans 224 90 0 0 ch_in[185]
port 94 nsew signal input
flabel metal1 s 403586 11200 403642 12000 0 FreeSans 224 90 0 0 ch_in[186]
port 95 nsew signal input
flabel metal1 s 404130 11200 404186 12000 0 FreeSans 224 90 0 0 ch_in[187]
port 96 nsew signal input
flabel metal1 s 440034 11200 440090 12000 0 FreeSans 224 90 0 0 ch_in[188]
port 97 nsew signal input
flabel metal1 s 440306 11200 440362 12000 0 FreeSans 224 90 0 0 ch_in[189]
port 98 nsew signal input
flabel metal1 s 19658 0 19714 800 0 FreeSans 224 90 0 0 ch_in[18]
port 99 nsew signal input
flabel metal1 s 440578 11200 440634 12000 0 FreeSans 224 90 0 0 ch_in[190]
port 100 nsew signal input
flabel metal1 s 440850 11200 440906 12000 0 FreeSans 224 90 0 0 ch_in[191]
port 101 nsew signal input
flabel metal1 s 441122 11200 441178 12000 0 FreeSans 224 90 0 0 ch_in[192]
port 102 nsew signal input
flabel metal1 s 441394 11200 441450 12000 0 FreeSans 224 90 0 0 ch_in[193]
port 103 nsew signal input
flabel metal1 s 441666 11200 441722 12000 0 FreeSans 224 90 0 0 ch_in[194]
port 104 nsew signal input
flabel metal1 s 441938 11200 441994 12000 0 FreeSans 224 90 0 0 ch_in[195]
port 105 nsew signal input
flabel metal1 s 442210 11200 442266 12000 0 FreeSans 224 90 0 0 ch_in[196]
port 106 nsew signal input
flabel metal1 s 442482 11200 442538 12000 0 FreeSans 224 90 0 0 ch_in[197]
port 107 nsew signal input
flabel metal1 s 442754 11200 442810 12000 0 FreeSans 224 90 0 0 ch_in[198]
port 108 nsew signal input
flabel metal1 s 443026 11200 443082 12000 0 FreeSans 224 90 0 0 ch_in[199]
port 109 nsew signal input
flabel metal1 s 20746 0 20802 800 0 FreeSans 224 90 0 0 ch_in[19]
port 110 nsew signal input
flabel metal1 s 1162 0 1218 800 0 FreeSans 224 90 0 0 ch_in[1]
port 111 nsew signal input
flabel metal1 s 443298 11200 443354 12000 0 FreeSans 224 90 0 0 ch_in[200]
port 112 nsew signal input
flabel metal1 s 443570 11200 443626 12000 0 FreeSans 224 90 0 0 ch_in[201]
port 113 nsew signal input
flabel metal1 s 443842 11200 443898 12000 0 FreeSans 224 90 0 0 ch_in[202]
port 114 nsew signal input
flabel metal1 s 444114 11200 444170 12000 0 FreeSans 224 90 0 0 ch_in[203]
port 115 nsew signal input
flabel metal1 s 444386 11200 444442 12000 0 FreeSans 224 90 0 0 ch_in[204]
port 116 nsew signal input
flabel metal1 s 444658 11200 444714 12000 0 FreeSans 224 90 0 0 ch_in[205]
port 117 nsew signal input
flabel metal1 s 444930 11200 444986 12000 0 FreeSans 224 90 0 0 ch_in[206]
port 118 nsew signal input
flabel metal1 s 445202 11200 445258 12000 0 FreeSans 224 90 0 0 ch_in[207]
port 119 nsew signal input
flabel metal1 s 445474 11200 445530 12000 0 FreeSans 224 90 0 0 ch_in[208]
port 120 nsew signal input
flabel metal1 s 445746 11200 445802 12000 0 FreeSans 224 90 0 0 ch_in[209]
port 121 nsew signal input
flabel metal1 s 210942 11200 210998 12000 0 FreeSans 224 90 0 0 ch_in[20]
port 122 nsew signal input
flabel metal1 s 446018 11200 446074 12000 0 FreeSans 224 90 0 0 ch_in[210]
port 123 nsew signal input
flabel metal1 s 446290 11200 446346 12000 0 FreeSans 224 90 0 0 ch_in[211]
port 124 nsew signal input
flabel metal1 s 446562 11200 446618 12000 0 FreeSans 224 90 0 0 ch_in[212]
port 125 nsew signal input
flabel metal1 s 446834 11200 446890 12000 0 FreeSans 224 90 0 0 ch_in[213]
port 126 nsew signal input
flabel metal1 s 447106 11200 447162 12000 0 FreeSans 224 90 0 0 ch_in[214]
port 127 nsew signal input
flabel metal1 s 447378 11200 447434 12000 0 FreeSans 224 90 0 0 ch_in[215]
port 128 nsew signal input
flabel metal1 s 447650 11200 447706 12000 0 FreeSans 224 90 0 0 ch_in[216]
port 129 nsew signal input
flabel metal1 s 447922 11200 447978 12000 0 FreeSans 224 90 0 0 ch_in[217]
port 130 nsew signal input
flabel metal1 s 448194 11200 448250 12000 0 FreeSans 224 90 0 0 ch_in[218]
port 131 nsew signal input
flabel metal1 s 448466 11200 448522 12000 0 FreeSans 224 90 0 0 ch_in[219]
port 132 nsew signal input
flabel metal1 s 22922 0 22978 800 0 FreeSans 224 90 0 0 ch_in[21]
port 133 nsew signal input
flabel metal1 s 480018 11200 480074 12000 0 FreeSans 224 90 0 0 ch_in[220]
port 134 nsew signal input
flabel metal1 s 480290 11200 480346 12000 0 FreeSans 224 90 0 0 ch_in[221]
port 135 nsew signal input
flabel metal1 s 480562 11200 480618 12000 0 FreeSans 224 90 0 0 ch_in[222]
port 136 nsew signal input
flabel metal1 s 480834 11200 480890 12000 0 FreeSans 224 90 0 0 ch_in[223]
port 137 nsew signal input
flabel metal1 s 481106 11200 481162 12000 0 FreeSans 224 90 0 0 ch_in[224]
port 138 nsew signal input
flabel metal1 s 481378 11200 481434 12000 0 FreeSans 224 90 0 0 ch_in[225]
port 139 nsew signal input
flabel metal1 s 481650 11200 481706 12000 0 FreeSans 224 90 0 0 ch_in[226]
port 140 nsew signal input
flabel metal1 s 481922 11200 481978 12000 0 FreeSans 224 90 0 0 ch_in[227]
port 141 nsew signal input
flabel metal1 s 482194 11200 482250 12000 0 FreeSans 224 90 0 0 ch_in[228]
port 142 nsew signal input
flabel metal1 s 482466 11200 482522 12000 0 FreeSans 224 90 0 0 ch_in[229]
port 143 nsew signal input
flabel metal1 s 24010 0 24066 800 0 FreeSans 224 90 0 0 ch_in[22]
port 144 nsew signal input
flabel metal1 s 482738 11200 482794 12000 0 FreeSans 224 90 0 0 ch_in[230]
port 145 nsew signal input
flabel metal1 s 483010 11200 483066 12000 0 FreeSans 224 90 0 0 ch_in[231]
port 146 nsew signal input
flabel metal1 s 483282 11200 483338 12000 0 FreeSans 224 90 0 0 ch_in[232]
port 147 nsew signal input
flabel metal1 s 483554 11200 483610 12000 0 FreeSans 224 90 0 0 ch_in[233]
port 148 nsew signal input
flabel metal1 s 483826 11200 483882 12000 0 FreeSans 224 90 0 0 ch_in[234]
port 149 nsew signal input
flabel metal1 s 484098 11200 484154 12000 0 FreeSans 224 90 0 0 ch_in[235]
port 150 nsew signal input
flabel metal1 s 484370 11200 484426 12000 0 FreeSans 224 90 0 0 ch_in[236]
port 151 nsew signal input
flabel metal1 s 484642 11200 484698 12000 0 FreeSans 224 90 0 0 ch_in[237]
port 152 nsew signal input
flabel metal1 s 484914 11200 484970 12000 0 FreeSans 224 90 0 0 ch_in[238]
port 153 nsew signal input
flabel metal1 s 485186 11200 485242 12000 0 FreeSans 224 90 0 0 ch_in[239]
port 154 nsew signal input
flabel metal1 s 25098 0 25154 800 0 FreeSans 224 90 0 0 ch_in[23]
port 155 nsew signal input
flabel metal1 s 485458 11200 485514 12000 0 FreeSans 224 90 0 0 ch_in[240]
port 156 nsew signal input
flabel metal1 s 485730 11200 485786 12000 0 FreeSans 224 90 0 0 ch_in[241]
port 157 nsew signal input
flabel metal1 s 486002 11200 486058 12000 0 FreeSans 224 90 0 0 ch_in[242]
port 158 nsew signal input
flabel metal1 s 486274 11200 486330 12000 0 FreeSans 224 90 0 0 ch_in[243]
port 159 nsew signal input
flabel metal1 s 486546 11200 486602 12000 0 FreeSans 224 90 0 0 ch_in[244]
port 160 nsew signal input
flabel metal1 s 486818 11200 486874 12000 0 FreeSans 224 90 0 0 ch_in[245]
port 161 nsew signal input
flabel metal1 s 487090 11200 487146 12000 0 FreeSans 224 90 0 0 ch_in[246]
port 162 nsew signal input
flabel metal1 s 487362 11200 487418 12000 0 FreeSans 224 90 0 0 ch_in[247]
port 163 nsew signal input
flabel metal1 s 487634 11200 487690 12000 0 FreeSans 224 90 0 0 ch_in[248]
port 164 nsew signal input
flabel metal1 s 487906 11200 487962 12000 0 FreeSans 224 90 0 0 ch_in[249]
port 165 nsew signal input
flabel metal1 s 213118 11200 213174 12000 0 FreeSans 224 90 0 0 ch_in[24]
port 166 nsew signal input
flabel metal1 s 488178 11200 488234 12000 0 FreeSans 224 90 0 0 ch_in[250]
port 167 nsew signal input
flabel metal1 s 488450 11200 488506 12000 0 FreeSans 224 90 0 0 ch_in[251]
port 168 nsew signal input
flabel metal1 s 499330 0 499386 800 0 FreeSans 224 90 0 0 ch_in[252]
port 169 nsew signal input
flabel metal1 s 27274 0 27330 800 0 FreeSans 224 90 0 0 ch_in[25]
port 170 nsew signal input
flabel metal1 s 28362 0 28418 800 0 FreeSans 224 90 0 0 ch_in[26]
port 171 nsew signal input
flabel metal1 s 214750 11200 214806 12000 0 FreeSans 224 90 0 0 ch_in[27]
port 172 nsew signal input
flabel metal1 s 30538 0 30594 800 0 FreeSans 224 90 0 0 ch_in[28]
port 173 nsew signal input
flabel metal1 s 31626 0 31682 800 0 FreeSans 224 90 0 0 ch_in[29]
port 174 nsew signal input
flabel metal1 s 201150 11200 201206 12000 0 FreeSans 224 90 0 0 ch_in[2]
port 175 nsew signal input
flabel metal1 s 216382 11200 216438 12000 0 FreeSans 224 90 0 0 ch_in[30]
port 176 nsew signal input
flabel metal1 s 33802 0 33858 800 0 FreeSans 224 90 0 0 ch_in[31]
port 177 nsew signal input
flabel metal1 s 34890 0 34946 800 0 FreeSans 224 90 0 0 ch_in[32]
port 178 nsew signal input
flabel metal1 s 218014 11200 218070 12000 0 FreeSans 224 90 0 0 ch_in[33]
port 179 nsew signal input
flabel metal1 s 37066 0 37122 800 0 FreeSans 224 90 0 0 ch_in[34]
port 180 nsew signal input
flabel metal1 s 38154 0 38210 800 0 FreeSans 224 90 0 0 ch_in[35]
port 181 nsew signal input
flabel metal1 s 219646 11200 219702 12000 0 FreeSans 224 90 0 0 ch_in[36]
port 182 nsew signal input
flabel metal1 s 40330 0 40386 800 0 FreeSans 224 90 0 0 ch_in[37]
port 183 nsew signal input
flabel metal1 s 41418 0 41474 800 0 FreeSans 224 90 0 0 ch_in[38]
port 184 nsew signal input
flabel metal1 s 221278 11200 221334 12000 0 FreeSans 224 90 0 0 ch_in[39]
port 185 nsew signal input
flabel metal1 s 3338 0 3394 800 0 FreeSans 224 90 0 0 ch_in[3]
port 186 nsew signal input
flabel metal1 s 43594 0 43650 800 0 FreeSans 224 90 0 0 ch_in[40]
port 187 nsew signal input
flabel metal1 s 44682 0 44738 800 0 FreeSans 224 90 0 0 ch_in[41]
port 188 nsew signal input
flabel metal1 s 222910 11200 222966 12000 0 FreeSans 224 90 0 0 ch_in[42]
port 189 nsew signal input
flabel metal1 s 46858 0 46914 800 0 FreeSans 224 90 0 0 ch_in[43]
port 190 nsew signal input
flabel metal1 s 47946 0 48002 800 0 FreeSans 224 90 0 0 ch_in[44]
port 191 nsew signal input
flabel metal1 s 224542 11200 224598 12000 0 FreeSans 224 90 0 0 ch_in[45]
port 192 nsew signal input
flabel metal1 s 50122 0 50178 800 0 FreeSans 224 90 0 0 ch_in[46]
port 193 nsew signal input
flabel metal1 s 51210 0 51266 800 0 FreeSans 224 90 0 0 ch_in[47]
port 194 nsew signal input
flabel metal1 s 226174 11200 226230 12000 0 FreeSans 224 90 0 0 ch_in[48]
port 195 nsew signal input
flabel metal1 s 53386 0 53442 800 0 FreeSans 224 90 0 0 ch_in[49]
port 196 nsew signal input
flabel metal1 s 4426 0 4482 800 0 FreeSans 224 90 0 0 ch_in[4]
port 197 nsew signal input
flabel metal1 s 54474 0 54530 800 0 FreeSans 224 90 0 0 ch_in[50]
port 198 nsew signal input
flabel metal1 s 227806 11200 227862 12000 0 FreeSans 224 90 0 0 ch_in[51]
port 199 nsew signal input
flabel metal1 s 56650 0 56706 800 0 FreeSans 224 90 0 0 ch_in[52]
port 200 nsew signal input
flabel metal1 s 57738 0 57794 800 0 FreeSans 224 90 0 0 ch_in[53]
port 201 nsew signal input
flabel metal1 s 229438 11200 229494 12000 0 FreeSans 224 90 0 0 ch_in[54]
port 202 nsew signal input
flabel metal1 s 59914 0 59970 800 0 FreeSans 224 90 0 0 ch_in[55]
port 203 nsew signal input
flabel metal1 s 61002 0 61058 800 0 FreeSans 224 90 0 0 ch_in[56]
port 204 nsew signal input
flabel metal1 s 231070 11200 231126 12000 0 FreeSans 224 90 0 0 ch_in[57]
port 205 nsew signal input
flabel metal1 s 63178 0 63234 800 0 FreeSans 224 90 0 0 ch_in[58]
port 206 nsew signal input
flabel metal1 s 64266 0 64322 800 0 FreeSans 224 90 0 0 ch_in[59]
port 207 nsew signal input
flabel metal1 s 5514 0 5570 800 0 FreeSans 224 90 0 0 ch_in[5]
port 208 nsew signal input
flabel metal1 s 232702 11200 232758 12000 0 FreeSans 224 90 0 0 ch_in[60]
port 209 nsew signal input
flabel metal1 s 66442 0 66498 800 0 FreeSans 224 90 0 0 ch_in[61]
port 210 nsew signal input
flabel metal1 s 67530 0 67586 800 0 FreeSans 224 90 0 0 ch_in[62]
port 211 nsew signal input
flabel metal1 s 234334 11200 234390 12000 0 FreeSans 224 90 0 0 ch_in[63]
port 212 nsew signal input
flabel metal1 s 69706 0 69762 800 0 FreeSans 224 90 0 0 ch_in[64]
port 213 nsew signal input
flabel metal1 s 70794 0 70850 800 0 FreeSans 224 90 0 0 ch_in[65]
port 214 nsew signal input
flabel metal1 s 235966 11200 236022 12000 0 FreeSans 224 90 0 0 ch_in[66]
port 215 nsew signal input
flabel metal1 s 72970 0 73026 800 0 FreeSans 224 90 0 0 ch_in[67]
port 216 nsew signal input
flabel metal1 s 74058 0 74114 800 0 FreeSans 224 90 0 0 ch_in[68]
port 217 nsew signal input
flabel metal1 s 237598 11200 237654 12000 0 FreeSans 224 90 0 0 ch_in[69]
port 218 nsew signal input
flabel metal1 s 6602 0 6658 800 0 FreeSans 224 90 0 0 ch_in[6]
port 219 nsew signal input
flabel metal1 s 76234 0 76290 800 0 FreeSans 224 90 0 0 ch_in[70]
port 220 nsew signal input
flabel metal1 s 77322 0 77378 800 0 FreeSans 224 90 0 0 ch_in[71]
port 221 nsew signal input
flabel metal1 s 239230 11200 239286 12000 0 FreeSans 224 90 0 0 ch_in[72]
port 222 nsew signal input
flabel metal1 s 79498 0 79554 800 0 FreeSans 224 90 0 0 ch_in[73]
port 223 nsew signal input
flabel metal1 s 80586 0 80642 800 0 FreeSans 224 90 0 0 ch_in[74]
port 224 nsew signal input
flabel metal1 s 240862 11200 240918 12000 0 FreeSans 224 90 0 0 ch_in[75]
port 225 nsew signal input
flabel metal1 s 82762 0 82818 800 0 FreeSans 224 90 0 0 ch_in[76]
port 226 nsew signal input
flabel metal1 s 83850 0 83906 800 0 FreeSans 224 90 0 0 ch_in[77]
port 227 nsew signal input
flabel metal1 s 242494 11200 242550 12000 0 FreeSans 224 90 0 0 ch_in[78]
port 228 nsew signal input
flabel metal1 s 86026 0 86082 800 0 FreeSans 224 90 0 0 ch_in[79]
port 229 nsew signal input
flabel metal1 s 7690 0 7746 800 0 FreeSans 224 90 0 0 ch_in[7]
port 230 nsew signal input
flabel metal1 s 87114 0 87170 800 0 FreeSans 224 90 0 0 ch_in[80]
port 231 nsew signal input
flabel metal1 s 244126 11200 244182 12000 0 FreeSans 224 90 0 0 ch_in[81]
port 232 nsew signal input
flabel metal1 s 89290 0 89346 800 0 FreeSans 224 90 0 0 ch_in[82]
port 233 nsew signal input
flabel metal1 s 90378 0 90434 800 0 FreeSans 224 90 0 0 ch_in[83]
port 234 nsew signal input
flabel metal1 s 245758 11200 245814 12000 0 FreeSans 224 90 0 0 ch_in[84]
port 235 nsew signal input
flabel metal1 s 92554 0 92610 800 0 FreeSans 224 90 0 0 ch_in[85]
port 236 nsew signal input
flabel metal1 s 93642 0 93698 800 0 FreeSans 224 90 0 0 ch_in[86]
port 237 nsew signal input
flabel metal1 s 247390 11200 247446 12000 0 FreeSans 224 90 0 0 ch_in[87]
port 238 nsew signal input
flabel metal1 s 95818 0 95874 800 0 FreeSans 224 90 0 0 ch_in[88]
port 239 nsew signal input
flabel metal1 s 96906 0 96962 800 0 FreeSans 224 90 0 0 ch_in[89]
port 240 nsew signal input
flabel metal1 s 204414 11200 204470 12000 0 FreeSans 224 90 0 0 ch_in[8]
port 241 nsew signal input
flabel metal1 s 249022 11200 249078 12000 0 FreeSans 224 90 0 0 ch_in[90]
port 242 nsew signal input
flabel metal1 s 99082 0 99138 800 0 FreeSans 224 90 0 0 ch_in[91]
port 243 nsew signal input
flabel metal1 s 100170 0 100226 800 0 FreeSans 224 90 0 0 ch_in[92]
port 244 nsew signal input
flabel metal1 s 250654 11200 250710 12000 0 FreeSans 224 90 0 0 ch_in[93]
port 245 nsew signal input
flabel metal1 s 102346 0 102402 800 0 FreeSans 224 90 0 0 ch_in[94]
port 246 nsew signal input
flabel metal1 s 103434 0 103490 800 0 FreeSans 224 90 0 0 ch_in[95]
port 247 nsew signal input
flabel metal1 s 252286 11200 252342 12000 0 FreeSans 224 90 0 0 ch_in[96]
port 248 nsew signal input
flabel metal1 s 105610 0 105666 800 0 FreeSans 224 90 0 0 ch_in[97]
port 249 nsew signal input
flabel metal1 s 106698 0 106754 800 0 FreeSans 224 90 0 0 ch_in[98]
port 250 nsew signal input
flabel metal1 s 253918 11200 253974 12000 0 FreeSans 224 90 0 0 ch_in[99]
port 251 nsew signal input
flabel metal1 s 9866 0 9922 800 0 FreeSans 224 90 0 0 ch_in[9]
port 252 nsew signal input
flabel metal1 s 200062 11200 200118 12000 0 FreeSans 224 90 0 0 ch_out[0]
port 253 nsew signal tristate
flabel metal1 s 254462 11200 254518 12000 0 FreeSans 224 90 0 0 ch_out[100]
port 254 nsew signal tristate
flabel metal1 s 255006 11200 255062 12000 0 FreeSans 224 90 0 0 ch_out[101]
port 255 nsew signal tristate
flabel metal1 s 111050 0 111106 800 0 FreeSans 224 90 0 0 ch_out[102]
port 256 nsew signal tristate
flabel metal1 s 256094 11200 256150 12000 0 FreeSans 224 90 0 0 ch_out[103]
port 257 nsew signal tristate
flabel metal1 s 256638 11200 256694 12000 0 FreeSans 224 90 0 0 ch_out[104]
port 258 nsew signal tristate
flabel metal1 s 114314 0 114370 800 0 FreeSans 224 90 0 0 ch_out[105]
port 259 nsew signal tristate
flabel metal1 s 360066 11200 360122 12000 0 FreeSans 224 90 0 0 ch_out[106]
port 260 nsew signal tristate
flabel metal1 s 122202 0 122258 800 0 FreeSans 224 90 0 0 ch_out[107]
port 261 nsew signal tristate
flabel metal1 s 361154 11200 361210 12000 0 FreeSans 224 90 0 0 ch_out[108]
port 262 nsew signal tristate
flabel metal1 s 126554 0 126610 800 0 FreeSans 224 90 0 0 ch_out[109]
port 263 nsew signal tristate
flabel metal1 s 205502 11200 205558 12000 0 FreeSans 224 90 0 0 ch_out[10]
port 264 nsew signal tristate
flabel metal1 s 362242 11200 362298 12000 0 FreeSans 224 90 0 0 ch_out[110]
port 265 nsew signal tristate
flabel metal1 s 130906 0 130962 800 0 FreeSans 224 90 0 0 ch_out[111]
port 266 nsew signal tristate
flabel metal1 s 363330 11200 363386 12000 0 FreeSans 224 90 0 0 ch_out[112]
port 267 nsew signal tristate
flabel metal1 s 135258 0 135314 800 0 FreeSans 224 90 0 0 ch_out[113]
port 268 nsew signal tristate
flabel metal1 s 364418 11200 364474 12000 0 FreeSans 224 90 0 0 ch_out[114]
port 269 nsew signal tristate
flabel metal1 s 139610 0 139666 800 0 FreeSans 224 90 0 0 ch_out[115]
port 270 nsew signal tristate
flabel metal1 s 365506 11200 365562 12000 0 FreeSans 224 90 0 0 ch_out[116]
port 271 nsew signal tristate
flabel metal1 s 143962 0 144018 800 0 FreeSans 224 90 0 0 ch_out[117]
port 272 nsew signal tristate
flabel metal1 s 366594 11200 366650 12000 0 FreeSans 224 90 0 0 ch_out[118]
port 273 nsew signal tristate
flabel metal1 s 148314 0 148370 800 0 FreeSans 224 90 0 0 ch_out[119]
port 274 nsew signal tristate
flabel metal1 s 206046 11200 206102 12000 0 FreeSans 224 90 0 0 ch_out[11]
port 275 nsew signal tristate
flabel metal1 s 367682 11200 367738 12000 0 FreeSans 224 90 0 0 ch_out[120]
port 276 nsew signal tristate
flabel metal1 s 152666 0 152722 800 0 FreeSans 224 90 0 0 ch_out[121]
port 277 nsew signal tristate
flabel metal1 s 368770 11200 368826 12000 0 FreeSans 224 90 0 0 ch_out[122]
port 278 nsew signal tristate
flabel metal1 s 157018 0 157074 800 0 FreeSans 224 90 0 0 ch_out[123]
port 279 nsew signal tristate
flabel metal1 s 369858 11200 369914 12000 0 FreeSans 224 90 0 0 ch_out[124]
port 280 nsew signal tristate
flabel metal1 s 161370 0 161426 800 0 FreeSans 224 90 0 0 ch_out[125]
port 281 nsew signal tristate
flabel metal1 s 370946 11200 371002 12000 0 FreeSans 224 90 0 0 ch_out[126]
port 282 nsew signal tristate
flabel metal1 s 164226 0 164282 800 0 FreeSans 224 90 0 0 ch_out[127]
port 283 nsew signal tristate
flabel metal1 s 372034 11200 372090 12000 0 FreeSans 224 90 0 0 ch_out[128]
port 284 nsew signal tristate
flabel metal1 s 168578 0 168634 800 0 FreeSans 224 90 0 0 ch_out[129]
port 285 nsew signal tristate
flabel metal1 s 13130 0 13186 800 0 FreeSans 224 90 0 0 ch_out[12]
port 286 nsew signal tristate
flabel metal1 s 373122 11200 373178 12000 0 FreeSans 224 90 0 0 ch_out[130]
port 287 nsew signal tristate
flabel metal1 s 172930 0 172986 800 0 FreeSans 224 90 0 0 ch_out[131]
port 288 nsew signal tristate
flabel metal1 s 374210 11200 374266 12000 0 FreeSans 224 90 0 0 ch_out[132]
port 289 nsew signal tristate
flabel metal1 s 177282 0 177338 800 0 FreeSans 224 90 0 0 ch_out[133]
port 290 nsew signal tristate
flabel metal1 s 375298 11200 375354 12000 0 FreeSans 224 90 0 0 ch_out[134]
port 291 nsew signal tristate
flabel metal1 s 181634 0 181690 800 0 FreeSans 224 90 0 0 ch_out[135]
port 292 nsew signal tristate
flabel metal1 s 376386 11200 376442 12000 0 FreeSans 224 90 0 0 ch_out[136]
port 293 nsew signal tristate
flabel metal1 s 185986 0 186042 800 0 FreeSans 224 90 0 0 ch_out[137]
port 294 nsew signal tristate
flabel metal1 s 377474 11200 377530 12000 0 FreeSans 224 90 0 0 ch_out[138]
port 295 nsew signal tristate
flabel metal1 s 190338 0 190394 800 0 FreeSans 224 90 0 0 ch_out[139]
port 296 nsew signal tristate
flabel metal1 s 207134 11200 207190 12000 0 FreeSans 224 90 0 0 ch_out[13]
port 297 nsew signal tristate
flabel metal1 s 378562 11200 378618 12000 0 FreeSans 224 90 0 0 ch_out[140]
port 298 nsew signal tristate
flabel metal1 s 194690 0 194746 800 0 FreeSans 224 90 0 0 ch_out[141]
port 299 nsew signal tristate
flabel metal1 s 220054 0 220110 800 0 FreeSans 224 90 0 0 ch_out[142]
port 300 nsew signal tristate
flabel metal1 s 222230 0 222286 800 0 FreeSans 224 90 0 0 ch_out[143]
port 301 nsew signal tristate
flabel metal1 s 224406 0 224462 800 0 FreeSans 224 90 0 0 ch_out[144]
port 302 nsew signal tristate
flabel metal1 s 226582 0 226638 800 0 FreeSans 224 90 0 0 ch_out[145]
port 303 nsew signal tristate
flabel metal1 s 228758 0 228814 800 0 FreeSans 224 90 0 0 ch_out[146]
port 304 nsew signal tristate
flabel metal1 s 230934 0 230990 800 0 FreeSans 224 90 0 0 ch_out[147]
port 305 nsew signal tristate
flabel metal1 s 233110 0 233166 800 0 FreeSans 224 90 0 0 ch_out[148]
port 306 nsew signal tristate
flabel metal1 s 235286 0 235342 800 0 FreeSans 224 90 0 0 ch_out[149]
port 307 nsew signal tristate
flabel metal1 s 207678 11200 207734 12000 0 FreeSans 224 90 0 0 ch_out[14]
port 308 nsew signal tristate
flabel metal1 s 237462 0 237518 800 0 FreeSans 224 90 0 0 ch_out[150]
port 309 nsew signal tristate
flabel metal1 s 239638 0 239694 800 0 FreeSans 224 90 0 0 ch_out[151]
port 310 nsew signal tristate
flabel metal1 s 241814 0 241870 800 0 FreeSans 224 90 0 0 ch_out[152]
port 311 nsew signal tristate
flabel metal1 s 243990 0 244046 800 0 FreeSans 224 90 0 0 ch_out[153]
port 312 nsew signal tristate
flabel metal1 s 246166 0 246222 800 0 FreeSans 224 90 0 0 ch_out[154]
port 313 nsew signal tristate
flabel metal1 s 248342 0 248398 800 0 FreeSans 224 90 0 0 ch_out[155]
port 314 nsew signal tristate
flabel metal1 s 250518 0 250574 800 0 FreeSans 224 90 0 0 ch_out[156]
port 315 nsew signal tristate
flabel metal1 s 252694 0 252750 800 0 FreeSans 224 90 0 0 ch_out[157]
port 316 nsew signal tristate
flabel metal1 s 254870 0 254926 800 0 FreeSans 224 90 0 0 ch_out[158]
port 317 nsew signal tristate
flabel metal1 s 257046 0 257102 800 0 FreeSans 224 90 0 0 ch_out[159]
port 318 nsew signal tristate
flabel metal1 s 208222 11200 208278 12000 0 FreeSans 224 90 0 0 ch_out[15]
port 319 nsew signal tristate
flabel metal1 s 259222 0 259278 800 0 FreeSans 224 90 0 0 ch_out[160]
port 320 nsew signal tristate
flabel metal1 s 261398 0 261454 800 0 FreeSans 224 90 0 0 ch_out[161]
port 321 nsew signal tristate
flabel metal1 s 263574 0 263630 800 0 FreeSans 224 90 0 0 ch_out[162]
port 322 nsew signal tristate
flabel metal1 s 265750 0 265806 800 0 FreeSans 224 90 0 0 ch_out[163]
port 323 nsew signal tristate
flabel metal1 s 267926 0 267982 800 0 FreeSans 224 90 0 0 ch_out[164]
port 324 nsew signal tristate
flabel metal1 s 270102 0 270158 800 0 FreeSans 224 90 0 0 ch_out[165]
port 325 nsew signal tristate
flabel metal1 s 272278 0 272334 800 0 FreeSans 224 90 0 0 ch_out[166]
port 326 nsew signal tristate
flabel metal1 s 274454 0 274510 800 0 FreeSans 224 90 0 0 ch_out[167]
port 327 nsew signal tristate
flabel metal1 s 276630 0 276686 800 0 FreeSans 224 90 0 0 ch_out[168]
port 328 nsew signal tristate
flabel metal1 s 278806 0 278862 800 0 FreeSans 224 90 0 0 ch_out[169]
port 329 nsew signal tristate
flabel metal1 s 17482 0 17538 800 0 FreeSans 224 90 0 0 ch_out[16]
port 330 nsew signal tristate
flabel metal1 s 280982 0 281038 800 0 FreeSans 224 90 0 0 ch_out[170]
port 331 nsew signal tristate
flabel metal1 s 283158 0 283214 800 0 FreeSans 224 90 0 0 ch_out[171]
port 332 nsew signal tristate
flabel metal1 s 285334 0 285390 800 0 FreeSans 224 90 0 0 ch_out[172]
port 333 nsew signal tristate
flabel metal1 s 287510 0 287566 800 0 FreeSans 224 90 0 0 ch_out[173]
port 334 nsew signal tristate
flabel metal1 s 289686 0 289742 800 0 FreeSans 224 90 0 0 ch_out[174]
port 335 nsew signal tristate
flabel metal1 s 291862 0 291918 800 0 FreeSans 224 90 0 0 ch_out[175]
port 336 nsew signal tristate
flabel metal1 s 294038 0 294094 800 0 FreeSans 224 90 0 0 ch_out[176]
port 337 nsew signal tristate
flabel metal1 s 296214 0 296270 800 0 FreeSans 224 90 0 0 ch_out[177]
port 338 nsew signal tristate
flabel metal1 s 298390 0 298446 800 0 FreeSans 224 90 0 0 ch_out[178]
port 339 nsew signal tristate
flabel metal1 s 300566 0 300622 800 0 FreeSans 224 90 0 0 ch_out[179]
port 340 nsew signal tristate
flabel metal1 s 209310 11200 209366 12000 0 FreeSans 224 90 0 0 ch_out[17]
port 341 nsew signal tristate
flabel metal1 s 302742 0 302798 800 0 FreeSans 224 90 0 0 ch_out[180]
port 342 nsew signal tristate
flabel metal1 s 304918 0 304974 800 0 FreeSans 224 90 0 0 ch_out[181]
port 343 nsew signal tristate
flabel metal1 s 307094 0 307150 800 0 FreeSans 224 90 0 0 ch_out[182]
port 344 nsew signal tristate
flabel metal1 s 309270 0 309326 800 0 FreeSans 224 90 0 0 ch_out[183]
port 345 nsew signal tristate
flabel metal1 s 311446 0 311502 800 0 FreeSans 224 90 0 0 ch_out[184]
port 346 nsew signal tristate
flabel metal1 s 313622 0 313678 800 0 FreeSans 224 90 0 0 ch_out[185]
port 347 nsew signal tristate
flabel metal1 s 315798 0 315854 800 0 FreeSans 224 90 0 0 ch_out[186]
port 348 nsew signal tristate
flabel metal1 s 317974 0 318030 800 0 FreeSans 224 90 0 0 ch_out[187]
port 349 nsew signal tristate
flabel metal1 s 360066 0 360122 800 0 FreeSans 224 90 0 0 ch_out[188]
port 350 nsew signal tristate
flabel metal1 s 362242 0 362298 800 0 FreeSans 224 90 0 0 ch_out[189]
port 351 nsew signal tristate
flabel metal1 s 209854 11200 209910 12000 0 FreeSans 224 90 0 0 ch_out[18]
port 352 nsew signal tristate
flabel metal1 s 364418 0 364474 800 0 FreeSans 224 90 0 0 ch_out[190]
port 353 nsew signal tristate
flabel metal1 s 366594 0 366650 800 0 FreeSans 224 90 0 0 ch_out[191]
port 354 nsew signal tristate
flabel metal1 s 368770 0 368826 800 0 FreeSans 224 90 0 0 ch_out[192]
port 355 nsew signal tristate
flabel metal1 s 370946 0 371002 800 0 FreeSans 224 90 0 0 ch_out[193]
port 356 nsew signal tristate
flabel metal1 s 373122 0 373178 800 0 FreeSans 224 90 0 0 ch_out[194]
port 357 nsew signal tristate
flabel metal1 s 375298 0 375354 800 0 FreeSans 224 90 0 0 ch_out[195]
port 358 nsew signal tristate
flabel metal1 s 377474 0 377530 800 0 FreeSans 224 90 0 0 ch_out[196]
port 359 nsew signal tristate
flabel metal1 s 379650 0 379706 800 0 FreeSans 224 90 0 0 ch_out[197]
port 360 nsew signal tristate
flabel metal1 s 381826 0 381882 800 0 FreeSans 224 90 0 0 ch_out[198]
port 361 nsew signal tristate
flabel metal1 s 384002 0 384058 800 0 FreeSans 224 90 0 0 ch_out[199]
port 362 nsew signal tristate
flabel metal1 s 210398 11200 210454 12000 0 FreeSans 224 90 0 0 ch_out[19]
port 363 nsew signal tristate
flabel metal1 s 200606 11200 200662 12000 0 FreeSans 224 90 0 0 ch_out[1]
port 364 nsew signal tristate
flabel metal1 s 386178 0 386234 800 0 FreeSans 224 90 0 0 ch_out[200]
port 365 nsew signal tristate
flabel metal1 s 388354 0 388410 800 0 FreeSans 224 90 0 0 ch_out[201]
port 366 nsew signal tristate
flabel metal1 s 390530 0 390586 800 0 FreeSans 224 90 0 0 ch_out[202]
port 367 nsew signal tristate
flabel metal1 s 392706 0 392762 800 0 FreeSans 224 90 0 0 ch_out[203]
port 368 nsew signal tristate
flabel metal1 s 394882 0 394938 800 0 FreeSans 224 90 0 0 ch_out[204]
port 369 nsew signal tristate
flabel metal1 s 397058 0 397114 800 0 FreeSans 224 90 0 0 ch_out[205]
port 370 nsew signal tristate
flabel metal1 s 399234 0 399290 800 0 FreeSans 224 90 0 0 ch_out[206]
port 371 nsew signal tristate
flabel metal1 s 401410 0 401466 800 0 FreeSans 224 90 0 0 ch_out[207]
port 372 nsew signal tristate
flabel metal1 s 403586 0 403642 800 0 FreeSans 224 90 0 0 ch_out[208]
port 373 nsew signal tristate
flabel metal1 s 405762 0 405818 800 0 FreeSans 224 90 0 0 ch_out[209]
port 374 nsew signal tristate
flabel metal1 s 21834 0 21890 800 0 FreeSans 224 90 0 0 ch_out[20]
port 375 nsew signal tristate
flabel metal1 s 407938 0 407994 800 0 FreeSans 224 90 0 0 ch_out[210]
port 376 nsew signal tristate
flabel metal1 s 410114 0 410170 800 0 FreeSans 224 90 0 0 ch_out[211]
port 377 nsew signal tristate
flabel metal1 s 412290 0 412346 800 0 FreeSans 224 90 0 0 ch_out[212]
port 378 nsew signal tristate
flabel metal1 s 414466 0 414522 800 0 FreeSans 224 90 0 0 ch_out[213]
port 379 nsew signal tristate
flabel metal1 s 416642 0 416698 800 0 FreeSans 224 90 0 0 ch_out[214]
port 380 nsew signal tristate
flabel metal1 s 418818 0 418874 800 0 FreeSans 224 90 0 0 ch_out[215]
port 381 nsew signal tristate
flabel metal1 s 420994 0 421050 800 0 FreeSans 224 90 0 0 ch_out[216]
port 382 nsew signal tristate
flabel metal1 s 423170 0 423226 800 0 FreeSans 224 90 0 0 ch_out[217]
port 383 nsew signal tristate
flabel metal1 s 425346 0 425402 800 0 FreeSans 224 90 0 0 ch_out[218]
port 384 nsew signal tristate
flabel metal1 s 427522 0 427578 800 0 FreeSans 224 90 0 0 ch_out[219]
port 385 nsew signal tristate
flabel metal1 s 211486 11200 211542 12000 0 FreeSans 224 90 0 0 ch_out[21]
port 386 nsew signal tristate
flabel metal1 s 429698 0 429754 800 0 FreeSans 224 90 0 0 ch_out[220]
port 387 nsew signal tristate
flabel metal1 s 431874 0 431930 800 0 FreeSans 224 90 0 0 ch_out[221]
port 388 nsew signal tristate
flabel metal1 s 434050 0 434106 800 0 FreeSans 224 90 0 0 ch_out[222]
port 389 nsew signal tristate
flabel metal1 s 436226 0 436282 800 0 FreeSans 224 90 0 0 ch_out[223]
port 390 nsew signal tristate
flabel metal1 s 438402 0 438458 800 0 FreeSans 224 90 0 0 ch_out[224]
port 391 nsew signal tristate
flabel metal1 s 440578 0 440634 800 0 FreeSans 224 90 0 0 ch_out[225]
port 392 nsew signal tristate
flabel metal1 s 442754 0 442810 800 0 FreeSans 224 90 0 0 ch_out[226]
port 393 nsew signal tristate
flabel metal1 s 444930 0 444986 800 0 FreeSans 224 90 0 0 ch_out[227]
port 394 nsew signal tristate
flabel metal1 s 447106 0 447162 800 0 FreeSans 224 90 0 0 ch_out[228]
port 395 nsew signal tristate
flabel metal1 s 449282 0 449338 800 0 FreeSans 224 90 0 0 ch_out[229]
port 396 nsew signal tristate
flabel metal1 s 212030 11200 212086 12000 0 FreeSans 224 90 0 0 ch_out[22]
port 397 nsew signal tristate
flabel metal1 s 451458 0 451514 800 0 FreeSans 224 90 0 0 ch_out[230]
port 398 nsew signal tristate
flabel metal1 s 453634 0 453690 800 0 FreeSans 224 90 0 0 ch_out[231]
port 399 nsew signal tristate
flabel metal1 s 455810 0 455866 800 0 FreeSans 224 90 0 0 ch_out[232]
port 400 nsew signal tristate
flabel metal1 s 457986 0 458042 800 0 FreeSans 224 90 0 0 ch_out[233]
port 401 nsew signal tristate
flabel metal1 s 460162 0 460218 800 0 FreeSans 224 90 0 0 ch_out[234]
port 402 nsew signal tristate
flabel metal1 s 462338 0 462394 800 0 FreeSans 224 90 0 0 ch_out[235]
port 403 nsew signal tristate
flabel metal1 s 464514 0 464570 800 0 FreeSans 224 90 0 0 ch_out[236]
port 404 nsew signal tristate
flabel metal1 s 466690 0 466746 800 0 FreeSans 224 90 0 0 ch_out[237]
port 405 nsew signal tristate
flabel metal1 s 468866 0 468922 800 0 FreeSans 224 90 0 0 ch_out[238]
port 406 nsew signal tristate
flabel metal1 s 471042 0 471098 800 0 FreeSans 224 90 0 0 ch_out[239]
port 407 nsew signal tristate
flabel metal1 s 212574 11200 212630 12000 0 FreeSans 224 90 0 0 ch_out[23]
port 408 nsew signal tristate
flabel metal1 s 473218 0 473274 800 0 FreeSans 224 90 0 0 ch_out[240]
port 409 nsew signal tristate
flabel metal1 s 475394 0 475450 800 0 FreeSans 224 90 0 0 ch_out[241]
port 410 nsew signal tristate
flabel metal1 s 477570 0 477626 800 0 FreeSans 224 90 0 0 ch_out[242]
port 411 nsew signal tristate
flabel metal1 s 479746 0 479802 800 0 FreeSans 224 90 0 0 ch_out[243]
port 412 nsew signal tristate
flabel metal1 s 481922 0 481978 800 0 FreeSans 224 90 0 0 ch_out[244]
port 413 nsew signal tristate
flabel metal1 s 484098 0 484154 800 0 FreeSans 224 90 0 0 ch_out[245]
port 414 nsew signal tristate
flabel metal1 s 486274 0 486330 800 0 FreeSans 224 90 0 0 ch_out[246]
port 415 nsew signal tristate
flabel metal1 s 488450 0 488506 800 0 FreeSans 224 90 0 0 ch_out[247]
port 416 nsew signal tristate
flabel metal1 s 490626 0 490682 800 0 FreeSans 224 90 0 0 ch_out[248]
port 417 nsew signal tristate
flabel metal1 s 492802 0 492858 800 0 FreeSans 224 90 0 0 ch_out[249]
port 418 nsew signal tristate
flabel metal1 s 26186 0 26242 800 0 FreeSans 224 90 0 0 ch_out[24]
port 419 nsew signal tristate
flabel metal1 s 494978 0 495034 800 0 FreeSans 224 90 0 0 ch_out[250]
port 420 nsew signal tristate
flabel metal1 s 497154 0 497210 800 0 FreeSans 224 90 0 0 ch_out[251]
port 421 nsew signal tristate
flabel metal1 s 488722 11200 488778 12000 0 FreeSans 224 90 0 0 ch_out[252]
port 422 nsew signal tristate
flabel metal1 s 213662 11200 213718 12000 0 FreeSans 224 90 0 0 ch_out[25]
port 423 nsew signal tristate
flabel metal1 s 214206 11200 214262 12000 0 FreeSans 224 90 0 0 ch_out[26]
port 424 nsew signal tristate
flabel metal1 s 29450 0 29506 800 0 FreeSans 224 90 0 0 ch_out[27]
port 425 nsew signal tristate
flabel metal1 s 215294 11200 215350 12000 0 FreeSans 224 90 0 0 ch_out[28]
port 426 nsew signal tristate
flabel metal1 s 215838 11200 215894 12000 0 FreeSans 224 90 0 0 ch_out[29]
port 427 nsew signal tristate
flabel metal1 s 2250 0 2306 800 0 FreeSans 224 90 0 0 ch_out[2]
port 428 nsew signal tristate
flabel metal1 s 32714 0 32770 800 0 FreeSans 224 90 0 0 ch_out[30]
port 429 nsew signal tristate
flabel metal1 s 216926 11200 216982 12000 0 FreeSans 224 90 0 0 ch_out[31]
port 430 nsew signal tristate
flabel metal1 s 217470 11200 217526 12000 0 FreeSans 224 90 0 0 ch_out[32]
port 431 nsew signal tristate
flabel metal1 s 35978 0 36034 800 0 FreeSans 224 90 0 0 ch_out[33]
port 432 nsew signal tristate
flabel metal1 s 218558 11200 218614 12000 0 FreeSans 224 90 0 0 ch_out[34]
port 433 nsew signal tristate
flabel metal1 s 219102 11200 219158 12000 0 FreeSans 224 90 0 0 ch_out[35]
port 434 nsew signal tristate
flabel metal1 s 39242 0 39298 800 0 FreeSans 224 90 0 0 ch_out[36]
port 435 nsew signal tristate
flabel metal1 s 220190 11200 220246 12000 0 FreeSans 224 90 0 0 ch_out[37]
port 436 nsew signal tristate
flabel metal1 s 220734 11200 220790 12000 0 FreeSans 224 90 0 0 ch_out[38]
port 437 nsew signal tristate
flabel metal1 s 42506 0 42562 800 0 FreeSans 224 90 0 0 ch_out[39]
port 438 nsew signal tristate
flabel metal1 s 201694 11200 201750 12000 0 FreeSans 224 90 0 0 ch_out[3]
port 439 nsew signal tristate
flabel metal1 s 221822 11200 221878 12000 0 FreeSans 224 90 0 0 ch_out[40]
port 440 nsew signal tristate
flabel metal1 s 222366 11200 222422 12000 0 FreeSans 224 90 0 0 ch_out[41]
port 441 nsew signal tristate
flabel metal1 s 45770 0 45826 800 0 FreeSans 224 90 0 0 ch_out[42]
port 442 nsew signal tristate
flabel metal1 s 223454 11200 223510 12000 0 FreeSans 224 90 0 0 ch_out[43]
port 443 nsew signal tristate
flabel metal1 s 223998 11200 224054 12000 0 FreeSans 224 90 0 0 ch_out[44]
port 444 nsew signal tristate
flabel metal1 s 49034 0 49090 800 0 FreeSans 224 90 0 0 ch_out[45]
port 445 nsew signal tristate
flabel metal1 s 225086 11200 225142 12000 0 FreeSans 224 90 0 0 ch_out[46]
port 446 nsew signal tristate
flabel metal1 s 225630 11200 225686 12000 0 FreeSans 224 90 0 0 ch_out[47]
port 447 nsew signal tristate
flabel metal1 s 52298 0 52354 800 0 FreeSans 224 90 0 0 ch_out[48]
port 448 nsew signal tristate
flabel metal1 s 226718 11200 226774 12000 0 FreeSans 224 90 0 0 ch_out[49]
port 449 nsew signal tristate
flabel metal1 s 202238 11200 202294 12000 0 FreeSans 224 90 0 0 ch_out[4]
port 450 nsew signal tristate
flabel metal1 s 227262 11200 227318 12000 0 FreeSans 224 90 0 0 ch_out[50]
port 451 nsew signal tristate
flabel metal1 s 55562 0 55618 800 0 FreeSans 224 90 0 0 ch_out[51]
port 452 nsew signal tristate
flabel metal1 s 228350 11200 228406 12000 0 FreeSans 224 90 0 0 ch_out[52]
port 453 nsew signal tristate
flabel metal1 s 228894 11200 228950 12000 0 FreeSans 224 90 0 0 ch_out[53]
port 454 nsew signal tristate
flabel metal1 s 58826 0 58882 800 0 FreeSans 224 90 0 0 ch_out[54]
port 455 nsew signal tristate
flabel metal1 s 229982 11200 230038 12000 0 FreeSans 224 90 0 0 ch_out[55]
port 456 nsew signal tristate
flabel metal1 s 230526 11200 230582 12000 0 FreeSans 224 90 0 0 ch_out[56]
port 457 nsew signal tristate
flabel metal1 s 62090 0 62146 800 0 FreeSans 224 90 0 0 ch_out[57]
port 458 nsew signal tristate
flabel metal1 s 231614 11200 231670 12000 0 FreeSans 224 90 0 0 ch_out[58]
port 459 nsew signal tristate
flabel metal1 s 232158 11200 232214 12000 0 FreeSans 224 90 0 0 ch_out[59]
port 460 nsew signal tristate
flabel metal1 s 202782 11200 202838 12000 0 FreeSans 224 90 0 0 ch_out[5]
port 461 nsew signal tristate
flabel metal1 s 65354 0 65410 800 0 FreeSans 224 90 0 0 ch_out[60]
port 462 nsew signal tristate
flabel metal1 s 233246 11200 233302 12000 0 FreeSans 224 90 0 0 ch_out[61]
port 463 nsew signal tristate
flabel metal1 s 233790 11200 233846 12000 0 FreeSans 224 90 0 0 ch_out[62]
port 464 nsew signal tristate
flabel metal1 s 68618 0 68674 800 0 FreeSans 224 90 0 0 ch_out[63]
port 465 nsew signal tristate
flabel metal1 s 234878 11200 234934 12000 0 FreeSans 224 90 0 0 ch_out[64]
port 466 nsew signal tristate
flabel metal1 s 235422 11200 235478 12000 0 FreeSans 224 90 0 0 ch_out[65]
port 467 nsew signal tristate
flabel metal1 s 71882 0 71938 800 0 FreeSans 224 90 0 0 ch_out[66]
port 468 nsew signal tristate
flabel metal1 s 236510 11200 236566 12000 0 FreeSans 224 90 0 0 ch_out[67]
port 469 nsew signal tristate
flabel metal1 s 237054 11200 237110 12000 0 FreeSans 224 90 0 0 ch_out[68]
port 470 nsew signal tristate
flabel metal1 s 75146 0 75202 800 0 FreeSans 224 90 0 0 ch_out[69]
port 471 nsew signal tristate
flabel metal1 s 203326 11200 203382 12000 0 FreeSans 224 90 0 0 ch_out[6]
port 472 nsew signal tristate
flabel metal1 s 238142 11200 238198 12000 0 FreeSans 224 90 0 0 ch_out[70]
port 473 nsew signal tristate
flabel metal1 s 238686 11200 238742 12000 0 FreeSans 224 90 0 0 ch_out[71]
port 474 nsew signal tristate
flabel metal1 s 78410 0 78466 800 0 FreeSans 224 90 0 0 ch_out[72]
port 475 nsew signal tristate
flabel metal1 s 239774 11200 239830 12000 0 FreeSans 224 90 0 0 ch_out[73]
port 476 nsew signal tristate
flabel metal1 s 240318 11200 240374 12000 0 FreeSans 224 90 0 0 ch_out[74]
port 477 nsew signal tristate
flabel metal1 s 81674 0 81730 800 0 FreeSans 224 90 0 0 ch_out[75]
port 478 nsew signal tristate
flabel metal1 s 241406 11200 241462 12000 0 FreeSans 224 90 0 0 ch_out[76]
port 479 nsew signal tristate
flabel metal1 s 241950 11200 242006 12000 0 FreeSans 224 90 0 0 ch_out[77]
port 480 nsew signal tristate
flabel metal1 s 84938 0 84994 800 0 FreeSans 224 90 0 0 ch_out[78]
port 481 nsew signal tristate
flabel metal1 s 243038 11200 243094 12000 0 FreeSans 224 90 0 0 ch_out[79]
port 482 nsew signal tristate
flabel metal1 s 203870 11200 203926 12000 0 FreeSans 224 90 0 0 ch_out[7]
port 483 nsew signal tristate
flabel metal1 s 243582 11200 243638 12000 0 FreeSans 224 90 0 0 ch_out[80]
port 484 nsew signal tristate
flabel metal1 s 88202 0 88258 800 0 FreeSans 224 90 0 0 ch_out[81]
port 485 nsew signal tristate
flabel metal1 s 244670 11200 244726 12000 0 FreeSans 224 90 0 0 ch_out[82]
port 486 nsew signal tristate
flabel metal1 s 245214 11200 245270 12000 0 FreeSans 224 90 0 0 ch_out[83]
port 487 nsew signal tristate
flabel metal1 s 91466 0 91522 800 0 FreeSans 224 90 0 0 ch_out[84]
port 488 nsew signal tristate
flabel metal1 s 246302 11200 246358 12000 0 FreeSans 224 90 0 0 ch_out[85]
port 489 nsew signal tristate
flabel metal1 s 246846 11200 246902 12000 0 FreeSans 224 90 0 0 ch_out[86]
port 490 nsew signal tristate
flabel metal1 s 94730 0 94786 800 0 FreeSans 224 90 0 0 ch_out[87]
port 491 nsew signal tristate
flabel metal1 s 247934 11200 247990 12000 0 FreeSans 224 90 0 0 ch_out[88]
port 492 nsew signal tristate
flabel metal1 s 248478 11200 248534 12000 0 FreeSans 224 90 0 0 ch_out[89]
port 493 nsew signal tristate
flabel metal1 s 8778 0 8834 800 0 FreeSans 224 90 0 0 ch_out[8]
port 494 nsew signal tristate
flabel metal1 s 97994 0 98050 800 0 FreeSans 224 90 0 0 ch_out[90]
port 495 nsew signal tristate
flabel metal1 s 249566 11200 249622 12000 0 FreeSans 224 90 0 0 ch_out[91]
port 496 nsew signal tristate
flabel metal1 s 250110 11200 250166 12000 0 FreeSans 224 90 0 0 ch_out[92]
port 497 nsew signal tristate
flabel metal1 s 101258 0 101314 800 0 FreeSans 224 90 0 0 ch_out[93]
port 498 nsew signal tristate
flabel metal1 s 251198 11200 251254 12000 0 FreeSans 224 90 0 0 ch_out[94]
port 499 nsew signal tristate
flabel metal1 s 251742 11200 251798 12000 0 FreeSans 224 90 0 0 ch_out[95]
port 500 nsew signal tristate
flabel metal1 s 104522 0 104578 800 0 FreeSans 224 90 0 0 ch_out[96]
port 501 nsew signal tristate
flabel metal1 s 252830 11200 252886 12000 0 FreeSans 224 90 0 0 ch_out[97]
port 502 nsew signal tristate
flabel metal1 s 253374 11200 253430 12000 0 FreeSans 224 90 0 0 ch_out[98]
port 503 nsew signal tristate
flabel metal1 s 107786 0 107842 800 0 FreeSans 224 90 0 0 ch_out[99]
port 504 nsew signal tristate
flabel metal1 s 204958 11200 205014 12000 0 FreeSans 224 90 0 0 ch_out[9]
port 505 nsew signal tristate
flabel metal2 s -416 656 -96 11312 0 FreeSans 1792 90 0 0 vccd1
port 506 nsew power bidirectional
flabel metal3 s -416 656 530336 976 0 FreeSans 1920 0 0 0 vccd1
port 506 nsew power bidirectional
flabel metal3 s -416 10992 530336 11312 0 FreeSans 1920 0 0 0 vccd1
port 506 nsew power bidirectional
flabel metal2 s 530016 656 530336 11312 0 FreeSans 1792 90 0 0 vccd1
port 506 nsew power bidirectional
flabel metal2 s 66908 -4 67228 11972 0 FreeSans 1792 90 0 0 vccd1
port 506 nsew power bidirectional
flabel metal2 s 198836 -4 199156 11972 0 FreeSans 1792 90 0 0 vccd1
port 506 nsew power bidirectional
flabel metal2 s 330764 -4 331084 11972 0 FreeSans 1792 90 0 0 vccd1
port 506 nsew power bidirectional
flabel metal2 s 462692 -4 463012 11972 0 FreeSans 1792 90 0 0 vccd1
port 506 nsew power bidirectional
flabel metal3 s -1076 2968 530996 3288 0 FreeSans 1920 0 0 0 vccd1
port 506 nsew power bidirectional
flabel metal3 s -1076 4872 530996 5192 0 FreeSans 1920 0 0 0 vccd1
port 506 nsew power bidirectional
flabel metal3 s -1076 6776 530996 7096 0 FreeSans 1920 0 0 0 vccd1
port 506 nsew power bidirectional
flabel metal3 s -1076 8680 530996 9000 0 FreeSans 1920 0 0 0 vccd1
port 506 nsew power bidirectional
flabel metal2 s -1076 -4 -756 11972 0 FreeSans 1792 90 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal3 s -1076 -4 530996 316 0 FreeSans 1920 0 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal3 s -1076 11652 530996 11972 0 FreeSans 1920 0 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal2 s 530676 -4 530996 11972 0 FreeSans 1792 90 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal2 s 67568 -4 67888 11972 0 FreeSans 1792 90 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal2 s 199496 -4 199816 11972 0 FreeSans 1792 90 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal2 s 331424 -4 331744 11972 0 FreeSans 1792 90 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal2 s 463352 -4 463672 11972 0 FreeSans 1792 90 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal3 s -1076 3628 530996 3948 0 FreeSans 1920 0 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal3 s -1076 5532 530996 5852 0 FreeSans 1920 0 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal3 s -1076 7436 530996 7756 0 FreeSans 1920 0 0 0 vssd1
port 507 nsew ground bidirectional
flabel metal3 s -1076 9340 530996 9660 0 FreeSans 1920 0 0 0 vssd1
port 507 nsew ground bidirectional
rlabel metal1 264960 9248 264960 9248 0 vccd1
rlabel metal1 264960 9792 264960 9792 0 vssd1
rlabel metal1 1426 2346 1426 2346 0 ch_in[0]
rlabel metal2 130686 2210 130686 2210 0 ch_in[100]
rlabel metal2 118634 1513 118634 1513 0 ch_in[101]
rlabel metal2 251206 9860 251206 9860 0 ch_in[102]
rlabel metal1 132894 3502 132894 3502 0 ch_in[103]
rlabel metal1 113650 646 113650 646 0 ch_in[104]
rlabel metal2 255714 10234 255714 10234 0 ch_in[105]
rlabel metal2 130778 1071 130778 1071 0 ch_in[106]
rlabel metal2 252586 5984 252586 5984 0 ch_in[107]
rlabel via1 137770 1173 137770 1173 0 ch_in[108]
rlabel metal2 257002 8976 257002 8976 0 ch_in[109]
rlabel metal1 12236 2346 12236 2346 0 ch_in[10]
rlabel metal1 137862 1224 137862 1224 0 ch_in[110]
rlabel metal2 262062 9248 262062 9248 0 ch_in[111]
rlabel metal1 134028 782 134028 782 0 ch_in[112]
rlabel metal2 267122 9214 267122 9214 0 ch_in[113]
rlabel via1 139334 595 139334 595 0 ch_in[114]
rlabel metal2 272182 9180 272182 9180 0 ch_in[115]
rlabel metal2 147982 119 147982 119 0 ch_in[116]
rlabel metal2 277150 9860 277150 9860 0 ch_in[117]
rlabel metal1 168912 2346 168912 2346 0 ch_in[118]
rlabel metal2 282302 9384 282302 9384 0 ch_in[119]
rlabel metal2 14306 1972 14306 1972 0 ch_in[11]
rlabel metal1 151462 714 151462 714 0 ch_in[120]
rlabel metal2 287454 9350 287454 9350 0 ch_in[121]
rlabel metal1 178618 2822 178618 2822 0 ch_in[122]
rlabel metal2 292606 9316 292606 9316 0 ch_in[123]
rlabel metal1 183954 2822 183954 2822 0 ch_in[124]
rlabel metal2 297758 9180 297758 9180 0 ch_in[125]
rlabel metal1 189290 2822 189290 2822 0 ch_in[126]
rlabel metal2 302450 9520 302450 9520 0 ch_in[127]
rlabel metal1 194902 2890 194902 2890 0 ch_in[128]
rlabel metal2 307510 9486 307510 9486 0 ch_in[129]
rlabel metal2 206218 10829 206218 10829 0 ch_in[12]
rlabel via1 200077 2414 200077 2414 0 ch_in[130]
rlabel metal2 312478 9452 312478 9452 0 ch_in[131]
rlabel metal1 205344 2414 205344 2414 0 ch_in[132]
rlabel metal2 317538 9350 317538 9350 0 ch_in[133]
rlabel metal1 210496 2414 210496 2414 0 ch_in[134]
rlabel metal2 322506 9554 322506 9554 0 ch_in[135]
rlabel metal1 215648 2414 215648 2414 0 ch_in[136]
rlabel metal1 327244 8942 327244 8942 0 ch_in[137]
rlabel metal1 220800 2414 220800 2414 0 ch_in[138]
rlabel metal2 332534 9520 332534 9520 0 ch_in[139]
rlabel metal2 16606 2142 16606 2142 0 ch_in[13]
rlabel metal2 219650 1088 219650 1088 0 ch_in[140]
rlabel metal2 337502 9486 337502 9486 0 ch_in[141]
rlabel metal2 340170 9792 340170 9792 0 ch_in[142]
rlabel metal2 342746 10404 342746 10404 0 ch_in[143]
rlabel metal1 345161 9622 345161 9622 0 ch_in[144]
rlabel metal2 347622 10438 347622 10438 0 ch_in[145]
rlabel metal2 350106 8942 350106 8942 0 ch_in[146]
rlabel metal2 382122 10472 382122 10472 0 ch_in[147]
rlabel metal2 364182 9860 364182 9860 0 ch_in[148]
rlabel metal2 383226 10812 383226 10812 0 ch_in[149]
rlabel metal1 19412 2346 19412 2346 0 ch_in[14]
rlabel metal2 380006 10030 380006 10030 0 ch_in[150]
rlabel metal2 362158 9180 362158 9180 0 ch_in[151]
rlabel metal1 365608 9486 365608 9486 0 ch_in[152]
rlabel metal2 367310 8942 367310 8942 0 ch_in[153]
rlabel metal2 382214 9962 382214 9962 0 ch_in[154]
rlabel metal2 382950 9520 382950 9520 0 ch_in[155]
rlabel metal2 385894 10098 385894 10098 0 ch_in[156]
rlabel metal2 388010 10200 388010 10200 0 ch_in[157]
rlabel metal2 387090 9860 387090 9860 0 ch_in[158]
rlabel metal1 383732 9418 383732 9418 0 ch_in[159]
rlabel metal1 19366 2822 19366 2822 0 ch_in[15]
rlabel metal1 386538 9622 386538 9622 0 ch_in[160]
rlabel metal1 280554 2414 280554 2414 0 ch_in[161]
rlabel metal2 283406 2516 283406 2516 0 ch_in[162]
rlabel metal1 285706 2414 285706 2414 0 ch_in[163]
rlabel metal1 288282 2414 288282 2414 0 ch_in[164]
rlabel metal1 290858 2414 290858 2414 0 ch_in[165]
rlabel metal1 293434 2414 293434 2414 0 ch_in[166]
rlabel metal2 364734 5644 364734 5644 0 ch_in[167]
rlabel metal1 298586 2414 298586 2414 0 ch_in[168]
rlabel metal1 301162 2414 301162 2414 0 ch_in[169]
rlabel metal2 189198 5270 189198 5270 0 ch_in[16]
rlabel metal1 303738 2414 303738 2414 0 ch_in[170]
rlabel metal1 306314 2414 306314 2414 0 ch_in[171]
rlabel metal1 308890 2414 308890 2414 0 ch_in[172]
rlabel metal1 349738 2414 349738 2414 0 ch_in[173]
rlabel metal2 361606 4182 361606 4182 0 ch_in[174]
rlabel metal1 318090 2618 318090 2618 0 ch_in[175]
rlabel metal2 367954 3944 367954 3944 0 ch_in[176]
rlabel metal2 322046 3604 322046 3604 0 ch_in[177]
rlabel metal2 324622 1904 324622 1904 0 ch_in[178]
rlabel metal1 326922 2414 326922 2414 0 ch_in[179]
rlabel metal2 21666 2278 21666 2278 0 ch_in[17]
rlabel metal2 329774 2108 329774 2108 0 ch_in[180]
rlabel metal2 332350 1836 332350 1836 0 ch_in[181]
rlabel metal2 334926 3536 334926 3536 0 ch_in[182]
rlabel metal2 337502 2006 337502 2006 0 ch_in[183]
rlabel metal2 340078 2176 340078 2176 0 ch_in[184]
rlabel via1 403084 10982 403084 10982 0 ch_in[185]
rlabel metal2 345230 1938 345230 1938 0 ch_in[186]
rlabel metal1 348450 2550 348450 2550 0 ch_in[187]
rlabel via2 350382 2363 350382 2363 0 ch_in[188]
rlabel via2 352958 2499 352958 2499 0 ch_in[189]
rlabel metal1 19688 1020 19688 1020 0 ch_in[18]
rlabel metal1 355258 2414 355258 2414 0 ch_in[190]
rlabel metal2 358110 2074 358110 2074 0 ch_in[191]
rlabel metal2 360686 2516 360686 2516 0 ch_in[192]
rlabel metal1 393300 2312 393300 2312 0 ch_in[193]
rlabel metal2 441646 8568 441646 8568 0 ch_in[194]
rlabel metal2 400430 3400 400430 3400 0 ch_in[195]
rlabel metal2 442106 7242 442106 7242 0 ch_in[196]
rlabel metal1 398130 2448 398130 2448 0 ch_in[197]
rlabel metal2 442658 8636 442658 8636 0 ch_in[198]
rlabel metal2 383778 2108 383778 2108 0 ch_in[199]
rlabel metal1 24242 2822 24242 2822 0 ch_in[19]
rlabel metal1 1472 2822 1472 2822 0 ch_in[1]
rlabel metal2 381294 1904 381294 1904 0 ch_in[200]
rlabel metal1 383916 2278 383916 2278 0 ch_in[201]
rlabel metal2 386446 1836 386446 1836 0 ch_in[202]
rlabel metal2 389022 2040 389022 2040 0 ch_in[203]
rlabel metal2 391598 2142 391598 2142 0 ch_in[204]
rlabel metal2 394174 2074 394174 2074 0 ch_in[205]
rlabel metal2 396750 2006 396750 2006 0 ch_in[206]
rlabel metal2 408526 4624 408526 4624 0 ch_in[207]
rlabel metal1 409722 2414 409722 2414 0 ch_in[208]
rlabel metal2 404386 3808 404386 3808 0 ch_in[209]
rlabel metal2 210726 9350 210726 9350 0 ch_in[20]
rlabel metal2 407054 1870 407054 1870 0 ch_in[210]
rlabel metal2 409630 2176 409630 2176 0 ch_in[211]
rlabel metal1 411930 2414 411930 2414 0 ch_in[212]
rlabel metal1 414506 2414 414506 2414 0 ch_in[213]
rlabel metal2 417358 2108 417358 2108 0 ch_in[214]
rlabel metal1 419658 2414 419658 2414 0 ch_in[215]
rlabel metal2 422510 2142 422510 2142 0 ch_in[216]
rlabel metal1 425638 2550 425638 2550 0 ch_in[217]
rlabel metal2 427662 1972 427662 1972 0 ch_in[218]
rlabel metal1 446982 8296 446982 8296 0 ch_in[219]
rlabel metal1 25553 3366 25553 3366 0 ch_in[21]
rlabel metal2 456826 3264 456826 3264 0 ch_in[220]
rlabel metal2 480378 7276 480378 7276 0 ch_in[221]
rlabel metal1 439783 2482 439783 2482 0 ch_in[222]
rlabel metal2 440542 2006 440542 2006 0 ch_in[223]
rlabel metal2 443118 2074 443118 2074 0 ch_in[224]
rlabel metal1 445418 2414 445418 2414 0 ch_in[225]
rlabel metal2 448270 1972 448270 1972 0 ch_in[226]
rlabel metal1 450570 2414 450570 2414 0 ch_in[227]
rlabel metal1 453100 2414 453100 2414 0 ch_in[228]
rlabel metal1 455722 2414 455722 2414 0 ch_in[229]
rlabel metal1 28704 2278 28704 2278 0 ch_in[22]
rlabel metal2 475410 2210 475410 2210 0 ch_in[230]
rlabel metal1 460874 2414 460874 2414 0 ch_in[231]
rlabel metal2 463726 2142 463726 2142 0 ch_in[232]
rlabel metal2 483644 11356 483644 11356 0 ch_in[233]
rlabel metal2 468878 2040 468878 2040 0 ch_in[234]
rlabel metal2 471454 2108 471454 2108 0 ch_in[235]
rlabel metal2 473938 1938 473938 1938 0 ch_in[236]
rlabel metal1 476330 2414 476330 2414 0 ch_in[237]
rlabel metal1 478630 2380 478630 2380 0 ch_in[238]
rlabel metal1 481482 2414 481482 2414 0 ch_in[239]
rlabel metal1 29348 2822 29348 2822 0 ch_in[23]
rlabel metal1 484058 2414 484058 2414 0 ch_in[240]
rlabel metal1 486082 2414 486082 2414 0 ch_in[241]
rlabel metal1 488934 2448 488934 2448 0 ch_in[242]
rlabel metal1 491280 2414 491280 2414 0 ch_in[243]
rlabel metal1 493856 2414 493856 2414 0 ch_in[244]
rlabel metal1 496432 2414 496432 2414 0 ch_in[245]
rlabel metal1 499008 2414 499008 2414 0 ch_in[246]
rlabel metal1 501584 2414 501584 2414 0 ch_in[247]
rlabel metal1 504160 2414 504160 2414 0 ch_in[248]
rlabel metal1 506736 2414 506736 2414 0 ch_in[249]
rlabel metal2 186346 9180 186346 9180 0 ch_in[24]
rlabel metal2 509082 2788 509082 2788 0 ch_in[250]
rlabel metal2 511658 3978 511658 3978 0 ch_in[251]
rlabel metal2 514234 1428 514234 1428 0 ch_in[252]
rlabel metal1 30682 3502 30682 3502 0 ch_in[25]
rlabel metal2 34868 2108 34868 2108 0 ch_in[26]
rlabel metal2 205850 10455 205850 10455 0 ch_in[27]
rlabel metal1 34914 1054 34914 1054 0 ch_in[28]
rlabel metal1 37582 3434 37582 3434 0 ch_in[29]
rlabel metal2 187910 8806 187910 8806 0 ch_in[2]
rlabel metal2 149730 9384 149730 9384 0 ch_in[30]
rlabel metal1 38548 2890 38548 2890 0 ch_in[31]
rlabel metal2 42826 2108 42826 2108 0 ch_in[32]
rlabel metal1 153134 8942 153134 8942 0 ch_in[33]
rlabel metal1 44344 2278 44344 2278 0 ch_in[34]
rlabel metal2 45862 3196 45862 3196 0 ch_in[35]
rlabel metal2 157918 9996 157918 9996 0 ch_in[36]
rlabel metal2 43194 2210 43194 2210 0 ch_in[37]
rlabel metal1 41821 782 41821 782 0 ch_in[38]
rlabel metal1 160770 8942 160770 8942 0 ch_in[39]
rlabel metal2 4002 1802 4002 1802 0 ch_in[3]
rlabel metal1 43638 782 43638 782 0 ch_in[40]
rlabel metal1 45133 782 45133 782 0 ch_in[41]
rlabel metal1 165232 8466 165232 8466 0 ch_in[42]
rlabel metal2 49036 1326 49036 1326 0 ch_in[43]
rlabel metal1 48399 782 48399 782 0 ch_in[44]
rlabel metal2 195270 11492 195270 11492 0 ch_in[45]
rlabel metal1 50538 714 50538 714 0 ch_in[46]
rlabel metal1 60122 2822 60122 2822 0 ch_in[47]
rlabel metal2 173098 9554 173098 9554 0 ch_in[48]
rlabel metal1 61916 3366 61916 3366 0 ch_in[49]
rlabel metal2 6026 1598 6026 1598 0 ch_in[4]
rlabel metal1 65642 2822 65642 2822 0 ch_in[50]
rlabel metal2 176318 9520 176318 9520 0 ch_in[51]
rlabel metal1 63434 1190 63434 1190 0 ch_in[52]
rlabel metal2 62790 1326 62790 1326 0 ch_in[53]
rlabel metal1 180274 8942 180274 8942 0 ch_in[54]
rlabel metal2 60766 1054 60766 1054 0 ch_in[55]
rlabel metal1 61463 782 61463 782 0 ch_in[56]
rlabel metal2 195638 11322 195638 11322 0 ch_in[57]
rlabel metal1 63602 782 63602 782 0 ch_in[58]
rlabel metal2 65090 884 65090 884 0 ch_in[59]
rlabel metal2 6210 2074 6210 2074 0 ch_in[5]
rlabel metal1 187634 8908 187634 8908 0 ch_in[60]
rlabel metal1 66661 782 66661 782 0 ch_in[61]
rlabel via1 76590 867 76590 867 0 ch_in[62]
rlabel metal2 191498 8874 191498 8874 0 ch_in[63]
rlabel metal2 75670 1394 75670 1394 0 ch_in[64]
rlabel metal2 83674 3230 83674 3230 0 ch_in[65]
rlabel metal2 195914 10506 195914 10506 0 ch_in[66]
rlabel metal1 75762 1020 75762 1020 0 ch_in[67]
rlabel metal2 75026 680 75026 680 0 ch_in[68]
rlabel metal1 199134 9350 199134 9350 0 ch_in[69]
rlabel metal1 6700 782 6700 782 0 ch_in[6]
rlabel metal1 76390 782 76390 782 0 ch_in[70]
rlabel metal1 77713 782 77713 782 0 ch_in[71]
rlabel metal1 205758 9996 205758 9996 0 ch_in[72]
rlabel metal2 89838 1598 89838 1598 0 ch_in[73]
rlabel metal1 96968 2346 96968 2346 0 ch_in[74]
rlabel metal1 206034 9554 206034 9554 0 ch_in[75]
rlabel metal1 83198 714 83198 714 0 ch_in[76]
rlabel metal1 99613 3434 99613 3434 0 ch_in[77]
rlabel metal2 211094 10302 211094 10302 0 ch_in[78]
rlabel metal1 102304 3434 102304 3434 0 ch_in[79]
rlabel metal1 8832 2822 8832 2822 0 ch_in[7]
rlabel metal1 89930 1122 89930 1122 0 ch_in[80]
rlabel metal2 213854 9724 213854 9724 0 ch_in[81]
rlabel metal2 90114 833 90114 833 0 ch_in[82]
rlabel metal2 107594 3230 107594 3230 0 ch_in[83]
rlabel metal1 225078 10540 225078 10540 0 ch_in[84]
rlabel metal1 92965 782 92965 782 0 ch_in[85]
rlabel metal1 94100 782 94100 782 0 ch_in[86]
rlabel metal1 225170 10812 225170 10812 0 ch_in[87]
rlabel metal2 115322 2108 115322 2108 0 ch_in[88]
rlabel metal1 114954 3434 114954 3434 0 ch_in[89]
rlabel metal2 122590 9248 122590 9248 0 ch_in[8]
rlabel metal1 225308 9554 225308 9554 0 ch_in[90]
rlabel metal2 110722 833 110722 833 0 ch_in[91]
rlabel metal1 100586 714 100586 714 0 ch_in[92]
rlabel metal2 229126 9214 229126 9214 0 ch_in[93]
rlabel metal1 102875 782 102875 782 0 ch_in[94]
rlabel metal2 110814 1122 110814 1122 0 ch_in[95]
rlabel metal1 232944 9554 232944 9554 0 ch_in[96]
rlabel metal1 106117 782 106117 782 0 ch_in[97]
rlabel metal2 114954 1122 114954 1122 0 ch_in[98]
rlabel metal2 236854 9214 236854 9214 0 ch_in[99]
rlabel metal2 11362 2108 11362 2108 0 ch_in[9]
rlabel metal2 92138 8364 92138 8364 0 ch_out[0]
rlabel metal2 194718 3434 194718 3434 0 ch_out[100]
rlabel metal1 148672 5134 148672 5134 0 ch_out[101]
rlabel metal1 111511 782 111511 782 0 ch_out[102]
rlabel metal2 255898 7922 255898 7922 0 ch_out[103]
rlabel metal1 151110 3978 151110 3978 0 ch_out[104]
rlabel metal1 115444 782 115444 782 0 ch_out[105]
rlabel metal2 250838 9010 250838 9010 0 ch_out[106]
rlabel metal2 136482 2176 136482 2176 0 ch_out[107]
rlabel metal2 252034 7106 252034 7106 0 ch_out[108]
rlabel metal2 144946 1836 144946 1836 0 ch_out[109]
rlabel metal2 195546 11220 195546 11220 0 ch_out[10]
rlabel metal2 362066 9248 362066 9248 0 ch_out[110]
rlabel metal2 147798 1360 147798 1360 0 ch_out[111]
rlabel via2 363170 11475 363170 11475 0 ch_out[112]
rlabel metal1 137770 782 137770 782 0 ch_out[113]
rlabel metal2 267674 7378 267674 7378 0 ch_out[114]
rlabel metal2 148074 1020 148074 1020 0 ch_out[115]
rlabel metal2 365286 9112 365286 9112 0 ch_out[116]
rlabel metal2 161966 2108 161966 2108 0 ch_out[117]
rlabel metal1 275954 7752 275954 7752 0 ch_out[118]
rlabel metal2 167026 1105 167026 1105 0 ch_out[119]
rlabel metal1 195454 10948 195454 10948 0 ch_out[11]
rlabel metal1 276138 7888 276138 7888 0 ch_out[120]
rlabel metal2 167210 1411 167210 1411 0 ch_out[121]
rlabel metal2 368690 9384 368690 9384 0 ch_out[122]
rlabel via1 159022 459 159022 459 0 ch_out[123]
rlabel metal2 362342 6936 362342 6936 0 ch_out[124]
rlabel metal2 176410 1309 176410 1309 0 ch_out[125]
rlabel metal1 273240 6188 273240 6188 0 ch_out[126]
rlabel metal2 174846 782 174846 782 0 ch_out[127]
rlabel metal1 269330 5746 269330 5746 0 ch_out[128]
rlabel metal2 196006 2006 196006 2006 0 ch_out[129]
rlabel metal2 17342 1632 17342 1632 0 ch_out[12]
rlabel metal1 269422 6256 269422 6256 0 ch_out[130]
rlabel metal2 202814 1292 202814 1292 0 ch_out[131]
rlabel metal2 368506 7072 368506 7072 0 ch_out[132]
rlabel metal2 207966 1224 207966 1224 0 ch_out[133]
rlabel metal1 270434 5678 270434 5678 0 ch_out[134]
rlabel metal2 213118 1734 213118 1734 0 ch_out[135]
rlabel metal1 269146 5814 269146 5814 0 ch_out[136]
rlabel metal2 218270 1632 218270 1632 0 ch_out[137]
rlabel metal2 373474 6528 373474 6528 0 ch_out[138]
rlabel metal2 219742 578 219742 578 0 ch_out[139]
rlabel metal2 195362 10982 195362 10982 0 ch_out[13]
rlabel metal2 293894 6358 293894 6358 0 ch_out[140]
rlabel metal1 219420 952 219420 952 0 ch_out[141]
rlabel metal1 221115 782 221115 782 0 ch_out[142]
rlabel metal1 223314 782 223314 782 0 ch_out[143]
rlabel metal2 226458 986 226458 986 0 ch_out[144]
rlabel metal1 227546 782 227546 782 0 ch_out[145]
rlabel metal1 229699 782 229699 782 0 ch_out[146]
rlabel metal1 231341 782 231341 782 0 ch_out[147]
rlabel metal2 235014 1054 235014 1054 0 ch_out[148]
rlabel metal1 244490 1088 244490 1088 0 ch_out[149]
rlabel metal2 99958 9010 99958 9010 0 ch_out[14]
rlabel metal1 238011 782 238011 782 0 ch_out[150]
rlabel metal2 253874 1700 253874 1700 0 ch_out[151]
rlabel metal2 244398 1105 244398 1105 0 ch_out[152]
rlabel metal1 254426 1292 254426 1292 0 ch_out[153]
rlabel metal2 248078 918 248078 918 0 ch_out[154]
rlabel metal2 263626 1241 263626 1241 0 ch_out[155]
rlabel metal2 267214 1700 267214 1700 0 ch_out[156]
rlabel metal2 268042 1734 268042 1734 0 ch_out[157]
rlabel metal2 267858 1326 267858 1326 0 ch_out[158]
rlabel metal1 273240 2312 273240 2312 0 ch_out[159]
rlabel metal1 100142 6698 100142 6698 0 ch_out[15]
rlabel metal2 271630 1258 271630 1258 0 ch_out[160]
rlabel metal2 274114 799 274114 799 0 ch_out[161]
rlabel metal1 264541 646 264541 646 0 ch_out[162]
rlabel metal1 266784 714 266784 714 0 ch_out[163]
rlabel metal1 268325 714 268325 714 0 ch_out[164]
rlabel metal1 270933 782 270933 782 0 ch_out[165]
rlabel metal2 289938 1836 289938 1836 0 ch_out[166]
rlabel metal2 291226 2108 291226 2108 0 ch_out[167]
rlabel metal2 295274 1870 295274 1870 0 ch_out[168]
rlabel metal2 291778 1666 291778 1666 0 ch_out[169]
rlabel metal1 17571 782 17571 782 0 ch_out[16]
rlabel metal1 302749 2618 302749 2618 0 ch_out[170]
rlabel metal1 284080 714 284080 714 0 ch_out[171]
rlabel metal1 286323 782 286323 782 0 ch_out[172]
rlabel via1 289754 901 289754 901 0 ch_out[173]
rlabel metal1 290428 782 290428 782 0 ch_out[174]
rlabel metal2 309258 1343 309258 1343 0 ch_out[175]
rlabel metal1 302450 884 302450 884 0 ch_out[176]
rlabel metal2 302358 1394 302358 1394 0 ch_out[177]
rlabel metal1 323886 2312 323886 2312 0 ch_out[178]
rlabel metal2 326462 1224 326462 1224 0 ch_out[179]
rlabel metal2 100694 9622 100694 9622 0 ch_out[17]
rlabel metal2 329038 1258 329038 1258 0 ch_out[180]
rlabel metal2 331246 1632 331246 1632 0 ch_out[181]
rlabel metal2 334190 1666 334190 1666 0 ch_out[182]
rlabel metal2 336766 1700 336766 1700 0 ch_out[183]
rlabel metal1 325680 816 325680 816 0 ch_out[184]
rlabel metal2 341918 1598 341918 1598 0 ch_out[185]
rlabel metal2 344494 1156 344494 1156 0 ch_out[186]
rlabel metal2 347070 1190 347070 1190 0 ch_out[187]
rlabel metal1 357758 782 357758 782 0 ch_out[188]
rlabel metal2 352222 2040 352222 2040 0 ch_out[189]
rlabel metal2 101982 8534 101982 8534 0 ch_out[18]
rlabel metal2 358018 1700 358018 1700 0 ch_out[190]
rlabel metal2 357374 1598 357374 1598 0 ch_out[191]
rlabel metal2 359950 1632 359950 1632 0 ch_out[192]
rlabel metal2 367126 1666 367126 1666 0 ch_out[193]
rlabel metal2 365102 1870 365102 1870 0 ch_out[194]
rlabel metal1 374387 782 374387 782 0 ch_out[195]
rlabel metal1 377459 782 377459 782 0 ch_out[196]
rlabel metal1 379654 782 379654 782 0 ch_out[197]
rlabel metal1 381379 782 381379 782 0 ch_out[198]
rlabel metal1 383943 782 383943 782 0 ch_out[199]
rlabel metal2 101890 7769 101890 7769 0 ch_out[19]
rlabel metal2 92230 9656 92230 9656 0 ch_out[1]
rlabel metal1 385634 782 385634 782 0 ch_out[200]
rlabel metal1 388095 782 388095 782 0 ch_out[201]
rlabel metal1 390625 782 390625 782 0 ch_out[202]
rlabel metal1 392350 782 392350 782 0 ch_out[203]
rlabel metal1 394489 782 394489 782 0 ch_out[204]
rlabel metal1 396168 782 396168 782 0 ch_out[205]
rlabel metal1 398459 782 398459 782 0 ch_out[206]
rlabel metal1 400837 782 400837 782 0 ch_out[207]
rlabel metal2 402454 1530 402454 1530 0 ch_out[208]
rlabel metal1 405877 714 405877 714 0 ch_out[209]
rlabel metal1 21972 782 21972 782 0 ch_out[20]
rlabel metal1 407139 782 407139 782 0 ch_out[210]
rlabel metal1 409508 782 409508 782 0 ch_out[211]
rlabel metal1 411887 782 411887 782 0 ch_out[212]
rlabel metal1 414269 782 414269 782 0 ch_out[213]
rlabel metal1 416592 782 416592 782 0 ch_out[214]
rlabel metal1 419029 782 419029 782 0 ch_out[215]
rlabel metal1 421405 782 421405 782 0 ch_out[216]
rlabel metal1 423414 782 423414 782 0 ch_out[217]
rlabel metal1 425737 782 425737 782 0 ch_out[218]
rlabel metal1 427659 782 427659 782 0 ch_out[219]
rlabel metal2 102902 8840 102902 8840 0 ch_out[21]
rlabel metal1 430130 782 430130 782 0 ch_out[220]
rlabel metal1 431841 782 431841 782 0 ch_out[221]
rlabel metal1 434373 782 434373 782 0 ch_out[222]
rlabel metal1 436570 782 436570 782 0 ch_out[223]
rlabel metal2 442382 1666 442382 1666 0 ch_out[224]
rlabel metal2 444406 1598 444406 1598 0 ch_out[225]
rlabel metal1 442872 782 442872 782 0 ch_out[226]
rlabel metal1 445885 782 445885 782 0 ch_out[227]
rlabel metal1 447150 782 447150 782 0 ch_out[228]
rlabel metal1 449243 714 449243 714 0 ch_out[229]
rlabel metal2 196374 646 196374 646 0 ch_out[22]
rlabel metal1 452509 782 452509 782 0 ch_out[230]
rlabel metal1 454602 782 454602 782 0 ch_out[231]
rlabel metal1 455773 782 455773 782 0 ch_out[232]
rlabel metal1 458075 782 458075 782 0 ch_out[233]
rlabel metal2 466486 1666 466486 1666 0 ch_out[234]
rlabel metal2 469246 1700 469246 1700 0 ch_out[235]
rlabel metal2 471914 1632 471914 1632 0 ch_out[236]
rlabel metal1 467666 714 467666 714 0 ch_out[237]
rlabel metal1 470810 850 470810 850 0 ch_out[238]
rlabel metal1 472005 782 472005 782 0 ch_out[239]
rlabel metal2 195270 10846 195270 10846 0 ch_out[23]
rlabel metal2 483598 1632 483598 1632 0 ch_out[240]
rlabel metal2 486174 1564 486174 1564 0 ch_out[241]
rlabel metal2 488750 1700 488750 1700 0 ch_out[242]
rlabel metal2 481574 1054 481574 1054 0 ch_out[243]
rlabel metal1 482869 782 482869 782 0 ch_out[244]
rlabel metal1 485065 782 485065 782 0 ch_out[245]
rlabel metal1 486282 714 486282 714 0 ch_out[246]
rlabel metal2 500342 1632 500342 1632 0 ch_out[247]
rlabel metal2 502366 1666 502366 1666 0 ch_out[248]
rlabel metal2 505126 1700 505126 1700 0 ch_out[249]
rlabel metal2 32798 1700 32798 1700 0 ch_out[24]
rlabel metal1 496025 782 496025 782 0 ch_out[250]
rlabel metal1 497750 782 497750 782 0 ch_out[251]
rlabel metal1 488750 2380 488750 2380 0 ch_out[252]
rlabel metal1 108514 6766 108514 6766 0 ch_out[25]
rlabel metal2 106214 8466 106214 8466 0 ch_out[26]
rlabel metal1 33626 3638 33626 3638 0 ch_out[27]
rlabel metal2 194994 10438 194994 10438 0 ch_out[28]
rlabel metal2 184230 9843 184230 9843 0 ch_out[29]
rlabel metal1 2779 782 2779 782 0 ch_out[2]
rlabel metal1 33150 714 33150 714 0 ch_out[30]
rlabel metal2 109526 6528 109526 6528 0 ch_out[31]
rlabel metal2 109894 8092 109894 8092 0 ch_out[32]
rlabel metal1 41124 3366 41124 3366 0 ch_out[33]
rlabel metal1 113298 6392 113298 6392 0 ch_out[34]
rlabel metal2 110906 6256 110906 6256 0 ch_out[35]
rlabel metal1 43378 918 43378 918 0 ch_out[36]
rlabel metal2 112838 8466 112838 8466 0 ch_out[37]
rlabel via1 113390 6443 113390 6443 0 ch_out[38]
rlabel metal1 42917 782 42917 782 0 ch_out[39]
rlabel metal2 92874 9520 92874 9520 0 ch_out[3]
rlabel metal2 114126 6052 114126 6052 0 ch_out[40]
rlabel metal2 114218 6647 114218 6647 0 ch_out[41]
rlabel metal1 46297 782 46297 782 0 ch_out[42]
rlabel metal1 117047 6834 117047 6834 0 ch_out[43]
rlabel metal1 130870 5678 130870 5678 0 ch_out[44]
rlabel metal1 57638 3366 57638 3366 0 ch_out[45]
rlabel metal2 224986 9044 224986 9044 0 ch_out[46]
rlabel metal2 225446 8976 225446 8976 0 ch_out[47]
rlabel metal1 61134 1462 61134 1462 0 ch_out[48]
rlabel metal2 118542 6698 118542 6698 0 ch_out[49]
rlabel metal2 186254 10081 186254 10081 0 ch_out[4]
rlabel metal1 135746 5814 135746 5814 0 ch_out[50]
rlabel metal2 63526 2312 63526 2312 0 ch_out[51]
rlabel metal1 135470 5746 135470 5746 0 ch_out[52]
rlabel metal2 228482 9588 228482 9588 0 ch_out[53]
rlabel metal2 63250 1122 63250 1122 0 ch_out[54]
rlabel metal2 229862 8772 229862 8772 0 ch_out[55]
rlabel metal2 230506 7565 230506 7565 0 ch_out[56]
rlabel metal1 62507 714 62507 714 0 ch_out[57]
rlabel metal2 231426 8704 231426 8704 0 ch_out[58]
rlabel metal2 231886 8806 231886 8806 0 ch_out[59]
rlabel metal2 93518 7667 93518 7667 0 ch_out[5]
rlabel metal1 76130 1224 76130 1224 0 ch_out[60]
rlabel metal2 233450 8789 233450 8789 0 ch_out[61]
rlabel metal1 148166 5168 148166 5168 0 ch_out[62]
rlabel metal2 75762 1326 75762 1326 0 ch_out[63]
rlabel metal2 128110 4658 128110 4658 0 ch_out[64]
rlabel metal2 186622 8704 186622 8704 0 ch_out[65]
rlabel metal1 75946 952 75946 952 0 ch_out[66]
rlabel metal2 236302 8738 236302 8738 0 ch_out[67]
rlabel metal2 130870 4964 130870 4964 0 ch_out[68]
rlabel metal1 75470 782 75470 782 0 ch_out[69]
rlabel metal2 176686 9231 176686 9231 0 ch_out[6]
rlabel metal1 131698 5100 131698 5100 0 ch_out[70]
rlabel metal2 130962 5933 130962 5933 0 ch_out[71]
rlabel metal1 78805 782 78805 782 0 ch_out[72]
rlabel metal2 132066 6766 132066 6766 0 ch_out[73]
rlabel metal2 133538 4913 133538 4913 0 ch_out[74]
rlabel metal1 82094 782 82094 782 0 ch_out[75]
rlabel metal1 134642 5304 134642 5304 0 ch_out[76]
rlabel metal2 134458 5882 134458 5882 0 ch_out[77]
rlabel metal1 85383 782 85383 782 0 ch_out[78]
rlabel metal2 135562 5899 135562 5899 0 ch_out[79]
rlabel metal2 186714 9146 186714 9146 0 ch_out[7]
rlabel metal2 138138 4726 138138 4726 0 ch_out[80]
rlabel metal1 99590 1020 99590 1020 0 ch_out[81]
rlabel metal2 244490 7888 244490 7888 0 ch_out[82]
rlabel metal2 137862 4777 137862 4777 0 ch_out[83]
rlabel metal1 91869 782 91869 782 0 ch_out[84]
rlabel metal2 246146 9622 246146 9622 0 ch_out[85]
rlabel metal2 246698 7956 246698 7956 0 ch_out[86]
rlabel metal1 95158 782 95158 782 0 ch_out[87]
rlabel metal2 247710 7990 247710 7990 0 ch_out[88]
rlabel metal2 248538 8245 248538 8245 0 ch_out[89]
rlabel metal1 9217 782 9217 782 0 ch_out[8]
rlabel metal1 98447 782 98447 782 0 ch_out[90]
rlabel metal2 249366 7752 249366 7752 0 ch_out[91]
rlabel metal2 250010 7106 250010 7106 0 ch_out[92]
rlabel metal2 109066 1972 109066 1972 0 ch_out[93]
rlabel metal1 151800 4080 151800 4080 0 ch_out[94]
rlabel metal2 251574 7769 251574 7769 0 ch_out[95]
rlabel metal2 109250 2040 109250 2040 0 ch_out[96]
rlabel metal2 252770 7905 252770 7905 0 ch_out[97]
rlabel via1 151202 3995 151202 3995 0 ch_out[98]
rlabel metal1 113850 782 113850 782 0 ch_out[99]
rlabel metal2 195178 10370 195178 10370 0 ch_out[9]
rlabel metal2 63526 6120 63526 6120 0 net1
rlabel metal2 112654 3604 112654 3604 0 net10
rlabel metal2 210266 9333 210266 9333 0 net100
rlabel metal2 114770 1003 114770 1003 0 net101
rlabel metal1 192878 2822 192878 2822 0 net102
rlabel via1 89654 3485 89654 3485 0 net103
rlabel metal2 194718 9316 194718 9316 0 net104
rlabel metal2 81926 3434 81926 3434 0 net105
rlabel metal2 79902 1921 79902 1921 0 net106
rlabel metal2 74750 6460 74750 6460 0 net107
rlabel metal2 179446 6222 179446 6222 0 net108
rlabel metal1 67160 3706 67160 3706 0 net109
rlabel metal2 109986 3944 109986 3944 0 net11
rlabel metal2 64446 2193 64446 2193 0 net110
rlabel metal1 59018 3502 59018 3502 0 net111
rlabel metal1 56396 2414 56396 2414 0 net112
rlabel metal2 160126 8568 160126 8568 0 net113
rlabel metal2 48990 2533 48990 2533 0 net114
rlabel metal1 43562 3502 43562 3502 0 net115
rlabel metal1 149132 8398 149132 8398 0 net116
rlabel metal2 5198 3910 5198 3910 0 net117
rlabel metal2 36110 3604 36110 3604 0 net118
rlabel metal1 33258 2414 33258 2414 0 net119
rlabel metal2 107502 3162 107502 3162 0 net12
rlabel metal2 136666 5083 136666 5083 0 net120
rlabel metal1 102166 7276 102166 7276 0 net121
rlabel metal2 283130 1326 283130 1326 0 net122
rlabel metal2 380834 9248 380834 9248 0 net123
rlabel metal1 272826 2414 272826 2414 0 net124
rlabel metal1 270250 2414 270250 2414 0 net125
rlabel metal2 267950 1768 267950 1768 0 net126
rlabel metal1 265098 2414 265098 2414 0 net127
rlabel metal2 368598 9758 368598 9758 0 net128
rlabel metal1 341642 9384 341642 9384 0 net129
rlabel metal2 137954 4352 137954 4352 0 net13
rlabel metal2 363722 6460 363722 6460 0 net130
rlabel metal1 360732 9486 360732 9486 0 net131
rlabel metal1 252172 2414 252172 2414 0 net132
rlabel metal1 249642 2414 249642 2414 0 net133
rlabel metal1 247020 2414 247020 2414 0 net134
rlabel metal2 312938 6562 312938 6562 0 net135
rlabel metal2 349370 9010 349370 9010 0 net136
rlabel metal2 346794 10438 346794 10438 0 net137
rlabel metal2 344126 8466 344126 8466 0 net138
rlabel metal1 341550 9452 341550 9452 0 net139
rlabel metal2 110814 1496 110814 1496 0 net14
rlabel metal2 338974 9316 338974 9316 0 net140
rlabel metal2 336306 10064 336306 10064 0 net141
rlabel metal1 326738 8840 326738 8840 0 net142
rlabel metal1 218684 2414 218684 2414 0 net143
rlabel metal1 213532 2414 213532 2414 0 net144
rlabel metal1 208380 2414 208380 2414 0 net145
rlabel metal2 311282 9928 311282 9928 0 net146
rlabel metal2 18078 3944 18078 3944 0 net147
rlabel metal1 198076 2414 198076 2414 0 net148
rlabel metal2 194672 3876 194672 3876 0 net149
rlabel metal2 9614 4488 9614 4488 0 net15
rlabel via1 195178 3621 195178 3621 0 net150
rlabel metal2 291226 7531 291226 7531 0 net151
rlabel metal1 195270 3604 195270 3604 0 net152
rlabel metal1 200100 680 200100 680 0 net153
rlabel metal2 276046 8126 276046 8126 0 net154
rlabel metal2 270986 7667 270986 7667 0 net155
rlabel metal2 196098 1258 196098 1258 0 net156
rlabel metal2 152030 2142 152030 2142 0 net157
rlabel via2 146878 2363 146878 2363 0 net158
rlabel metal2 187358 2159 187358 2159 0 net159
rlabel metal2 102350 3910 102350 3910 0 net16
rlabel metal1 136298 3502 136298 3502 0 net160
rlabel metal2 133998 1972 133998 1972 0 net161
rlabel metal2 99774 3230 99774 3230 0 net17
rlabel metal2 134366 4828 134366 4828 0 net18
rlabel metal2 97198 3672 97198 3672 0 net19
rlabel metal2 132388 1462 132388 1462 0 net2
rlabel metal2 94622 3264 94622 3264 0 net20
rlabel metal2 92046 3128 92046 3128 0 net21
rlabel metal1 92230 2618 92230 2618 0 net22
rlabel metal2 59202 3672 59202 3672 0 net23
rlabel metal2 94162 3536 94162 3536 0 net24
rlabel metal2 86894 3230 86894 3230 0 net25
rlabel metal2 84318 3740 84318 3740 0 net26
rlabel metal2 84318 1904 84318 1904 0 net27
rlabel metal2 81742 3655 81742 3655 0 net28
rlabel metal2 79074 3740 79074 3740 0 net29
rlabel metal1 133170 3604 133170 3604 0 net3
rlabel metal2 6854 4420 6854 4420 0 net30
rlabel metal2 76498 3706 76498 3706 0 net31
rlabel metal2 76590 3842 76590 3842 0 net32
rlabel metal2 74014 3706 74014 3706 0 net33
rlabel metal2 71438 3638 71438 3638 0 net34
rlabel metal2 120474 4998 120474 4998 0 net35
rlabel metal2 68862 3842 68862 3842 0 net36
rlabel metal2 66286 1870 66286 1870 0 net37
rlabel metal2 75578 2074 75578 2074 0 net38
rlabel metal1 117576 6086 117576 6086 0 net39
rlabel metal2 133170 3808 133170 3808 0 net4
rlabel metal1 61134 3604 61134 3604 0 net40
rlabel metal2 61134 2890 61134 2890 0 net41
rlabel metal2 58558 2108 58558 2108 0 net42
rlabel metal2 55982 3077 55982 3077 0 net43
rlabel via1 62974 3451 62974 3451 0 net44
rlabel metal2 53406 2142 53406 2142 0 net45
rlabel metal2 4462 3842 4462 3842 0 net46
rlabel metal2 50830 1938 50830 1938 0 net47
rlabel metal2 48254 3876 48254 3876 0 net48
rlabel metal1 99498 6290 99498 6290 0 net49
rlabel metal2 122958 2108 122958 2108 0 net5
rlabel metal1 110124 6290 110124 6290 0 net50
rlabel metal1 44321 2550 44321 2550 0 net51
rlabel metal1 60030 3672 60030 3672 0 net52
rlabel metal2 47426 4590 47426 4590 0 net53
rlabel metal1 106766 5678 106766 5678 0 net54
rlabel metal2 105110 5814 105110 5814 0 net55
rlabel metal2 32798 3417 32798 3417 0 net56
rlabel metal1 102442 6800 102442 6800 0 net57
rlabel metal2 102626 5984 102626 5984 0 net58
rlabel metal2 101246 4794 101246 4794 0 net59
rlabel metal2 120382 2074 120382 2074 0 net6
rlabel metal2 1886 4930 1886 4930 0 net60
rlabel metal2 35926 5814 35926 5814 0 net61
rlabel metal1 100188 6086 100188 6086 0 net62
rlabel metal2 22494 5814 22494 5814 0 net63
rlabel metal2 19918 4726 19918 4726 0 net64
rlabel metal2 42918 4318 42918 4318 0 net65
rlabel metal2 225998 2040 225998 2040 0 net66
rlabel metal2 17342 4998 17342 4998 0 net67
rlabel metal2 220846 2074 220846 2074 0 net68
rlabel metal2 215694 2108 215694 2108 0 net69
rlabel metal2 133078 3808 133078 3808 0 net7
rlabel metal2 210542 2856 210542 2856 0 net70
rlabel metal2 210450 3910 210450 3910 0 net71
rlabel metal2 200238 2142 200238 2142 0 net72
rlabel metal2 195086 2176 195086 2176 0 net73
rlabel metal2 195362 1904 195362 1904 0 net74
rlabel metal1 222778 2550 222778 2550 0 net75
rlabel metal2 179630 1904 179630 1904 0 net76
rlabel metal2 174478 2193 174478 2193 0 net77
rlabel metal2 14766 5712 14766 5712 0 net78
rlabel via2 169326 2261 169326 2261 0 net79
rlabel metal2 115138 4420 115138 4420 0 net8
rlabel metal2 164174 2465 164174 2465 0 net80
rlabel metal2 158930 2465 158930 2465 0 net81
rlabel metal1 203918 2482 203918 2482 0 net82
rlabel metal2 148626 1972 148626 1972 0 net83
rlabel metal2 14766 2040 14766 2040 0 net84
rlabel metal2 191130 1955 191130 1955 0 net85
rlabel metal1 249596 7174 249596 7174 0 net86
rlabel metal1 136022 2346 136022 2346 0 net87
rlabel metal2 149178 3808 149178 3808 0 net88
rlabel metal2 148074 5100 148074 5100 0 net89
rlabel metal2 115230 1938 115230 1938 0 net9
rlabel metal1 148212 3570 148212 3570 0 net90
rlabel metal1 33626 2380 33626 2380 0 net91
rlabel metal1 135838 3400 135838 3400 0 net92
rlabel metal1 232162 9486 232162 9486 0 net93
rlabel metal2 228298 6137 228298 6137 0 net94
rlabel metal1 118266 2414 118266 2414 0 net95
rlabel metal2 43010 7004 43010 7004 0 net96
rlabel metal1 112838 3536 112838 3536 0 net97
rlabel metal1 110538 2414 110538 2414 0 net98
rlabel via2 105662 3451 105662 3451 0 net99
<< properties >>
string FIXED_BBOX 0 0 530000 12000
<< end >>
